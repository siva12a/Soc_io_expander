magic
tech sky130A
magscale 1 2
timestamp 1623941690
<< obsli1 >>
rect 1104 17 98808 39627
<< obsm1 >>
rect 106 8 99898 39636
<< metal2 >>
rect 386 39200 442 40000
rect 1214 39200 1270 40000
rect 2134 39200 2190 40000
rect 2962 39200 3018 40000
rect 3882 39200 3938 40000
rect 4710 39200 4766 40000
rect 5630 39200 5686 40000
rect 6458 39200 6514 40000
rect 7378 39200 7434 40000
rect 8206 39200 8262 40000
rect 9126 39200 9182 40000
rect 9954 39200 10010 40000
rect 10874 39200 10930 40000
rect 11702 39200 11758 40000
rect 12622 39200 12678 40000
rect 13542 39200 13598 40000
rect 14370 39200 14426 40000
rect 15290 39200 15346 40000
rect 16118 39200 16174 40000
rect 17038 39200 17094 40000
rect 17866 39200 17922 40000
rect 18786 39200 18842 40000
rect 19614 39200 19670 40000
rect 20534 39200 20590 40000
rect 21362 39200 21418 40000
rect 22282 39200 22338 40000
rect 23110 39200 23166 40000
rect 24030 39200 24086 40000
rect 24858 39200 24914 40000
rect 25778 39200 25834 40000
rect 26698 39200 26754 40000
rect 27526 39200 27582 40000
rect 28446 39200 28502 40000
rect 29274 39200 29330 40000
rect 30194 39200 30250 40000
rect 31022 39200 31078 40000
rect 31942 39200 31998 40000
rect 32770 39200 32826 40000
rect 33690 39200 33746 40000
rect 34518 39200 34574 40000
rect 35438 39200 35494 40000
rect 36266 39200 36322 40000
rect 37186 39200 37242 40000
rect 38106 39200 38162 40000
rect 38934 39200 38990 40000
rect 39854 39200 39910 40000
rect 40682 39200 40738 40000
rect 41602 39200 41658 40000
rect 42430 39200 42486 40000
rect 43350 39200 43406 40000
rect 44178 39200 44234 40000
rect 45098 39200 45154 40000
rect 45926 39200 45982 40000
rect 46846 39200 46902 40000
rect 47674 39200 47730 40000
rect 48594 39200 48650 40000
rect 49422 39200 49478 40000
rect 50342 39200 50398 40000
rect 51262 39200 51318 40000
rect 52090 39200 52146 40000
rect 53010 39200 53066 40000
rect 53838 39200 53894 40000
rect 54758 39200 54814 40000
rect 55586 39200 55642 40000
rect 56506 39200 56562 40000
rect 57334 39200 57390 40000
rect 58254 39200 58310 40000
rect 59082 39200 59138 40000
rect 60002 39200 60058 40000
rect 60830 39200 60886 40000
rect 61750 39200 61806 40000
rect 62578 39200 62634 40000
rect 63498 39200 63554 40000
rect 64418 39200 64474 40000
rect 65246 39200 65302 40000
rect 66166 39200 66222 40000
rect 66994 39200 67050 40000
rect 67914 39200 67970 40000
rect 68742 39200 68798 40000
rect 69662 39200 69718 40000
rect 70490 39200 70546 40000
rect 71410 39200 71466 40000
rect 72238 39200 72294 40000
rect 73158 39200 73214 40000
rect 73986 39200 74042 40000
rect 74906 39200 74962 40000
rect 75826 39200 75882 40000
rect 76654 39200 76710 40000
rect 77574 39200 77630 40000
rect 78402 39200 78458 40000
rect 79322 39200 79378 40000
rect 80150 39200 80206 40000
rect 81070 39200 81126 40000
rect 81898 39200 81954 40000
rect 82818 39200 82874 40000
rect 83646 39200 83702 40000
rect 84566 39200 84622 40000
rect 85394 39200 85450 40000
rect 86314 39200 86370 40000
rect 87142 39200 87198 40000
rect 88062 39200 88118 40000
rect 88982 39200 89038 40000
rect 89810 39200 89866 40000
rect 90730 39200 90786 40000
rect 91558 39200 91614 40000
rect 92478 39200 92534 40000
rect 93306 39200 93362 40000
rect 94226 39200 94282 40000
rect 95054 39200 95110 40000
rect 95974 39200 96030 40000
rect 96802 39200 96858 40000
rect 97722 39200 97778 40000
rect 98550 39200 98606 40000
rect 99470 39200 99526 40000
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 13910 0 13966 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19338 0 19394 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36450 0 36506 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38658 0 38714 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40130 0 40186 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62026 0 62082 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63498 0 63554 800
rect 63682 0 63738 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65338 0 65394 800
rect 65522 0 65578 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67546 0 67602 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70766 0 70822 800
rect 71042 0 71098 800
rect 71226 0 71282 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73250 0 73306 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73802 0 73858 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74906 0 74962 800
rect 75090 0 75146 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76286 0 76342 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78770 0 78826 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81346 0 81402 800
rect 81530 0 81586 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83002 0 83058 800
rect 83186 0 83242 800
rect 83370 0 83426 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85026 0 85082 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88522 0 88578 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89258 0 89314 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 92938 0 92994 800
rect 93122 0 93178 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95146 0 95202 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< obsm2 >>
rect 112 39144 330 39642
rect 498 39144 1158 39642
rect 1326 39144 2078 39642
rect 2246 39144 2906 39642
rect 3074 39144 3826 39642
rect 3994 39144 4654 39642
rect 4822 39144 5574 39642
rect 5742 39144 6402 39642
rect 6570 39144 7322 39642
rect 7490 39144 8150 39642
rect 8318 39144 9070 39642
rect 9238 39144 9898 39642
rect 10066 39144 10818 39642
rect 10986 39144 11646 39642
rect 11814 39144 12566 39642
rect 12734 39144 13486 39642
rect 13654 39144 14314 39642
rect 14482 39144 15234 39642
rect 15402 39144 16062 39642
rect 16230 39144 16982 39642
rect 17150 39144 17810 39642
rect 17978 39144 18730 39642
rect 18898 39144 19558 39642
rect 19726 39144 20478 39642
rect 20646 39144 21306 39642
rect 21474 39144 22226 39642
rect 22394 39144 23054 39642
rect 23222 39144 23974 39642
rect 24142 39144 24802 39642
rect 24970 39144 25722 39642
rect 25890 39144 26642 39642
rect 26810 39144 27470 39642
rect 27638 39144 28390 39642
rect 28558 39144 29218 39642
rect 29386 39144 30138 39642
rect 30306 39144 30966 39642
rect 31134 39144 31886 39642
rect 32054 39144 32714 39642
rect 32882 39144 33634 39642
rect 33802 39144 34462 39642
rect 34630 39144 35382 39642
rect 35550 39144 36210 39642
rect 36378 39144 37130 39642
rect 37298 39144 38050 39642
rect 38218 39144 38878 39642
rect 39046 39144 39798 39642
rect 39966 39144 40626 39642
rect 40794 39144 41546 39642
rect 41714 39144 42374 39642
rect 42542 39144 43294 39642
rect 43462 39144 44122 39642
rect 44290 39144 45042 39642
rect 45210 39144 45870 39642
rect 46038 39144 46790 39642
rect 46958 39144 47618 39642
rect 47786 39144 48538 39642
rect 48706 39144 49366 39642
rect 49534 39144 50286 39642
rect 50454 39144 51206 39642
rect 51374 39144 52034 39642
rect 52202 39144 52954 39642
rect 53122 39144 53782 39642
rect 53950 39144 54702 39642
rect 54870 39144 55530 39642
rect 55698 39144 56450 39642
rect 56618 39144 57278 39642
rect 57446 39144 58198 39642
rect 58366 39144 59026 39642
rect 59194 39144 59946 39642
rect 60114 39144 60774 39642
rect 60942 39144 61694 39642
rect 61862 39144 62522 39642
rect 62690 39144 63442 39642
rect 63610 39144 64362 39642
rect 64530 39144 65190 39642
rect 65358 39144 66110 39642
rect 66278 39144 66938 39642
rect 67106 39144 67858 39642
rect 68026 39144 68686 39642
rect 68854 39144 69606 39642
rect 69774 39144 70434 39642
rect 70602 39144 71354 39642
rect 71522 39144 72182 39642
rect 72350 39144 73102 39642
rect 73270 39144 73930 39642
rect 74098 39144 74850 39642
rect 75018 39144 75770 39642
rect 75938 39144 76598 39642
rect 76766 39144 77518 39642
rect 77686 39144 78346 39642
rect 78514 39144 79266 39642
rect 79434 39144 80094 39642
rect 80262 39144 81014 39642
rect 81182 39144 81842 39642
rect 82010 39144 82762 39642
rect 82930 39144 83590 39642
rect 83758 39144 84510 39642
rect 84678 39144 85338 39642
rect 85506 39144 86258 39642
rect 86426 39144 87086 39642
rect 87254 39144 88006 39642
rect 88174 39144 88926 39642
rect 89094 39144 89754 39642
rect 89922 39144 90674 39642
rect 90842 39144 91502 39642
rect 91670 39144 92422 39642
rect 92590 39144 93250 39642
rect 93418 39144 94170 39642
rect 94338 39144 94998 39642
rect 95166 39144 95918 39642
rect 96086 39144 96746 39642
rect 96914 39144 97666 39642
rect 97834 39144 98494 39642
rect 98662 39144 99414 39642
rect 99582 39144 99892 39642
rect 112 856 99892 39144
rect 222 2 238 856
rect 406 2 422 856
rect 590 2 606 856
rect 774 2 790 856
rect 958 2 1066 856
rect 1234 2 1250 856
rect 1418 2 1434 856
rect 1602 2 1618 856
rect 1786 2 1802 856
rect 1970 2 2078 856
rect 2246 2 2262 856
rect 2430 2 2446 856
rect 2614 2 2630 856
rect 2798 2 2814 856
rect 2982 2 3090 856
rect 3258 2 3274 856
rect 3442 2 3458 856
rect 3626 2 3642 856
rect 3810 2 3826 856
rect 3994 2 4102 856
rect 4270 2 4286 856
rect 4454 2 4470 856
rect 4638 2 4654 856
rect 4822 2 4930 856
rect 5098 2 5114 856
rect 5282 2 5298 856
rect 5466 2 5482 856
rect 5650 2 5666 856
rect 5834 2 5942 856
rect 6110 2 6126 856
rect 6294 2 6310 856
rect 6478 2 6494 856
rect 6662 2 6678 856
rect 6846 2 6954 856
rect 7122 2 7138 856
rect 7306 2 7322 856
rect 7490 2 7506 856
rect 7674 2 7690 856
rect 7858 2 7966 856
rect 8134 2 8150 856
rect 8318 2 8334 856
rect 8502 2 8518 856
rect 8686 2 8794 856
rect 8962 2 8978 856
rect 9146 2 9162 856
rect 9330 2 9346 856
rect 9514 2 9530 856
rect 9698 2 9806 856
rect 9974 2 9990 856
rect 10158 2 10174 856
rect 10342 2 10358 856
rect 10526 2 10542 856
rect 10710 2 10818 856
rect 10986 2 11002 856
rect 11170 2 11186 856
rect 11354 2 11370 856
rect 11538 2 11554 856
rect 11722 2 11830 856
rect 11998 2 12014 856
rect 12182 2 12198 856
rect 12366 2 12382 856
rect 12550 2 12566 856
rect 12734 2 12842 856
rect 13010 2 13026 856
rect 13194 2 13210 856
rect 13378 2 13394 856
rect 13562 2 13670 856
rect 13838 2 13854 856
rect 14022 2 14038 856
rect 14206 2 14222 856
rect 14390 2 14406 856
rect 14574 2 14682 856
rect 14850 2 14866 856
rect 15034 2 15050 856
rect 15218 2 15234 856
rect 15402 2 15418 856
rect 15586 2 15694 856
rect 15862 2 15878 856
rect 16046 2 16062 856
rect 16230 2 16246 856
rect 16414 2 16430 856
rect 16598 2 16706 856
rect 16874 2 16890 856
rect 17058 2 17074 856
rect 17242 2 17258 856
rect 17426 2 17534 856
rect 17702 2 17718 856
rect 17886 2 17902 856
rect 18070 2 18086 856
rect 18254 2 18270 856
rect 18438 2 18546 856
rect 18714 2 18730 856
rect 18898 2 18914 856
rect 19082 2 19098 856
rect 19266 2 19282 856
rect 19450 2 19558 856
rect 19726 2 19742 856
rect 19910 2 19926 856
rect 20094 2 20110 856
rect 20278 2 20294 856
rect 20462 2 20570 856
rect 20738 2 20754 856
rect 20922 2 20938 856
rect 21106 2 21122 856
rect 21290 2 21306 856
rect 21474 2 21582 856
rect 21750 2 21766 856
rect 21934 2 21950 856
rect 22118 2 22134 856
rect 22302 2 22410 856
rect 22578 2 22594 856
rect 22762 2 22778 856
rect 22946 2 22962 856
rect 23130 2 23146 856
rect 23314 2 23422 856
rect 23590 2 23606 856
rect 23774 2 23790 856
rect 23958 2 23974 856
rect 24142 2 24158 856
rect 24326 2 24434 856
rect 24602 2 24618 856
rect 24786 2 24802 856
rect 24970 2 24986 856
rect 25154 2 25170 856
rect 25338 2 25446 856
rect 25614 2 25630 856
rect 25798 2 25814 856
rect 25982 2 25998 856
rect 26166 2 26274 856
rect 26442 2 26458 856
rect 26626 2 26642 856
rect 26810 2 26826 856
rect 26994 2 27010 856
rect 27178 2 27286 856
rect 27454 2 27470 856
rect 27638 2 27654 856
rect 27822 2 27838 856
rect 28006 2 28022 856
rect 28190 2 28298 856
rect 28466 2 28482 856
rect 28650 2 28666 856
rect 28834 2 28850 856
rect 29018 2 29034 856
rect 29202 2 29310 856
rect 29478 2 29494 856
rect 29662 2 29678 856
rect 29846 2 29862 856
rect 30030 2 30046 856
rect 30214 2 30322 856
rect 30490 2 30506 856
rect 30674 2 30690 856
rect 30858 2 30874 856
rect 31042 2 31150 856
rect 31318 2 31334 856
rect 31502 2 31518 856
rect 31686 2 31702 856
rect 31870 2 31886 856
rect 32054 2 32162 856
rect 32330 2 32346 856
rect 32514 2 32530 856
rect 32698 2 32714 856
rect 32882 2 32898 856
rect 33066 2 33174 856
rect 33342 2 33358 856
rect 33526 2 33542 856
rect 33710 2 33726 856
rect 33894 2 33910 856
rect 34078 2 34186 856
rect 34354 2 34370 856
rect 34538 2 34554 856
rect 34722 2 34738 856
rect 34906 2 35014 856
rect 35182 2 35198 856
rect 35366 2 35382 856
rect 35550 2 35566 856
rect 35734 2 35750 856
rect 35918 2 36026 856
rect 36194 2 36210 856
rect 36378 2 36394 856
rect 36562 2 36578 856
rect 36746 2 36762 856
rect 36930 2 37038 856
rect 37206 2 37222 856
rect 37390 2 37406 856
rect 37574 2 37590 856
rect 37758 2 37774 856
rect 37942 2 38050 856
rect 38218 2 38234 856
rect 38402 2 38418 856
rect 38586 2 38602 856
rect 38770 2 38786 856
rect 38954 2 39062 856
rect 39230 2 39246 856
rect 39414 2 39430 856
rect 39598 2 39614 856
rect 39782 2 39890 856
rect 40058 2 40074 856
rect 40242 2 40258 856
rect 40426 2 40442 856
rect 40610 2 40626 856
rect 40794 2 40902 856
rect 41070 2 41086 856
rect 41254 2 41270 856
rect 41438 2 41454 856
rect 41622 2 41638 856
rect 41806 2 41914 856
rect 42082 2 42098 856
rect 42266 2 42282 856
rect 42450 2 42466 856
rect 42634 2 42650 856
rect 42818 2 42926 856
rect 43094 2 43110 856
rect 43278 2 43294 856
rect 43462 2 43478 856
rect 43646 2 43754 856
rect 43922 2 43938 856
rect 44106 2 44122 856
rect 44290 2 44306 856
rect 44474 2 44490 856
rect 44658 2 44766 856
rect 44934 2 44950 856
rect 45118 2 45134 856
rect 45302 2 45318 856
rect 45486 2 45502 856
rect 45670 2 45778 856
rect 45946 2 45962 856
rect 46130 2 46146 856
rect 46314 2 46330 856
rect 46498 2 46514 856
rect 46682 2 46790 856
rect 46958 2 46974 856
rect 47142 2 47158 856
rect 47326 2 47342 856
rect 47510 2 47526 856
rect 47694 2 47802 856
rect 47970 2 47986 856
rect 48154 2 48170 856
rect 48338 2 48354 856
rect 48522 2 48630 856
rect 48798 2 48814 856
rect 48982 2 48998 856
rect 49166 2 49182 856
rect 49350 2 49366 856
rect 49534 2 49642 856
rect 49810 2 49826 856
rect 49994 2 50010 856
rect 50178 2 50194 856
rect 50362 2 50378 856
rect 50546 2 50654 856
rect 50822 2 50838 856
rect 51006 2 51022 856
rect 51190 2 51206 856
rect 51374 2 51390 856
rect 51558 2 51666 856
rect 51834 2 51850 856
rect 52018 2 52034 856
rect 52202 2 52218 856
rect 52386 2 52494 856
rect 52662 2 52678 856
rect 52846 2 52862 856
rect 53030 2 53046 856
rect 53214 2 53230 856
rect 53398 2 53506 856
rect 53674 2 53690 856
rect 53858 2 53874 856
rect 54042 2 54058 856
rect 54226 2 54242 856
rect 54410 2 54518 856
rect 54686 2 54702 856
rect 54870 2 54886 856
rect 55054 2 55070 856
rect 55238 2 55254 856
rect 55422 2 55530 856
rect 55698 2 55714 856
rect 55882 2 55898 856
rect 56066 2 56082 856
rect 56250 2 56266 856
rect 56434 2 56542 856
rect 56710 2 56726 856
rect 56894 2 56910 856
rect 57078 2 57094 856
rect 57262 2 57370 856
rect 57538 2 57554 856
rect 57722 2 57738 856
rect 57906 2 57922 856
rect 58090 2 58106 856
rect 58274 2 58382 856
rect 58550 2 58566 856
rect 58734 2 58750 856
rect 58918 2 58934 856
rect 59102 2 59118 856
rect 59286 2 59394 856
rect 59562 2 59578 856
rect 59746 2 59762 856
rect 59930 2 59946 856
rect 60114 2 60130 856
rect 60298 2 60406 856
rect 60574 2 60590 856
rect 60758 2 60774 856
rect 60942 2 60958 856
rect 61126 2 61234 856
rect 61402 2 61418 856
rect 61586 2 61602 856
rect 61770 2 61786 856
rect 61954 2 61970 856
rect 62138 2 62246 856
rect 62414 2 62430 856
rect 62598 2 62614 856
rect 62782 2 62798 856
rect 62966 2 62982 856
rect 63150 2 63258 856
rect 63426 2 63442 856
rect 63610 2 63626 856
rect 63794 2 63810 856
rect 63978 2 63994 856
rect 64162 2 64270 856
rect 64438 2 64454 856
rect 64622 2 64638 856
rect 64806 2 64822 856
rect 64990 2 65006 856
rect 65174 2 65282 856
rect 65450 2 65466 856
rect 65634 2 65650 856
rect 65818 2 65834 856
rect 66002 2 66110 856
rect 66278 2 66294 856
rect 66462 2 66478 856
rect 66646 2 66662 856
rect 66830 2 66846 856
rect 67014 2 67122 856
rect 67290 2 67306 856
rect 67474 2 67490 856
rect 67658 2 67674 856
rect 67842 2 67858 856
rect 68026 2 68134 856
rect 68302 2 68318 856
rect 68486 2 68502 856
rect 68670 2 68686 856
rect 68854 2 68870 856
rect 69038 2 69146 856
rect 69314 2 69330 856
rect 69498 2 69514 856
rect 69682 2 69698 856
rect 69866 2 69974 856
rect 70142 2 70158 856
rect 70326 2 70342 856
rect 70510 2 70526 856
rect 70694 2 70710 856
rect 70878 2 70986 856
rect 71154 2 71170 856
rect 71338 2 71354 856
rect 71522 2 71538 856
rect 71706 2 71722 856
rect 71890 2 71998 856
rect 72166 2 72182 856
rect 72350 2 72366 856
rect 72534 2 72550 856
rect 72718 2 72734 856
rect 72902 2 73010 856
rect 73178 2 73194 856
rect 73362 2 73378 856
rect 73546 2 73562 856
rect 73730 2 73746 856
rect 73914 2 74022 856
rect 74190 2 74206 856
rect 74374 2 74390 856
rect 74558 2 74574 856
rect 74742 2 74850 856
rect 75018 2 75034 856
rect 75202 2 75218 856
rect 75386 2 75402 856
rect 75570 2 75586 856
rect 75754 2 75862 856
rect 76030 2 76046 856
rect 76214 2 76230 856
rect 76398 2 76414 856
rect 76582 2 76598 856
rect 76766 2 76874 856
rect 77042 2 77058 856
rect 77226 2 77242 856
rect 77410 2 77426 856
rect 77594 2 77610 856
rect 77778 2 77886 856
rect 78054 2 78070 856
rect 78238 2 78254 856
rect 78422 2 78438 856
rect 78606 2 78714 856
rect 78882 2 78898 856
rect 79066 2 79082 856
rect 79250 2 79266 856
rect 79434 2 79450 856
rect 79618 2 79726 856
rect 79894 2 79910 856
rect 80078 2 80094 856
rect 80262 2 80278 856
rect 80446 2 80462 856
rect 80630 2 80738 856
rect 80906 2 80922 856
rect 81090 2 81106 856
rect 81274 2 81290 856
rect 81458 2 81474 856
rect 81642 2 81750 856
rect 81918 2 81934 856
rect 82102 2 82118 856
rect 82286 2 82302 856
rect 82470 2 82486 856
rect 82654 2 82762 856
rect 82930 2 82946 856
rect 83114 2 83130 856
rect 83298 2 83314 856
rect 83482 2 83590 856
rect 83758 2 83774 856
rect 83942 2 83958 856
rect 84126 2 84142 856
rect 84310 2 84326 856
rect 84494 2 84602 856
rect 84770 2 84786 856
rect 84954 2 84970 856
rect 85138 2 85154 856
rect 85322 2 85338 856
rect 85506 2 85614 856
rect 85782 2 85798 856
rect 85966 2 85982 856
rect 86150 2 86166 856
rect 86334 2 86350 856
rect 86518 2 86626 856
rect 86794 2 86810 856
rect 86978 2 86994 856
rect 87162 2 87178 856
rect 87346 2 87454 856
rect 87622 2 87638 856
rect 87806 2 87822 856
rect 87990 2 88006 856
rect 88174 2 88190 856
rect 88358 2 88466 856
rect 88634 2 88650 856
rect 88818 2 88834 856
rect 89002 2 89018 856
rect 89186 2 89202 856
rect 89370 2 89478 856
rect 89646 2 89662 856
rect 89830 2 89846 856
rect 90014 2 90030 856
rect 90198 2 90214 856
rect 90382 2 90490 856
rect 90658 2 90674 856
rect 90842 2 90858 856
rect 91026 2 91042 856
rect 91210 2 91226 856
rect 91394 2 91502 856
rect 91670 2 91686 856
rect 91854 2 91870 856
rect 92038 2 92054 856
rect 92222 2 92330 856
rect 92498 2 92514 856
rect 92682 2 92698 856
rect 92866 2 92882 856
rect 93050 2 93066 856
rect 93234 2 93342 856
rect 93510 2 93526 856
rect 93694 2 93710 856
rect 93878 2 93894 856
rect 94062 2 94078 856
rect 94246 2 94354 856
rect 94522 2 94538 856
rect 94706 2 94722 856
rect 94890 2 94906 856
rect 95074 2 95090 856
rect 95258 2 95366 856
rect 95534 2 95550 856
rect 95718 2 95734 856
rect 95902 2 95918 856
rect 96086 2 96194 856
rect 96362 2 96378 856
rect 96546 2 96562 856
rect 96730 2 96746 856
rect 96914 2 96930 856
rect 97098 2 97206 856
rect 97374 2 97390 856
rect 97558 2 97574 856
rect 97742 2 97758 856
rect 97926 2 97942 856
rect 98110 2 98218 856
rect 98386 2 98402 856
rect 98570 2 98586 856
rect 98754 2 98770 856
rect 98938 2 98954 856
rect 99122 2 99230 856
rect 99398 2 99414 856
rect 99582 2 99598 856
rect 99766 2 99782 856
<< metal3 >>
rect 0 20000 800 20120
rect 99200 20000 100000 20120
<< obsm3 >>
rect 800 20200 99200 37569
rect 880 19920 99120 20200
rect 800 171 99200 19920
<< metal4 >>
rect 4208 2128 4528 37584
rect 4868 2176 5188 37536
rect 5528 2176 5848 37536
rect 6188 2176 6508 37536
rect 19568 2128 19888 37584
rect 20228 2176 20548 37536
rect 20888 2176 21208 37536
rect 21548 2176 21868 37536
rect 34928 2128 35248 37584
rect 35588 2176 35908 37536
rect 36248 2176 36568 37536
rect 36908 2176 37228 37536
rect 50288 2128 50608 37584
rect 50948 2176 51268 37536
rect 51608 2176 51928 37536
rect 52268 2176 52588 37536
rect 65648 2128 65968 37584
rect 66308 2176 66628 37536
rect 66968 2176 67288 37536
rect 67628 2176 67948 37536
rect 81008 2128 81328 37584
rect 81668 2176 81988 37536
rect 82328 2176 82648 37536
rect 82988 2176 83308 37536
rect 96368 2128 96688 37584
rect 97028 2176 97348 37536
rect 97688 2176 98008 37536
<< obsm4 >>
rect 38515 11051 38765 26621
<< labels >>
rlabel metal2 s 386 39200 442 40000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 26698 39200 26754 40000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 29274 39200 29330 40000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 31942 39200 31998 40000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 34518 39200 34574 40000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 37186 39200 37242 40000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 39854 39200 39910 40000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 42430 39200 42486 40000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 45098 39200 45154 40000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 47674 39200 47730 40000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 50342 39200 50398 40000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2962 39200 3018 40000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 53010 39200 53066 40000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 55586 39200 55642 40000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 58254 39200 58310 40000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 60830 39200 60886 40000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 63498 39200 63554 40000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 66166 39200 66222 40000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 68742 39200 68798 40000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 71410 39200 71466 40000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 73986 39200 74042 40000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 76654 39200 76710 40000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5630 39200 5686 40000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 79322 39200 79378 40000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 81898 39200 81954 40000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 84566 39200 84622 40000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 87142 39200 87198 40000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 89810 39200 89866 40000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 92478 39200 92534 40000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 95054 39200 95110 40000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 97722 39200 97778 40000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8206 39200 8262 40000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10874 39200 10930 40000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13542 39200 13598 40000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 16118 39200 16174 40000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 18786 39200 18842 40000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 21362 39200 21418 40000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 24030 39200 24086 40000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1214 39200 1270 40000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 27526 39200 27582 40000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 30194 39200 30250 40000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 32770 39200 32826 40000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 35438 39200 35494 40000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 38106 39200 38162 40000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 40682 39200 40738 40000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 43350 39200 43406 40000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 45926 39200 45982 40000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 48594 39200 48650 40000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 51262 39200 51318 40000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3882 39200 3938 40000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 53838 39200 53894 40000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 56506 39200 56562 40000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 59082 39200 59138 40000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 61750 39200 61806 40000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 64418 39200 64474 40000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 66994 39200 67050 40000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 69662 39200 69718 40000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 72238 39200 72294 40000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 74906 39200 74962 40000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 77574 39200 77630 40000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6458 39200 6514 40000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 80150 39200 80206 40000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 82818 39200 82874 40000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 85394 39200 85450 40000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 88062 39200 88118 40000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 90730 39200 90786 40000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 93306 39200 93362 40000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 95974 39200 96030 40000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 98550 39200 98606 40000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9126 39200 9182 40000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 11702 39200 11758 40000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 14370 39200 14426 40000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 17038 39200 17094 40000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 19614 39200 19670 40000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 22282 39200 22338 40000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 24858 39200 24914 40000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2134 39200 2190 40000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 28446 39200 28502 40000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 31022 39200 31078 40000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 33690 39200 33746 40000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 36266 39200 36322 40000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 38934 39200 38990 40000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 41602 39200 41658 40000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 44178 39200 44234 40000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 46846 39200 46902 40000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 49422 39200 49478 40000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 52090 39200 52146 40000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4710 39200 4766 40000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 54758 39200 54814 40000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 57334 39200 57390 40000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 60002 39200 60058 40000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 62578 39200 62634 40000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 65246 39200 65302 40000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 67914 39200 67970 40000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 70490 39200 70546 40000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 73158 39200 73214 40000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 75826 39200 75882 40000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 78402 39200 78458 40000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7378 39200 7434 40000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 81070 39200 81126 40000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 83646 39200 83702 40000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 86314 39200 86370 40000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 88982 39200 89038 40000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 91558 39200 91614 40000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 94226 39200 94282 40000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 96802 39200 96858 40000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 99470 39200 99526 40000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9954 39200 10010 40000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 12622 39200 12678 40000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 15290 39200 15346 40000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 17866 39200 17922 40000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 20534 39200 20590 40000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 23110 39200 23166 40000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 25778 39200 25834 40000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 99200 20000 100000 20120 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 97446 0 97502 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 80334 0 80390 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 user_clock2
port 502 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 503 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 504 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 505 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[0]
port 506 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[10]
port 507 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[11]
port 508 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[12]
port 509 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[13]
port 510 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[14]
port 511 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[15]
port 512 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[16]
port 513 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[17]
port 514 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[18]
port 515 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_adr_i[19]
port 516 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[1]
port 517 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[20]
port 518 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[21]
port 519 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[22]
port 520 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[23]
port 521 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[24]
port 522 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[25]
port 523 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[26]
port 524 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[27]
port 525 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[28]
port 526 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[29]
port 527 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 528 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[30]
port 529 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[31]
port 530 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[3]
port 531 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[4]
port 532 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[5]
port 533 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[6]
port 534 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[7]
port 535 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[8]
port 536 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[9]
port 537 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 538 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 539 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[10]
port 540 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[11]
port 541 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[12]
port 542 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[13]
port 543 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[14]
port 544 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[15]
port 545 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[16]
port 546 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[17]
port 547 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[18]
port 548 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[19]
port 549 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[1]
port 550 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[20]
port 551 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[21]
port 552 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[22]
port 553 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[23]
port 554 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[24]
port 555 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[25]
port 556 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[26]
port 557 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[27]
port 558 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[28]
port 559 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[29]
port 560 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[2]
port 561 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[30]
port 562 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[31]
port 563 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[3]
port 564 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[4]
port 565 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[5]
port 566 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[6]
port 567 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[7]
port 568 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[8]
port 569 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[9]
port 570 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 571 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[10]
port 572 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[11]
port 573 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[12]
port 574 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[13]
port 575 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[14]
port 576 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[15]
port 577 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[16]
port 578 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[17]
port 579 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[18]
port 580 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[19]
port 581 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[1]
port 582 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[20]
port 583 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[21]
port 584 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[22]
port 585 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[23]
port 586 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[24]
port 587 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[25]
port 588 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[26]
port 589 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[27]
port 590 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[28]
port 591 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[29]
port 592 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[2]
port 593 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[30]
port 594 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[31]
port 595 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[3]
port 596 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[4]
port 597 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[5]
port 598 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[6]
port 599 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[7]
port 600 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[8]
port 601 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[9]
port 602 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 603 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 604 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[2]
port 605 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_sel_i[3]
port 606 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 607 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 608 nsew signal input
rlabel metal4 s 96368 2128 96688 37584 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 81008 2128 81328 37584 6 vssd1
port 613 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 97028 2176 97348 37536 6 vccd2
port 616 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 37536 6 vccd2
port 617 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 37536 6 vccd2
port 618 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 37536 6 vccd2
port 619 nsew power bidirectional
rlabel metal4 s 81668 2176 81988 37536 6 vssd2
port 620 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 37536 6 vssd2
port 621 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 37536 6 vssd2
port 622 nsew ground bidirectional
rlabel metal4 s 97688 2176 98008 37536 6 vdda1
port 623 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 37536 6 vdda1
port 624 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 37536 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 37536 6 vdda1
port 626 nsew power bidirectional
rlabel metal4 s 82328 2176 82648 37536 6 vssa1
port 627 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 37536 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 37536 6 vssa1
port 629 nsew ground bidirectional
rlabel metal4 s 67628 2176 67948 37536 6 vdda2
port 630 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 37536 6 vdda2
port 631 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 37536 6 vdda2
port 632 nsew power bidirectional
rlabel metal4 s 82988 2176 83308 37536 6 vssa2
port 633 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 37536 6 vssa2
port 634 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 37536 6 vssa2
port 635 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 100000 40000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 4501790
string GDS_START 312884
<< end >>

