magic
tech sky130A
magscale 1 2
timestamp 1623941680
<< locali >>
rect 5733 37723 5767 38641
rect 17233 37723 17267 38029
rect 26525 37723 26559 38301
rect 31401 37723 31435 39321
rect 36461 38335 36495 38573
rect 40049 37723 40083 39185
rect 41705 37791 41739 38845
rect 42349 37791 42383 38913
rect 47961 37655 47995 38029
rect 48513 37655 48547 38845
rect 52377 37655 52411 39117
rect 54217 38539 54251 39117
rect 56149 37859 56183 38505
rect 57897 37655 57931 38029
rect 63785 37655 63819 39185
rect 74273 37723 74307 38913
rect 80161 37655 80195 39593
rect 84393 37655 84427 38981
rect 87153 37655 87187 38777
rect 89913 37655 89947 39049
rect 40969 37111 41003 37213
rect 46765 36567 46799 36873
rect 12817 36023 12851 36261
rect 50905 36023 50939 36329
rect 85865 34935 85899 35037
rect 31401 32215 31435 32317
rect 32505 32215 32539 32521
rect 42993 32283 43027 32521
rect 19441 31875 19475 31977
rect 88901 31807 88935 31977
rect 94697 31807 94731 31909
rect 59645 31195 59679 31365
rect 85865 30651 85899 30753
rect 79701 29087 79735 29257
rect 37013 28407 37047 28713
rect 19441 26367 19475 26537
rect 35449 26435 35483 26537
rect 20361 24191 20395 24293
rect 36093 24055 36127 24293
rect 65257 24055 65291 24293
rect 25697 23171 25731 23273
rect 84761 21879 84795 21981
rect 43729 21335 43763 21641
rect 58725 21539 58759 21641
rect 60565 21403 60599 21641
rect 38335 20009 38427 20043
rect 38393 19839 38427 20009
rect 38301 19703 38335 19805
rect 72985 18207 73019 18309
rect 61393 17527 61427 17697
rect 31309 15895 31343 16133
rect 58633 13855 58667 13957
rect 85221 12631 85255 12801
rect 58357 12087 58391 12257
rect 14197 11135 14231 11305
rect 69029 11203 69063 11305
rect 95985 11203 96019 11305
rect 26617 11067 26651 11169
rect 66361 10523 66395 10625
rect 29929 10115 29963 10217
rect 57437 9979 57471 10217
rect 57529 10115 57563 10217
rect 50629 9367 50663 9469
rect 61117 8415 61151 8517
rect 67281 8347 67315 8585
rect 27169 7259 27203 7429
rect 7389 5559 7423 5797
rect 6285 5083 6319 5253
rect 6469 5151 6503 5321
rect 38485 5015 38519 5253
rect 79701 5151 79735 5321
rect 54125 4675 54159 4777
rect 54217 4539 54251 4777
rect 40417 3451 40451 3689
rect 22017 2907 22051 3077
rect 69489 2975 69523 3077
rect 76389 2975 76423 3145
rect 80713 2839 80747 3145
rect 90465 2975 90499 3145
rect 78689 2295 78723 2465
rect 31033 51 31067 901
rect 40601 867 40635 1105
rect 40693 935 40727 1105
rect 40785 867 40819 901
rect 40601 833 40819 867
rect 44741 493 45017 527
rect 44741 459 44775 493
rect 46121 119 46155 561
rect 49433 459 49467 1241
rect 51549 1207 51583 2057
rect 58173 1071 58207 1309
<< viali >>
rect 80161 39593 80195 39627
rect 31401 39321 31435 39355
rect 5733 38641 5767 38675
rect 26525 38301 26559 38335
rect 5733 37689 5767 37723
rect 17233 38029 17267 38063
rect 17233 37689 17267 37723
rect 26525 37689 26559 37723
rect 40049 39185 40083 39219
rect 36461 38573 36495 38607
rect 36461 38301 36495 38335
rect 31401 37689 31435 37723
rect 63785 39185 63819 39219
rect 52377 39117 52411 39151
rect 42349 38913 42383 38947
rect 41705 38845 41739 38879
rect 41705 37757 41739 37791
rect 48513 38845 48547 38879
rect 42349 37757 42383 37791
rect 47961 38029 47995 38063
rect 40049 37689 40083 37723
rect 47961 37621 47995 37655
rect 48513 37621 48547 37655
rect 54217 39117 54251 39151
rect 54217 38505 54251 38539
rect 56149 38505 56183 38539
rect 56149 37825 56183 37859
rect 57897 38029 57931 38063
rect 52377 37621 52411 37655
rect 57897 37621 57931 37655
rect 74273 38913 74307 38947
rect 74273 37689 74307 37723
rect 63785 37621 63819 37655
rect 89913 39049 89947 39083
rect 80161 37621 80195 37655
rect 84393 38981 84427 39015
rect 84393 37621 84427 37655
rect 87153 38777 87187 38811
rect 87153 37621 87187 37655
rect 89913 37621 89947 37655
rect 4445 37417 4479 37451
rect 7849 37417 7883 37451
rect 8585 37417 8619 37451
rect 9505 37417 9539 37451
rect 11069 37417 11103 37451
rect 12449 37417 12483 37451
rect 14841 37417 14875 37451
rect 16497 37417 16531 37451
rect 17785 37417 17819 37451
rect 21557 37417 21591 37451
rect 23121 37417 23155 37451
rect 25789 37417 25823 37451
rect 27261 37417 27295 37451
rect 29193 37417 29227 37451
rect 31125 37417 31159 37451
rect 32137 37417 32171 37451
rect 33793 37417 33827 37451
rect 34713 37417 34747 37451
rect 36461 37417 36495 37451
rect 37381 37417 37415 37451
rect 39129 37417 39163 37451
rect 40049 37417 40083 37451
rect 41797 37417 41831 37451
rect 42533 37417 42567 37451
rect 44465 37417 44499 37451
rect 45293 37417 45327 37451
rect 47133 37417 47167 37451
rect 47869 37417 47903 37451
rect 48605 37417 48639 37451
rect 50537 37417 50571 37451
rect 51273 37417 51307 37451
rect 55873 37417 55907 37451
rect 56609 37417 56643 37451
rect 57805 37417 57839 37451
rect 61761 37417 61795 37451
rect 64429 37417 64463 37451
rect 67097 37417 67131 37451
rect 69673 37417 69707 37451
rect 79149 37417 79183 37451
rect 80345 37417 80379 37451
rect 83013 37417 83047 37451
rect 92397 37417 92431 37451
rect 96169 37417 96203 37451
rect 97641 37417 97675 37451
rect 1869 37349 1903 37383
rect 7021 37349 7055 37383
rect 8493 37349 8527 37383
rect 9597 37349 9631 37383
rect 9781 37349 9815 37383
rect 12357 37349 12391 37383
rect 13829 37349 13863 37383
rect 14933 37349 14967 37383
rect 15117 37349 15151 37383
rect 16221 37349 16255 37383
rect 17693 37349 17727 37383
rect 18889 37349 18923 37383
rect 19257 37349 19291 37383
rect 20545 37349 20579 37383
rect 21465 37349 21499 37383
rect 23029 37349 23063 37383
rect 26341 37349 26375 37383
rect 26525 37349 26559 37383
rect 28549 37349 28583 37383
rect 30021 37349 30055 37383
rect 31033 37349 31067 37383
rect 32045 37349 32079 37383
rect 34621 37349 34655 37383
rect 36369 37349 36403 37383
rect 43361 37349 43395 37383
rect 47777 37349 47811 37383
rect 48513 37349 48547 37383
rect 50445 37349 50479 37383
rect 52561 37349 52595 37383
rect 53113 37349 53147 37383
rect 55229 37349 55263 37383
rect 57713 37349 57747 37383
rect 60933 37349 60967 37383
rect 61117 37349 61151 37383
rect 63601 37349 63635 37383
rect 63785 37349 63819 37383
rect 66269 37349 66303 37383
rect 66453 37349 66487 37383
rect 71513 37349 71547 37383
rect 72433 37349 72467 37383
rect 74089 37349 74123 37383
rect 75009 37349 75043 37383
rect 76757 37349 76791 37383
rect 82001 37349 82035 37383
rect 84577 37349 84611 37383
rect 85221 37349 85255 37383
rect 85405 37349 85439 37383
rect 87245 37349 87279 37383
rect 87889 37349 87923 37383
rect 88073 37349 88107 37383
rect 89453 37349 89487 37383
rect 89637 37349 89671 37383
rect 90557 37349 90591 37383
rect 90741 37349 90775 37383
rect 93317 37349 93351 37383
rect 96077 37349 96111 37383
rect 97917 37349 97951 37383
rect 98101 37349 98135 37383
rect 2973 37281 3007 37315
rect 4353 37281 4387 37315
rect 5365 37281 5399 37315
rect 5733 37281 5767 37315
rect 7205 37281 7239 37315
rect 7757 37281 7791 37315
rect 10885 37281 10919 37315
rect 13553 37281 13587 37315
rect 20361 37281 20395 37315
rect 23857 37281 23891 37315
rect 24133 37281 24167 37315
rect 25697 37281 25731 37315
rect 26249 37281 26283 37315
rect 27169 37281 27203 37315
rect 28365 37281 28399 37315
rect 29101 37281 29135 37315
rect 29837 37281 29871 37315
rect 33701 37281 33735 37315
rect 37197 37281 37231 37315
rect 39037 37281 39071 37315
rect 39865 37281 39899 37315
rect 41705 37281 41739 37315
rect 42441 37281 42475 37315
rect 43177 37281 43211 37315
rect 44373 37281 44407 37315
rect 45109 37281 45143 37315
rect 47041 37281 47075 37315
rect 49709 37281 49743 37315
rect 49893 37281 49927 37315
rect 51181 37281 51215 37315
rect 52377 37281 52411 37315
rect 53481 37281 53515 37315
rect 55045 37281 55079 37315
rect 55781 37281 55815 37315
rect 56517 37281 56551 37315
rect 58449 37281 58483 37315
rect 58909 37281 58943 37315
rect 61669 37281 61703 37315
rect 64337 37281 64371 37315
rect 67005 37281 67039 37315
rect 68753 37281 68787 37315
rect 69581 37281 69615 37315
rect 72249 37281 72283 37315
rect 74273 37281 74307 37315
rect 74825 37281 74859 37315
rect 77493 37281 77527 37315
rect 77677 37281 77711 37315
rect 79057 37281 79091 37315
rect 80253 37281 80287 37315
rect 82185 37281 82219 37315
rect 82921 37281 82955 37315
rect 84393 37281 84427 37315
rect 85589 37281 85623 37315
rect 87061 37281 87095 37315
rect 88257 37281 88291 37315
rect 89821 37281 89855 37315
rect 90925 37281 90959 37315
rect 91109 37281 91143 37315
rect 92489 37281 92523 37315
rect 92673 37281 92707 37315
rect 93225 37281 93259 37315
rect 93501 37281 93535 37315
rect 95065 37281 95099 37315
rect 95249 37281 95283 37315
rect 98193 37281 98227 37315
rect 40969 37213 41003 37247
rect 76941 37213 76975 37247
rect 1685 37145 1719 37179
rect 2145 37145 2179 37179
rect 2421 37145 2455 37179
rect 68937 37145 68971 37179
rect 92121 37145 92155 37179
rect 3157 37077 3191 37111
rect 40969 37077 41003 37111
rect 71605 37077 71639 37111
rect 46765 36873 46799 36907
rect 47041 36873 47075 36907
rect 54953 36873 54987 36907
rect 55321 36873 55355 36907
rect 55505 36873 55539 36907
rect 57529 36873 57563 36907
rect 60197 36873 60231 36907
rect 62773 36873 62807 36907
rect 70685 36873 70719 36907
rect 72985 36873 73019 36907
rect 2145 36805 2179 36839
rect 7665 36805 7699 36839
rect 10241 36805 10275 36839
rect 12909 36805 12943 36839
rect 15577 36805 15611 36839
rect 17877 36805 17911 36839
rect 19441 36805 19475 36839
rect 20821 36805 20855 36839
rect 33977 36805 34011 36839
rect 36553 36805 36587 36839
rect 3249 36737 3283 36771
rect 4629 36737 4663 36771
rect 2053 36669 2087 36703
rect 2329 36669 2363 36703
rect 2973 36669 3007 36703
rect 8217 36669 8251 36703
rect 15393 36669 15427 36703
rect 18705 36669 18739 36703
rect 19257 36669 19291 36703
rect 19533 36669 19567 36703
rect 26709 36669 26743 36703
rect 28641 36669 28675 36703
rect 29929 36669 29963 36703
rect 31401 36669 31435 36703
rect 31677 36669 31711 36703
rect 42441 36669 42475 36703
rect 43545 36669 43579 36703
rect 43821 36669 43855 36703
rect 7481 36601 7515 36635
rect 10057 36601 10091 36635
rect 12725 36601 12759 36635
rect 17785 36601 17819 36635
rect 18061 36601 18095 36635
rect 20637 36601 20671 36635
rect 29009 36601 29043 36635
rect 33793 36601 33827 36635
rect 36369 36601 36403 36635
rect 94237 36805 94271 36839
rect 96813 36805 96847 36839
rect 98101 36805 98135 36839
rect 56149 36669 56183 36703
rect 65441 36669 65475 36703
rect 68661 36669 68695 36703
rect 70593 36669 70627 36703
rect 73721 36669 73755 36703
rect 73997 36669 74031 36703
rect 76113 36669 76147 36703
rect 78505 36669 78539 36703
rect 78689 36669 78723 36703
rect 79149 36669 79183 36703
rect 84393 36669 84427 36703
rect 87153 36669 87187 36703
rect 89637 36669 89671 36703
rect 92489 36669 92523 36703
rect 46949 36601 46983 36635
rect 54861 36601 54895 36635
rect 57437 36601 57471 36635
rect 60105 36601 60139 36635
rect 62681 36601 62715 36635
rect 65809 36601 65843 36635
rect 68017 36601 68051 36635
rect 68201 36601 68235 36635
rect 72893 36601 72927 36635
rect 75929 36601 75963 36635
rect 94145 36601 94179 36635
rect 94421 36601 94455 36635
rect 96997 36601 97031 36635
rect 97641 36601 97675 36635
rect 97917 36601 97951 36635
rect 98193 36601 98227 36635
rect 8401 36533 8435 36567
rect 19073 36533 19107 36567
rect 26893 36533 26927 36567
rect 29745 36533 29779 36567
rect 42625 36533 42659 36567
rect 45109 36533 45143 36567
rect 46765 36533 46799 36567
rect 56333 36533 56367 36567
rect 68477 36533 68511 36567
rect 73537 36533 73571 36567
rect 73905 36533 73939 36567
rect 79333 36533 79367 36567
rect 96629 36533 96663 36567
rect 50905 36329 50939 36363
rect 12817 36261 12851 36295
rect 5273 36193 5307 36227
rect 5641 36193 5675 36227
rect 5733 36193 5767 36227
rect 6009 36193 6043 36227
rect 6101 36125 6135 36159
rect 13001 36193 13035 36227
rect 18429 36193 18463 36227
rect 18705 36193 18739 36227
rect 27445 36193 27479 36227
rect 27813 36193 27847 36227
rect 28181 36193 28215 36227
rect 47225 36193 47259 36227
rect 13553 36125 13587 36159
rect 27629 36125 27663 36159
rect 28089 36125 28123 36159
rect 28733 36125 28767 36159
rect 47501 36125 47535 36159
rect 37197 36057 37231 36091
rect 37473 36057 37507 36091
rect 47133 36057 47167 36091
rect 48789 36057 48823 36091
rect 6469 35989 6503 36023
rect 12817 35989 12851 36023
rect 55597 36261 55631 36295
rect 52193 36193 52227 36227
rect 54861 36193 54895 36227
rect 55044 36193 55078 36227
rect 55229 36193 55263 36227
rect 55413 36193 55447 36227
rect 65349 36193 65383 36227
rect 73905 36193 73939 36227
rect 93501 36193 93535 36227
rect 95065 36193 95099 36227
rect 97549 36193 97583 36227
rect 52745 36125 52779 36159
rect 55137 36125 55171 36159
rect 63141 36125 63175 36159
rect 63417 36125 63451 36159
rect 74273 36125 74307 36159
rect 94053 36125 94087 36159
rect 65533 36057 65567 36091
rect 50905 35989 50939 36023
rect 64521 35989 64555 36023
rect 74043 35989 74077 36023
rect 74181 35989 74215 36023
rect 74549 35989 74583 36023
rect 24501 35785 24535 35819
rect 57069 35785 57103 35819
rect 39589 35649 39623 35683
rect 82277 35649 82311 35683
rect 18889 35581 18923 35615
rect 19165 35581 19199 35615
rect 24685 35581 24719 35615
rect 24869 35581 24903 35615
rect 25237 35581 25271 35615
rect 25421 35581 25455 35615
rect 39859 35581 39893 35615
rect 55689 35581 55723 35615
rect 55965 35581 55999 35615
rect 81909 35581 81943 35615
rect 82057 35581 82091 35615
rect 82185 35581 82219 35615
rect 82461 35581 82495 35615
rect 39405 35445 39439 35479
rect 40969 35445 41003 35479
rect 82553 35445 82587 35479
rect 43545 35173 43579 35207
rect 44005 35173 44039 35207
rect 46949 35173 46983 35207
rect 47041 35173 47075 35207
rect 85957 35173 85991 35207
rect 17417 35105 17451 35139
rect 36553 35105 36587 35139
rect 36829 35105 36863 35139
rect 43729 35105 43763 35139
rect 43913 35105 43947 35139
rect 46765 35105 46799 35139
rect 47138 35105 47172 35139
rect 47334 35105 47368 35139
rect 54125 35105 54159 35139
rect 62037 35105 62071 35139
rect 68109 35105 68143 35139
rect 68477 35105 68511 35139
rect 68845 35105 68879 35139
rect 78873 35105 78907 35139
rect 86141 35105 86175 35139
rect 86324 35105 86358 35139
rect 86693 35105 86727 35139
rect 95065 35105 95099 35139
rect 62313 35037 62347 35071
rect 68293 35037 68327 35071
rect 68753 35037 68787 35071
rect 79149 35037 79183 35071
rect 85865 35037 85899 35071
rect 86417 35037 86451 35071
rect 86509 35037 86543 35071
rect 95433 35037 95467 35071
rect 67741 34969 67775 35003
rect 67925 34969 67959 35003
rect 69213 34969 69247 35003
rect 69581 34969 69615 35003
rect 69765 34969 69799 35003
rect 54401 34901 54435 34935
rect 61853 34901 61887 34935
rect 63601 34901 63635 34935
rect 85865 34901 85899 34935
rect 86785 34901 86819 34935
rect 95203 34901 95237 34935
rect 95341 34901 95375 34935
rect 95525 34901 95559 34935
rect 27721 34697 27755 34731
rect 27997 34697 28031 34731
rect 40785 34629 40819 34663
rect 34529 34493 34563 34527
rect 34805 34493 34839 34527
rect 39405 34493 39439 34527
rect 39661 34493 39695 34527
rect 59369 34493 59403 34527
rect 59737 34493 59771 34527
rect 67189 34493 67223 34527
rect 67465 34493 67499 34527
rect 73721 34493 73755 34527
rect 73997 34493 74031 34527
rect 81725 34493 81759 34527
rect 82277 34493 82311 34527
rect 94237 34493 94271 34527
rect 94605 34493 94639 34527
rect 71053 34153 71087 34187
rect 17877 34085 17911 34119
rect 93409 34085 93443 34119
rect 9965 34017 9999 34051
rect 10333 34017 10367 34051
rect 18429 34017 18463 34051
rect 18705 34017 18739 34051
rect 42257 34017 42291 34051
rect 42441 34017 42475 34051
rect 42533 34017 42567 34051
rect 70409 34017 70443 34051
rect 77769 34017 77803 34051
rect 10425 33949 10459 33983
rect 18245 33949 18279 33983
rect 21557 33949 21591 33983
rect 21833 33949 21867 33983
rect 42073 33949 42107 33983
rect 70777 33949 70811 33983
rect 78045 33949 78079 33983
rect 94789 33949 94823 33983
rect 95065 33949 95099 33983
rect 9781 33881 9815 33915
rect 18613 33881 18647 33915
rect 23121 33813 23155 33847
rect 27629 33813 27663 33847
rect 27905 33813 27939 33847
rect 70547 33813 70581 33847
rect 70685 33813 70719 33847
rect 93225 33813 93259 33847
rect 19625 33541 19659 33575
rect 17601 33473 17635 33507
rect 60841 33473 60875 33507
rect 17325 33405 17359 33439
rect 20269 33405 20303 33439
rect 20637 33405 20671 33439
rect 20729 33405 20763 33439
rect 21005 33405 21039 33439
rect 21189 33405 21223 33439
rect 24501 33405 24535 33439
rect 30205 33405 30239 33439
rect 30389 33405 30423 33439
rect 30477 33405 30511 33439
rect 30619 33405 30653 33439
rect 39957 33405 39991 33439
rect 40141 33405 40175 33439
rect 40417 33405 40451 33439
rect 49249 33405 49283 33439
rect 59369 33405 59403 33439
rect 60473 33405 60507 33439
rect 60621 33405 60655 33439
rect 60749 33405 60783 33439
rect 60979 33405 61013 33439
rect 24869 33337 24903 33371
rect 41797 33337 41831 33371
rect 49525 33337 49559 33371
rect 59737 33337 59771 33371
rect 18705 33269 18739 33303
rect 19809 33269 19843 33303
rect 19901 33269 19935 33303
rect 20085 33269 20119 33303
rect 21465 33269 21499 33303
rect 21741 33269 21775 33303
rect 21925 33269 21959 33303
rect 22293 33269 22327 33303
rect 30757 33269 30791 33303
rect 61117 33269 61151 33303
rect 90649 33065 90683 33099
rect 22109 32929 22143 32963
rect 39037 32929 39071 32963
rect 39221 32929 39255 32963
rect 39313 32929 39347 32963
rect 39589 32929 39623 32963
rect 42073 32929 42107 32963
rect 42257 32929 42291 32963
rect 42349 32929 42383 32963
rect 46949 32929 46983 32963
rect 90465 32929 90499 32963
rect 90741 32929 90775 32963
rect 22661 32861 22695 32895
rect 39405 32861 39439 32895
rect 47225 32861 47259 32895
rect 6469 32793 6503 32827
rect 6745 32793 6779 32827
rect 39773 32793 39807 32827
rect 13369 32725 13403 32759
rect 13645 32725 13679 32759
rect 38853 32725 38887 32759
rect 41889 32725 41923 32759
rect 90281 32725 90315 32759
rect 31585 32521 31619 32555
rect 31861 32521 31895 32555
rect 32505 32521 32539 32555
rect 13461 32453 13495 32487
rect 13737 32453 13771 32487
rect 23029 32453 23063 32487
rect 22477 32385 22511 32419
rect 22569 32317 22603 32351
rect 22845 32317 22879 32351
rect 27905 32317 27939 32351
rect 31401 32317 31435 32351
rect 28457 32249 28491 32283
rect 22661 32181 22695 32215
rect 31401 32181 31435 32215
rect 42993 32521 43027 32555
rect 40141 32317 40175 32351
rect 40417 32317 40451 32351
rect 56609 32385 56643 32419
rect 55781 32317 55815 32351
rect 55965 32317 55999 32351
rect 56149 32317 56183 32351
rect 56517 32317 56551 32351
rect 41797 32249 41831 32283
rect 42993 32249 43027 32283
rect 32505 32181 32539 32215
rect 56977 32181 57011 32215
rect 13829 31977 13863 32011
rect 19441 31977 19475 32011
rect 58633 31977 58667 32011
rect 88901 31977 88935 32011
rect 88993 31977 89027 32011
rect 90373 31977 90407 32011
rect 16773 31909 16807 31943
rect 13093 31841 13127 31875
rect 13277 31841 13311 31875
rect 13645 31841 13679 31875
rect 19441 31841 19475 31875
rect 33720 31841 33754 31875
rect 33885 31841 33919 31875
rect 33977 31841 34011 31875
rect 45017 31841 45051 31875
rect 45293 31841 45327 31875
rect 57988 31841 58022 31875
rect 58328 31841 58362 31875
rect 94697 31909 94731 31943
rect 89177 31841 89211 31875
rect 89361 31841 89395 31875
rect 89545 31841 89579 31875
rect 89913 31841 89947 31875
rect 95893 31841 95927 31875
rect 96261 31841 96295 31875
rect 96629 31841 96663 31875
rect 13369 31773 13403 31807
rect 13461 31773 13495 31807
rect 16920 31773 16954 31807
rect 17141 31773 17175 31807
rect 33517 31773 33551 31807
rect 52837 31773 52871 31807
rect 53113 31773 53147 31807
rect 88901 31773 88935 31807
rect 89821 31773 89855 31807
rect 90833 31773 90867 31807
rect 91017 31773 91051 31807
rect 94697 31773 94731 31807
rect 94881 31773 94915 31807
rect 96077 31773 96111 31807
rect 96537 31773 96571 31807
rect 96997 31773 97031 31807
rect 97365 31773 97399 31807
rect 97549 31773 97583 31807
rect 97733 31773 97767 31807
rect 97917 31773 97951 31807
rect 17049 31705 17083 31739
rect 17233 31705 17267 31739
rect 54217 31705 54251 31739
rect 94973 31705 95007 31739
rect 95157 31705 95191 31739
rect 95341 31705 95375 31739
rect 95525 31705 95559 31739
rect 95709 31705 95743 31739
rect 58127 31637 58161 31671
rect 58265 31637 58299 31671
rect 43913 31433 43947 31467
rect 44189 31433 44223 31467
rect 17601 31365 17635 31399
rect 27721 31365 27755 31399
rect 27997 31365 28031 31399
rect 59645 31365 59679 31399
rect 94605 31365 94639 31399
rect 19073 31297 19107 31331
rect 19349 31229 19383 31263
rect 54769 31229 54803 31263
rect 55045 31229 55079 31263
rect 59921 31297 59955 31331
rect 60473 31297 60507 31331
rect 60197 31229 60231 31263
rect 60380 31229 60414 31263
rect 60565 31229 60599 31263
rect 60749 31229 60783 31263
rect 60933 31229 60967 31263
rect 87245 31229 87279 31263
rect 94053 31229 94087 31263
rect 94426 31229 94460 31263
rect 19533 31161 19567 31195
rect 59645 31161 59679 31195
rect 93961 31161 93995 31195
rect 94237 31161 94271 31195
rect 94329 31161 94363 31195
rect 94789 31161 94823 31195
rect 17785 31093 17819 31127
rect 56149 31093 56183 31127
rect 60013 31093 60047 31127
rect 61117 31093 61151 31127
rect 87153 31093 87187 31127
rect 86049 30889 86083 30923
rect 72709 30821 72743 30855
rect 86417 30821 86451 30855
rect 43637 30753 43671 30787
rect 43913 30753 43947 30787
rect 46581 30753 46615 30787
rect 46848 30753 46882 30787
rect 46949 30753 46983 30787
rect 47133 30753 47167 30787
rect 72433 30753 72467 30787
rect 72526 30753 72560 30787
rect 72801 30753 72835 30787
rect 72939 30753 72973 30787
rect 85865 30753 85899 30787
rect 86233 30753 86267 30787
rect 86509 30753 86543 30787
rect 86606 30753 86640 30787
rect 46397 30685 46431 30719
rect 46765 30685 46799 30719
rect 85865 30617 85899 30651
rect 23765 30549 23799 30583
rect 24041 30549 24075 30583
rect 46305 30549 46339 30583
rect 67005 30549 67039 30583
rect 67189 30549 67223 30583
rect 73077 30549 73111 30583
rect 86785 30549 86819 30583
rect 88625 30549 88659 30583
rect 88809 30549 88843 30583
rect 70961 30345 70995 30379
rect 10149 30209 10183 30243
rect 12357 30209 12391 30243
rect 87889 30209 87923 30243
rect 9965 30141 9999 30175
rect 12081 30141 12115 30175
rect 24133 30141 24167 30175
rect 43637 30141 43671 30175
rect 62497 30141 62531 30175
rect 62681 30141 62715 30175
rect 71237 30141 71271 30175
rect 80253 30141 80287 30175
rect 80529 30141 80563 30175
rect 87613 30141 87647 30175
rect 91017 30141 91051 30175
rect 91293 30141 91327 30175
rect 13737 30073 13771 30107
rect 24685 30073 24719 30107
rect 44005 30073 44039 30107
rect 81909 30073 81943 30107
rect 92673 30073 92707 30107
rect 88993 30005 89027 30039
rect 39129 29733 39163 29767
rect 46673 29733 46707 29767
rect 88349 29733 88383 29767
rect 36369 29665 36403 29699
rect 38025 29665 38059 29699
rect 38209 29665 38243 29699
rect 38393 29665 38427 29699
rect 38577 29665 38611 29699
rect 39405 29665 39439 29699
rect 46489 29665 46523 29699
rect 46765 29665 46799 29699
rect 20821 29597 20855 29631
rect 21097 29597 21131 29631
rect 38301 29597 38335 29631
rect 38761 29597 38795 29631
rect 67005 29597 67039 29631
rect 67189 29597 67223 29631
rect 67465 29597 67499 29631
rect 89729 29597 89763 29631
rect 90005 29597 90039 29631
rect 2237 29529 2271 29563
rect 2513 29529 2547 29563
rect 36185 29529 36219 29563
rect 46305 29529 46339 29563
rect 36921 29461 36955 29495
rect 37197 29461 37231 29495
rect 68569 29461 68603 29495
rect 88165 29461 88199 29495
rect 9689 29257 9723 29291
rect 17325 29257 17359 29291
rect 68201 29257 68235 29291
rect 79701 29257 79735 29291
rect 26157 29189 26191 29223
rect 37013 29189 37047 29223
rect 42165 29189 42199 29223
rect 42441 29189 42475 29223
rect 67925 29189 67959 29223
rect 75929 29189 75963 29223
rect 76113 29189 76147 29223
rect 8401 29121 8435 29155
rect 68569 29121 68603 29155
rect 86969 29121 87003 29155
rect 88533 29121 88567 29155
rect 96905 29121 96939 29155
rect 97181 29121 97215 29155
rect 8125 29053 8159 29087
rect 14013 29053 14047 29087
rect 15577 29053 15611 29087
rect 15853 29053 15887 29087
rect 17509 29053 17543 29087
rect 23949 29053 23983 29087
rect 24225 29053 24259 29087
rect 26341 29053 26375 29087
rect 35633 29053 35667 29087
rect 68293 29053 68327 29087
rect 68477 29053 68511 29087
rect 68662 29053 68696 29087
rect 68845 29053 68879 29087
rect 71237 29053 71271 29087
rect 79701 29053 79735 29087
rect 86693 29053 86727 29087
rect 88257 29053 88291 29087
rect 97273 29053 97307 29087
rect 97641 29053 97675 29087
rect 14565 28985 14599 29019
rect 35900 28985 35934 29019
rect 98101 28985 98135 29019
rect 71053 28917 71087 28951
rect 37013 28713 37047 28747
rect 37381 28713 37415 28747
rect 33241 28645 33275 28679
rect 33609 28645 33643 28679
rect 1685 28577 1719 28611
rect 15669 28577 15703 28611
rect 20821 28577 20855 28611
rect 33333 28577 33367 28611
rect 33517 28577 33551 28611
rect 33701 28577 33735 28611
rect 1961 28509 1995 28543
rect 15209 28509 15243 28543
rect 15393 28509 15427 28543
rect 15577 28509 15611 28543
rect 15945 28509 15979 28543
rect 21097 28509 21131 28543
rect 37749 28645 37783 28679
rect 37289 28577 37323 28611
rect 37565 28577 37599 28611
rect 62129 28577 62163 28611
rect 78413 28577 78447 28611
rect 78682 28577 78716 28611
rect 78782 28577 78816 28611
rect 78965 28577 78999 28611
rect 81081 28577 81115 28611
rect 49157 28509 49191 28543
rect 49433 28509 49467 28543
rect 78045 28509 78079 28543
rect 78597 28509 78631 28543
rect 47869 28441 47903 28475
rect 78229 28441 78263 28475
rect 3249 28373 3283 28407
rect 5457 28373 5491 28407
rect 5733 28373 5767 28407
rect 17233 28373 17267 28407
rect 17509 28373 17543 28407
rect 17693 28373 17727 28407
rect 17785 28373 17819 28407
rect 33885 28373 33919 28407
rect 37013 28373 37047 28407
rect 37105 28373 37139 28407
rect 47593 28373 47627 28407
rect 61945 28373 61979 28407
rect 80897 28373 80931 28407
rect 3617 28169 3651 28203
rect 14473 28169 14507 28203
rect 38945 28169 38979 28203
rect 39221 28169 39255 28203
rect 19947 28101 19981 28135
rect 20085 28101 20119 28135
rect 17417 28033 17451 28067
rect 20177 28033 20211 28067
rect 87061 28033 87095 28067
rect 87429 28033 87463 28067
rect 87521 28033 87555 28067
rect 3801 27965 3835 27999
rect 4077 27965 4111 27999
rect 14289 27965 14323 27999
rect 17049 27965 17083 27999
rect 17141 27965 17175 27999
rect 18705 27965 18739 27999
rect 18981 27965 19015 27999
rect 33149 27965 33183 27999
rect 87245 27965 87279 27999
rect 87613 27965 87647 27999
rect 87797 27965 87831 27999
rect 3525 27897 3559 27931
rect 14013 27897 14047 27931
rect 19809 27897 19843 27931
rect 33609 27897 33643 27931
rect 3985 27829 4019 27863
rect 13921 27829 13955 27863
rect 14105 27829 14139 27863
rect 19165 27829 19199 27863
rect 20453 27829 20487 27863
rect 86969 27829 87003 27863
rect 29101 27625 29135 27659
rect 53849 27625 53883 27659
rect 11805 27557 11839 27591
rect 11069 27489 11103 27523
rect 11253 27489 11287 27523
rect 11529 27489 11563 27523
rect 11713 27489 11747 27523
rect 12265 27489 12299 27523
rect 12449 27489 12483 27523
rect 12817 27489 12851 27523
rect 16129 27489 16163 27523
rect 23673 27489 23707 27523
rect 27813 27489 27847 27523
rect 38945 27489 38979 27523
rect 39129 27489 39163 27523
rect 39221 27489 39255 27523
rect 39497 27489 39531 27523
rect 41245 27489 41279 27523
rect 41521 27489 41555 27523
rect 41797 27489 41831 27523
rect 41889 27489 41923 27523
rect 42073 27489 42107 27523
rect 53205 27489 53239 27523
rect 53388 27489 53422 27523
rect 53757 27489 53791 27523
rect 12541 27421 12575 27455
rect 12633 27421 12667 27455
rect 15853 27421 15887 27455
rect 27537 27421 27571 27455
rect 39313 27421 39347 27455
rect 39681 27421 39715 27455
rect 41705 27421 41739 27455
rect 53481 27421 53515 27455
rect 53573 27421 53607 27455
rect 79333 27421 79367 27455
rect 79609 27421 79643 27455
rect 13001 27285 13035 27319
rect 15025 27285 15059 27319
rect 15301 27285 15335 27319
rect 17417 27285 17451 27319
rect 41337 27285 41371 27319
rect 80713 27285 80747 27319
rect 78505 27013 78539 27047
rect 94789 27013 94823 27047
rect 59645 26945 59679 26979
rect 61209 26945 61243 26979
rect 86325 26945 86359 26979
rect 86601 26945 86635 26979
rect 97365 26945 97399 26979
rect 39313 26877 39347 26911
rect 39865 26877 39899 26911
rect 59921 26877 59955 26911
rect 77861 26877 77895 26911
rect 78091 26877 78125 26911
rect 78229 26877 78263 26911
rect 94237 26877 94271 26911
rect 94513 26877 94547 26911
rect 94605 26877 94639 26911
rect 96721 26877 96755 26911
rect 96905 26877 96939 26911
rect 97089 26877 97123 26911
rect 97457 26877 97491 26911
rect 94421 26809 94455 26843
rect 78137 26741 78171 26775
rect 87705 26741 87739 26775
rect 97917 26741 97951 26775
rect 5365 26537 5399 26571
rect 16681 26537 16715 26571
rect 19441 26537 19475 26571
rect 30573 26537 30607 26571
rect 35449 26537 35483 26571
rect 35541 26537 35575 26571
rect 36369 26537 36403 26571
rect 90465 26537 90499 26571
rect 4721 26401 4755 26435
rect 4904 26401 4938 26435
rect 5004 26401 5038 26435
rect 5273 26401 5307 26435
rect 6653 26401 6687 26435
rect 6929 26401 6963 26435
rect 15393 26401 15427 26435
rect 20637 26469 20671 26503
rect 50169 26469 50203 26503
rect 20085 26401 20119 26435
rect 30389 26401 30423 26435
rect 30481 26401 30515 26435
rect 30757 26401 30791 26435
rect 30941 26401 30975 26435
rect 35449 26401 35483 26435
rect 35725 26401 35759 26435
rect 35873 26401 35907 26435
rect 36001 26401 36035 26435
rect 36277 26401 36311 26435
rect 47869 26401 47903 26435
rect 48237 26401 48271 26435
rect 48605 26401 48639 26435
rect 49985 26401 50019 26435
rect 50261 26401 50295 26435
rect 50353 26401 50387 26435
rect 73353 26401 73387 26435
rect 73518 26401 73552 26435
rect 73767 26401 73801 26435
rect 73905 26401 73939 26435
rect 74089 26401 74123 26435
rect 86049 26401 86083 26435
rect 86417 26401 86451 26435
rect 86555 26401 86589 26435
rect 86693 26401 86727 26435
rect 86821 26401 86855 26435
rect 86969 26401 87003 26435
rect 91293 26401 91327 26435
rect 91661 26401 91695 26435
rect 91845 26401 91879 26435
rect 5089 26333 5123 26367
rect 15117 26333 15151 26367
rect 19441 26333 19475 26367
rect 36093 26333 36127 26367
rect 48053 26333 48087 26367
rect 48513 26333 48547 26367
rect 73629 26333 73663 26367
rect 87981 26333 88015 26367
rect 88165 26333 88199 26367
rect 90649 26333 90683 26367
rect 91385 26333 91419 26367
rect 4629 26265 4663 26299
rect 48973 26265 49007 26299
rect 86233 26265 86267 26299
rect 50537 26197 50571 26231
rect 68753 25925 68787 25959
rect 19073 25789 19107 25823
rect 22937 25789 22971 25823
rect 39228 25789 39262 25823
rect 39405 25789 39439 25823
rect 39589 25789 39623 25823
rect 39865 25789 39899 25823
rect 39957 25789 39991 25823
rect 61669 25789 61703 25823
rect 66361 25789 66395 25823
rect 67189 25789 67223 25823
rect 67465 25789 67499 25823
rect 80437 25789 80471 25823
rect 19340 25721 19374 25755
rect 20453 25653 20487 25687
rect 40417 25653 40451 25687
rect 21649 25449 21683 25483
rect 43545 25449 43579 25483
rect 52377 25449 52411 25483
rect 42625 25381 42659 25415
rect 21557 25313 21591 25347
rect 21833 25313 21867 25347
rect 41245 25313 41279 25347
rect 43637 25313 43671 25347
rect 43913 25313 43947 25347
rect 44041 25313 44075 25347
rect 44189 25313 44223 25347
rect 51641 25313 51675 25347
rect 51825 25313 51859 25347
rect 52193 25313 52227 25347
rect 53021 25313 53055 25347
rect 53205 25313 53239 25347
rect 53297 25313 53331 25347
rect 73629 25313 73663 25347
rect 90649 25313 90683 25347
rect 91017 25313 91051 25347
rect 91385 25313 91419 25347
rect 40969 25245 41003 25279
rect 43821 25245 43855 25279
rect 51917 25245 51951 25279
rect 52009 25245 52043 25279
rect 74365 25245 74399 25279
rect 90833 25245 90867 25279
rect 91293 25245 91327 25279
rect 21465 25109 21499 25143
rect 22017 25109 22051 25143
rect 27721 25109 27755 25143
rect 43361 25109 43395 25143
rect 52837 25109 52871 25143
rect 90097 25109 90131 25143
rect 90281 25109 90315 25143
rect 90465 25109 90499 25143
rect 91845 25109 91879 25143
rect 92121 25109 92155 25143
rect 92305 25109 92339 25143
rect 92489 25109 92523 25143
rect 2237 24837 2271 24871
rect 71421 24837 71455 24871
rect 1869 24769 1903 24803
rect 3433 24769 3467 24803
rect 1501 24701 1535 24735
rect 1684 24701 1718 24735
rect 1777 24701 1811 24735
rect 2053 24701 2087 24735
rect 2421 24701 2455 24735
rect 3341 24701 3375 24735
rect 3709 24701 3743 24735
rect 3893 24701 3927 24735
rect 12173 24701 12207 24735
rect 12449 24701 12483 24735
rect 30665 24701 30699 24735
rect 43545 24701 43579 24735
rect 43821 24701 43855 24735
rect 45201 24701 45235 24735
rect 50905 24701 50939 24735
rect 51181 24701 51215 24735
rect 78045 24701 78079 24735
rect 78321 24701 78355 24735
rect 29837 24633 29871 24667
rect 76665 24633 76699 24667
rect 78413 24633 78447 24667
rect 78597 24633 78631 24667
rect 78781 24633 78815 24667
rect 2605 24565 2639 24599
rect 2973 24565 3007 24599
rect 52469 24565 52503 24599
rect 76113 24565 76147 24599
rect 76297 24565 76331 24599
rect 76481 24565 76515 24599
rect 17601 24361 17635 24395
rect 21833 24361 21867 24395
rect 20361 24293 20395 24327
rect 3249 24225 3283 24259
rect 16773 24225 16807 24259
rect 16865 24225 16899 24259
rect 17141 24225 17175 24259
rect 17325 24225 17359 24259
rect 17509 24225 17543 24259
rect 36093 24293 36127 24327
rect 46397 24293 46431 24327
rect 46489 24293 46523 24327
rect 65257 24293 65291 24327
rect 75837 24293 75871 24327
rect 22569 24225 22603 24259
rect 16037 24157 16071 24191
rect 20361 24157 20395 24191
rect 20453 24157 20487 24191
rect 20729 24157 20763 24191
rect 23305 24157 23339 24191
rect 16405 24089 16439 24123
rect 40969 24225 41003 24259
rect 46213 24225 46247 24259
rect 46581 24225 46615 24259
rect 41153 24089 41187 24123
rect 46765 24089 46799 24123
rect 75377 24225 75411 24259
rect 75561 24225 75595 24259
rect 75745 24225 75779 24259
rect 75929 24225 75963 24259
rect 83013 24225 83047 24259
rect 83196 24225 83230 24259
rect 83565 24225 83599 24259
rect 76297 24157 76331 24191
rect 83289 24157 83323 24191
rect 83381 24157 83415 24191
rect 3249 24021 3283 24055
rect 36093 24021 36127 24055
rect 36369 24021 36403 24055
rect 65257 24021 65291 24055
rect 65533 24021 65567 24055
rect 76113 24021 76147 24055
rect 83657 24021 83691 24055
rect 76941 23817 76975 23851
rect 80069 23817 80103 23851
rect 80253 23817 80287 23851
rect 25237 23749 25271 23783
rect 50169 23749 50203 23783
rect 66361 23749 66395 23783
rect 69949 23749 69983 23783
rect 72157 23749 72191 23783
rect 95341 23749 95375 23783
rect 95617 23749 95651 23783
rect 95801 23749 95835 23783
rect 25329 23681 25363 23715
rect 48789 23681 48823 23715
rect 49065 23681 49099 23715
rect 96261 23681 96295 23715
rect 97733 23681 97767 23715
rect 97917 23681 97951 23715
rect 98101 23681 98135 23715
rect 4813 23613 4847 23647
rect 14473 23613 14507 23647
rect 25108 23613 25142 23647
rect 66085 23613 66119 23647
rect 72249 23613 72283 23647
rect 72525 23613 72559 23647
rect 75009 23613 75043 23647
rect 76757 23613 76791 23647
rect 77125 23613 77159 23647
rect 77309 23613 77343 23647
rect 77401 23613 77435 23647
rect 79149 23613 79183 23647
rect 95985 23613 96019 23647
rect 4537 23545 4571 23579
rect 24961 23545 24995 23579
rect 65809 23545 65843 23579
rect 75254 23545 75288 23579
rect 25605 23477 25639 23511
rect 65533 23477 65567 23511
rect 65901 23477 65935 23511
rect 76389 23477 76423 23511
rect 97365 23477 97399 23511
rect 25697 23273 25731 23307
rect 26525 23273 26559 23307
rect 48513 23273 48547 23307
rect 73261 23273 73295 23307
rect 11161 23205 11195 23239
rect 61853 23205 61887 23239
rect 72433 23205 72467 23239
rect 14749 23137 14783 23171
rect 14933 23137 14967 23171
rect 15025 23137 15059 23171
rect 15117 23137 15151 23171
rect 25697 23137 25731 23171
rect 25789 23137 25823 23171
rect 25973 23137 26007 23171
rect 26203 23137 26237 23171
rect 26341 23137 26375 23171
rect 47501 23137 47535 23171
rect 48421 23137 48455 23171
rect 61945 23137 61979 23171
rect 62129 23137 62163 23171
rect 62497 23137 62531 23171
rect 70133 23137 70167 23171
rect 70685 23137 70719 23171
rect 72617 23137 72651 23171
rect 72765 23137 72799 23171
rect 72985 23137 73019 23171
rect 73169 23137 73203 23171
rect 9505 23069 9539 23103
rect 9781 23069 9815 23103
rect 26065 23069 26099 23103
rect 47685 23069 47719 23103
rect 48053 23069 48087 23103
rect 62221 23069 62255 23103
rect 62313 23069 62347 23103
rect 67465 23069 67499 23103
rect 67741 23069 67775 23103
rect 72893 23069 72927 23103
rect 15301 23001 15335 23035
rect 47317 23001 47351 23035
rect 48697 23001 48731 23035
rect 48145 22933 48179 22967
rect 48283 22933 48317 22967
rect 62681 22933 62715 22967
rect 69029 22933 69063 22967
rect 73445 22933 73479 22967
rect 14657 22729 14691 22763
rect 14933 22729 14967 22763
rect 65901 22661 65935 22695
rect 33701 22593 33735 22627
rect 64981 22593 65015 22627
rect 65533 22593 65567 22627
rect 33517 22525 33551 22559
rect 33977 22525 34011 22559
rect 65165 22525 65199 22559
rect 65349 22525 65383 22559
rect 65441 22525 65475 22559
rect 65717 22525 65751 22559
rect 75009 22525 75043 22559
rect 76113 22525 76147 22559
rect 75285 22457 75319 22491
rect 35265 22389 35299 22423
rect 38389 22117 38423 22151
rect 52469 22117 52503 22151
rect 9873 22049 9907 22083
rect 38117 22049 38151 22083
rect 38301 22049 38335 22083
rect 38485 22049 38519 22083
rect 43545 22049 43579 22083
rect 43637 22049 43671 22083
rect 43821 22049 43855 22083
rect 52193 22049 52227 22083
rect 75377 22049 75411 22083
rect 85037 22049 85071 22083
rect 85405 22049 85439 22083
rect 85773 22049 85807 22083
rect 10425 21981 10459 22015
rect 44005 21981 44039 22015
rect 84761 21981 84795 22015
rect 85313 21981 85347 22015
rect 85681 21981 85715 22015
rect 43453 21913 43487 21947
rect 38025 21845 38059 21879
rect 38669 21845 38703 21879
rect 58633 21845 58667 21879
rect 84761 21845 84795 21879
rect 84853 21845 84887 21879
rect 86233 21845 86267 21879
rect 43729 21641 43763 21675
rect 32873 21573 32907 21607
rect 33241 21573 33275 21607
rect 12449 21505 12483 21539
rect 12081 21437 12115 21471
rect 12265 21437 12299 21471
rect 12357 21437 12391 21471
rect 12633 21437 12667 21471
rect 12817 21437 12851 21471
rect 25881 21437 25915 21471
rect 26029 21437 26063 21471
rect 26157 21437 26191 21471
rect 26249 21437 26283 21471
rect 26433 21437 26467 21471
rect 39681 21437 39715 21471
rect 41153 21437 41187 21471
rect 41429 21437 41463 21471
rect 39773 21369 39807 21403
rect 58725 21641 58759 21675
rect 44005 21573 44039 21607
rect 52285 21505 52319 21539
rect 54033 21505 54067 21539
rect 58725 21505 58759 21539
rect 60565 21641 60599 21675
rect 51917 21437 51951 21471
rect 52101 21437 52135 21471
rect 52193 21437 52227 21471
rect 52469 21437 52503 21471
rect 54309 21437 54343 21471
rect 55689 21437 55723 21471
rect 65165 21505 65199 21539
rect 60657 21437 60691 21471
rect 60841 21437 60875 21471
rect 60936 21437 60970 21471
rect 61025 21437 61059 21471
rect 61192 21437 61226 21471
rect 82553 21437 82587 21471
rect 60565 21369 60599 21403
rect 26525 21301 26559 21335
rect 43729 21301 43763 21335
rect 52653 21301 52687 21335
rect 61393 21301 61427 21335
rect 1869 21097 1903 21131
rect 2697 21097 2731 21131
rect 17509 21097 17543 21131
rect 1685 21029 1719 21063
rect 4997 21029 5031 21063
rect 6193 21029 6227 21063
rect 63417 21029 63451 21063
rect 81725 21029 81759 21063
rect 95341 21029 95375 21063
rect 1501 20961 1535 20995
rect 1961 20961 1995 20995
rect 2237 20961 2271 20995
rect 2365 20961 2399 20995
rect 2513 20961 2547 20995
rect 5457 20961 5491 20995
rect 5861 20961 5895 20995
rect 6009 20961 6043 20995
rect 15945 20961 15979 20995
rect 18613 20961 18647 20995
rect 44281 20961 44315 20995
rect 63233 20961 63267 20995
rect 63509 20961 63543 20995
rect 67373 20961 67407 20995
rect 80345 20961 80379 20995
rect 93961 20961 93995 20995
rect 95433 20961 95467 20995
rect 95617 20961 95651 20995
rect 95801 20961 95835 20995
rect 95985 20961 96019 20995
rect 96169 20961 96203 20995
rect 2145 20893 2179 20927
rect 5181 20893 5215 20927
rect 5641 20893 5675 20927
rect 5733 20893 5767 20927
rect 16221 20893 16255 20927
rect 18797 20893 18831 20927
rect 44557 20893 44591 20927
rect 80069 20893 80103 20927
rect 93685 20893 93719 20927
rect 5365 20757 5399 20791
rect 63049 20757 63083 20791
rect 64153 20757 64187 20791
rect 92765 20757 92799 20791
rect 93133 20757 93167 20791
rect 93317 20757 93351 20791
rect 93501 20757 93535 20791
rect 22753 20553 22787 20587
rect 94237 20553 94271 20587
rect 70593 20485 70627 20519
rect 71421 20485 71455 20519
rect 71789 20485 71823 20519
rect 70225 20417 70259 20451
rect 72709 20417 72743 20451
rect 97457 20417 97491 20451
rect 15669 20349 15703 20383
rect 34253 20349 34287 20383
rect 52009 20349 52043 20383
rect 64521 20349 64555 20383
rect 69857 20349 69891 20383
rect 70005 20349 70039 20383
rect 70133 20349 70167 20383
rect 70409 20349 70443 20383
rect 71973 20349 72007 20383
rect 72157 20349 72191 20383
rect 72525 20349 72559 20383
rect 72893 20349 72927 20383
rect 81633 20349 81667 20383
rect 81817 20349 81851 20383
rect 81955 20349 81989 20383
rect 82093 20349 82127 20383
rect 82186 20349 82220 20383
rect 82369 20349 82403 20383
rect 93501 20349 93535 20383
rect 93685 20349 93719 20383
rect 93786 20349 93820 20383
rect 93915 20349 93949 20383
rect 94053 20349 94087 20383
rect 97089 20349 97123 20383
rect 52285 20281 52319 20315
rect 64788 20281 64822 20315
rect 65901 20213 65935 20247
rect 72985 20213 73019 20247
rect 81449 20213 81483 20247
rect 38301 20009 38335 20043
rect 38485 20009 38519 20043
rect 97641 20009 97675 20043
rect 1409 19873 1443 19907
rect 28825 19873 28859 19907
rect 33425 19873 33459 19907
rect 54861 19941 54895 19975
rect 54953 19941 54987 19975
rect 97365 19941 97399 19975
rect 97549 19941 97583 19975
rect 38669 19873 38703 19907
rect 48789 19873 48823 19907
rect 54677 19873 54711 19907
rect 55045 19873 55079 19907
rect 59461 19873 59495 19907
rect 64613 19873 64647 19907
rect 73997 19873 74031 19907
rect 75653 19873 75687 19907
rect 75837 19873 75871 19907
rect 29101 19805 29135 19839
rect 38301 19805 38335 19839
rect 38393 19805 38427 19839
rect 50537 19805 50571 19839
rect 74733 19805 74767 19839
rect 76205 19805 76239 19839
rect 55229 19737 55263 19771
rect 59277 19737 59311 19771
rect 33241 19669 33275 19703
rect 38301 19669 38335 19703
rect 64429 19669 64463 19703
rect 50077 19465 50111 19499
rect 49341 19397 49375 19431
rect 44373 19329 44407 19363
rect 50537 19329 50571 19363
rect 61025 19329 61059 19363
rect 98101 19329 98135 19363
rect 35909 19261 35943 19295
rect 36092 19261 36126 19295
rect 36185 19261 36219 19295
rect 36323 19261 36357 19295
rect 36461 19261 36495 19295
rect 45845 19261 45879 19295
rect 46121 19261 46155 19295
rect 50261 19261 50295 19295
rect 50445 19261 50479 19295
rect 50629 19261 50663 19295
rect 50813 19261 50847 19295
rect 52377 19261 52411 19295
rect 60473 19261 60507 19295
rect 52653 19193 52687 19227
rect 36553 19125 36587 19159
rect 44741 19125 44775 19159
rect 50997 19125 51031 19159
rect 59553 18921 59587 18955
rect 7021 18853 7055 18887
rect 7205 18853 7239 18887
rect 71053 18853 71087 18887
rect 4997 18785 5031 18819
rect 5181 18785 5215 18819
rect 6653 18785 6687 18819
rect 6929 18785 6963 18819
rect 15577 18785 15611 18819
rect 52561 18785 52595 18819
rect 52965 18785 52999 18819
rect 53113 18785 53147 18819
rect 59553 18785 59587 18819
rect 70777 18785 70811 18819
rect 15853 18717 15887 18751
rect 52745 18717 52779 18751
rect 52837 18717 52871 18751
rect 52377 18649 52411 18683
rect 5365 18581 5399 18615
rect 16957 18581 16991 18615
rect 52285 18581 52319 18615
rect 74641 18581 74675 18615
rect 3157 18377 3191 18411
rect 3341 18377 3375 18411
rect 3525 18377 3559 18411
rect 3801 18377 3835 18411
rect 5181 18377 5215 18411
rect 5365 18377 5399 18411
rect 5549 18377 5583 18411
rect 35173 18309 35207 18343
rect 72985 18309 73019 18343
rect 73215 18309 73249 18343
rect 73353 18309 73387 18343
rect 4353 18241 4387 18275
rect 34069 18241 34103 18275
rect 39596 18241 39630 18275
rect 73445 18241 73479 18275
rect 73721 18241 73755 18275
rect 89545 18241 89579 18275
rect 92949 18241 92983 18275
rect 4261 18173 4295 18207
rect 4629 18173 4663 18207
rect 4813 18173 4847 18207
rect 4997 18173 5031 18207
rect 33793 18173 33827 18207
rect 39313 18173 39347 18207
rect 39496 18173 39530 18207
rect 39681 18173 39715 18207
rect 39865 18173 39899 18207
rect 62681 18173 62715 18207
rect 69765 18173 69799 18207
rect 70041 18173 70075 18207
rect 72985 18173 73019 18207
rect 75929 18173 75963 18207
rect 89269 18173 89303 18207
rect 92673 18173 92707 18207
rect 39129 18105 39163 18139
rect 63233 18105 63267 18139
rect 71421 18105 71455 18139
rect 73077 18105 73111 18139
rect 91293 18105 91327 18139
rect 39957 18037 39991 18071
rect 91201 18037 91235 18071
rect 2513 17697 2547 17731
rect 2881 17697 2915 17731
rect 3065 17697 3099 17731
rect 61393 17697 61427 17731
rect 2145 17629 2179 17663
rect 2421 17629 2455 17663
rect 28365 17629 28399 17663
rect 59185 17629 59219 17663
rect 59461 17629 59495 17663
rect 57897 17561 57931 17595
rect 57621 17493 57655 17527
rect 61393 17493 61427 17527
rect 77953 17289 77987 17323
rect 78689 17289 78723 17323
rect 93961 17289 93995 17323
rect 94421 17289 94455 17323
rect 94053 17221 94087 17255
rect 94605 17221 94639 17255
rect 34529 17153 34563 17187
rect 94145 17153 94179 17187
rect 13553 17085 13587 17119
rect 13829 17085 13863 17119
rect 34345 17085 34379 17119
rect 34713 17085 34747 17119
rect 35081 17085 35115 17119
rect 35265 17085 35299 17119
rect 35633 17085 35667 17119
rect 77677 17085 77711 17119
rect 78045 17085 78079 17119
rect 78229 17085 78263 17119
rect 78321 17085 78355 17119
rect 78449 17085 78483 17119
rect 78597 17085 78631 17119
rect 87521 17085 87555 17119
rect 93593 17085 93627 17119
rect 93225 17017 93259 17051
rect 34253 16949 34287 16983
rect 93409 16949 93443 16983
rect 67925 16745 67959 16779
rect 27537 16677 27571 16711
rect 28825 16677 28859 16711
rect 57161 16677 57195 16711
rect 84485 16677 84519 16711
rect 25881 16609 25915 16643
rect 27997 16609 28031 16643
rect 41061 16609 41095 16643
rect 41429 16609 41463 16643
rect 56793 16609 56827 16643
rect 67741 16609 67775 16643
rect 69038 16609 69072 16643
rect 69305 16609 69339 16643
rect 84117 16609 84151 16643
rect 26151 16541 26185 16575
rect 6745 16201 6779 16235
rect 7021 16201 7055 16235
rect 25881 16201 25915 16235
rect 31401 16201 31435 16235
rect 31585 16201 31619 16235
rect 76941 16201 76975 16235
rect 31309 16133 31343 16167
rect 34069 16133 34103 16167
rect 17785 16065 17819 16099
rect 17536 15997 17570 16031
rect 17693 15997 17727 16031
rect 17878 15997 17912 16031
rect 18061 15997 18095 16031
rect 17325 15929 17359 15963
rect 72525 16065 72559 16099
rect 75561 16065 75595 16099
rect 31723 15997 31757 16031
rect 31861 15997 31895 16031
rect 32137 15997 32171 16031
rect 56333 15997 56367 16031
rect 66177 15997 66211 16031
rect 70869 15997 70903 16031
rect 71145 15997 71179 16031
rect 75837 15997 75871 16031
rect 31953 15929 31987 15963
rect 17233 15861 17267 15895
rect 31309 15861 31343 15895
rect 40969 15589 41003 15623
rect 41429 15589 41463 15623
rect 49065 15589 49099 15623
rect 54677 15589 54711 15623
rect 69673 15589 69707 15623
rect 17049 15521 17083 15555
rect 17325 15521 17359 15555
rect 17601 15521 17635 15555
rect 17693 15521 17727 15555
rect 17877 15521 17911 15555
rect 18429 15521 18463 15555
rect 18797 15521 18831 15555
rect 41337 15521 41371 15555
rect 41521 15521 41555 15555
rect 41705 15521 41739 15555
rect 48789 15521 48823 15555
rect 48882 15521 48916 15555
rect 49157 15521 49191 15555
rect 49295 15521 49329 15555
rect 54493 15521 54527 15555
rect 54769 15521 54803 15555
rect 54861 15521 54895 15555
rect 58541 15521 58575 15555
rect 69121 15521 69155 15555
rect 83933 15521 83967 15555
rect 84117 15521 84151 15555
rect 84301 15521 84335 15555
rect 89729 15521 89763 15555
rect 90051 15521 90085 15555
rect 90189 15521 90223 15555
rect 17509 15453 17543 15487
rect 59001 15453 59035 15487
rect 89269 15453 89303 15487
rect 83749 15385 83783 15419
rect 17141 15317 17175 15351
rect 41153 15317 41187 15351
rect 41889 15317 41923 15351
rect 49433 15317 49467 15351
rect 54033 15317 54067 15351
rect 54309 15317 54343 15351
rect 55045 15317 55079 15351
rect 12265 15113 12299 15147
rect 19441 15113 19475 15147
rect 52561 15113 52595 15147
rect 92213 15113 92247 15147
rect 93961 15113 93995 15147
rect 69949 15045 69983 15079
rect 19901 14977 19935 15011
rect 35909 14977 35943 15011
rect 9413 14909 9447 14943
rect 9689 14909 9723 14943
rect 18429 14909 18463 14943
rect 19533 14909 19567 14943
rect 19717 14909 19751 14943
rect 19809 14909 19843 14943
rect 20085 14909 20119 14943
rect 33149 14909 33183 14943
rect 34069 14909 34103 14943
rect 35541 14909 35575 14943
rect 35724 14909 35758 14943
rect 35817 14909 35851 14943
rect 36093 14909 36127 14943
rect 60473 14909 60507 14943
rect 70041 14909 70075 14943
rect 70317 14909 70351 14943
rect 72801 14909 72835 14943
rect 92397 14909 92431 14943
rect 92673 14909 92707 14943
rect 18981 14841 19015 14875
rect 20269 14841 20303 14875
rect 61025 14841 61059 14875
rect 71697 14841 71731 14875
rect 73353 14841 73387 14875
rect 36185 14773 36219 14807
rect 31861 14569 31895 14603
rect 41061 14569 41095 14603
rect 60289 14569 60323 14603
rect 70409 14501 70443 14535
rect 5089 14433 5123 14467
rect 10241 14433 10275 14467
rect 10425 14433 10459 14467
rect 10609 14433 10643 14467
rect 10793 14433 10827 14467
rect 30481 14433 30515 14467
rect 40785 14433 40819 14467
rect 42174 14433 42208 14467
rect 59645 14433 59679 14467
rect 59793 14433 59827 14467
rect 60013 14433 60047 14467
rect 60197 14433 60231 14467
rect 70225 14433 70259 14467
rect 70501 14433 70535 14467
rect 70645 14433 70679 14467
rect 96997 14433 97031 14467
rect 97181 14433 97215 14467
rect 97549 14433 97583 14467
rect 5365 14365 5399 14399
rect 10885 14365 10919 14399
rect 11161 14365 11195 14399
rect 30757 14365 30791 14399
rect 42441 14365 42475 14399
rect 59921 14365 59955 14399
rect 96721 14365 96755 14399
rect 97457 14365 97491 14399
rect 12449 14297 12483 14331
rect 6653 14229 6687 14263
rect 12725 14229 12759 14263
rect 12909 14229 12943 14263
rect 13093 14229 13127 14263
rect 70777 14229 70811 14263
rect 40877 14025 40911 14059
rect 44097 14025 44131 14059
rect 73905 14025 73939 14059
rect 97825 14025 97859 14059
rect 58633 13957 58667 13991
rect 96445 13957 96479 13991
rect 10333 13889 10367 13923
rect 56517 13889 56551 13923
rect 65993 13889 66027 13923
rect 73353 13889 73387 13923
rect 96813 13889 96847 13923
rect 97273 13889 97307 13923
rect 9781 13821 9815 13855
rect 43545 13821 43579 13855
rect 43729 13821 43763 13855
rect 43965 13821 43999 13855
rect 49525 13821 49559 13855
rect 55413 13821 55447 13855
rect 55965 13821 55999 13855
rect 56241 13821 56275 13855
rect 58633 13821 58667 13855
rect 66177 13821 66211 13855
rect 66453 13821 66487 13855
rect 69949 13821 69983 13855
rect 72709 13821 72743 13855
rect 72893 13821 72927 13855
rect 73077 13821 73111 13855
rect 73445 13821 73479 13855
rect 82001 13821 82035 13855
rect 82829 13821 82863 13855
rect 96629 13821 96663 13855
rect 96997 13821 97031 13855
rect 97365 13821 97399 13855
rect 43821 13753 43855 13787
rect 66637 13753 66671 13787
rect 66269 13685 66303 13719
rect 27169 13413 27203 13447
rect 26893 13345 26927 13379
rect 27077 13345 27111 13379
rect 27261 13345 27295 13379
rect 72801 13345 72835 13379
rect 73169 13345 73203 13379
rect 83059 13345 83093 13379
rect 83289 13277 83323 13311
rect 95249 13277 95283 13311
rect 27445 13141 27479 13175
rect 52101 13141 52135 13175
rect 81633 13141 81667 13175
rect 22385 12937 22419 12971
rect 7941 12801 7975 12835
rect 12633 12801 12667 12835
rect 13093 12801 13127 12835
rect 43453 12801 43487 12835
rect 43821 12801 43855 12835
rect 71329 12801 71363 12835
rect 85221 12801 85255 12835
rect 85773 12801 85807 12835
rect 86325 12801 86359 12835
rect 7665 12733 7699 12767
rect 12909 12733 12943 12767
rect 13185 12733 13219 12767
rect 13277 12733 13311 12767
rect 13461 12733 13495 12767
rect 22753 12733 22787 12767
rect 23029 12733 23063 12767
rect 43545 12733 43579 12767
rect 66453 12733 66487 12767
rect 71605 12733 71639 12767
rect 75653 12733 75687 12767
rect 9321 12665 9355 12699
rect 66821 12665 66855 12699
rect 85497 12733 85531 12767
rect 85681 12733 85715 12767
rect 85865 12733 85899 12767
rect 86049 12733 86083 12767
rect 96537 12733 96571 12767
rect 86233 12665 86267 12699
rect 12725 12597 12759 12631
rect 44925 12597 44959 12631
rect 72709 12597 72743 12631
rect 75469 12597 75503 12631
rect 85221 12597 85255 12631
rect 85405 12597 85439 12631
rect 59645 12393 59679 12427
rect 65809 12393 65843 12427
rect 42717 12325 42751 12359
rect 42809 12325 42843 12359
rect 10609 12257 10643 12291
rect 10885 12257 10919 12291
rect 17693 12257 17727 12291
rect 42533 12257 42567 12291
rect 42901 12257 42935 12291
rect 46489 12257 46523 12291
rect 58357 12257 58391 12291
rect 58449 12257 58483 12291
rect 58817 12257 58851 12291
rect 59093 12257 59127 12291
rect 59185 12257 59219 12291
rect 62221 12257 62255 12291
rect 65993 12257 66027 12291
rect 72617 12257 72651 12291
rect 18245 12189 18279 12223
rect 46213 12189 46247 12223
rect 47593 12189 47627 12223
rect 58909 12189 58943 12223
rect 62497 12189 62531 12223
rect 4445 12053 4479 12087
rect 43085 12053 43119 12087
rect 57713 12053 57747 12087
rect 58357 12053 58391 12087
rect 65349 12053 65383 12087
rect 67373 12053 67407 12087
rect 97641 11849 97675 11883
rect 10333 11781 10367 11815
rect 85497 11781 85531 11815
rect 91017 11781 91051 11815
rect 7113 11713 7147 11747
rect 13001 11713 13035 11747
rect 28641 11713 28675 11747
rect 75561 11713 75595 11747
rect 6837 11645 6871 11679
rect 12817 11645 12851 11679
rect 15209 11645 15243 11679
rect 27813 11645 27847 11679
rect 35081 11645 35115 11679
rect 38209 11645 38243 11679
rect 38393 11645 38427 11679
rect 38576 11645 38610 11679
rect 38669 11645 38703 11679
rect 38807 11645 38841 11679
rect 38945 11645 38979 11679
rect 75101 11645 75135 11679
rect 85681 11645 85715 11679
rect 39129 11577 39163 11611
rect 8401 11509 8435 11543
rect 15025 11509 15059 11543
rect 34897 11509 34931 11543
rect 12173 11305 12207 11339
rect 14197 11305 14231 11339
rect 13369 11237 13403 11271
rect 6469 11169 6503 11203
rect 12357 11169 12391 11203
rect 12633 11169 12667 11203
rect 12909 11169 12943 11203
rect 13037 11169 13071 11203
rect 13185 11169 13219 11203
rect 69029 11305 69063 11339
rect 28365 11237 28399 11271
rect 67189 11237 67223 11271
rect 67925 11237 67959 11271
rect 95985 11305 96019 11339
rect 97549 11305 97583 11339
rect 69397 11237 69431 11271
rect 21465 11169 21499 11203
rect 21741 11169 21775 11203
rect 25421 11169 25455 11203
rect 26617 11169 26651 11203
rect 38209 11169 38243 11203
rect 38393 11169 38427 11203
rect 38577 11169 38611 11203
rect 38945 11169 38979 11203
rect 39129 11169 39163 11203
rect 42625 11169 42659 11203
rect 69029 11169 69063 11203
rect 69121 11169 69155 11203
rect 95985 11169 96019 11203
rect 96353 11169 96387 11203
rect 96721 11169 96755 11203
rect 96997 11169 97031 11203
rect 97089 11169 97123 11203
rect 6745 11101 6779 11135
rect 8125 11101 8159 11135
rect 12817 11101 12851 11135
rect 14197 11101 14231 11135
rect 26709 11101 26743 11135
rect 26985 11101 27019 11135
rect 37749 11101 37783 11135
rect 96169 11101 96203 11135
rect 96537 11101 96571 11135
rect 26617 11033 26651 11067
rect 39405 11033 39439 11067
rect 12541 10965 12575 10999
rect 25237 10965 25271 10999
rect 44833 10761 44867 10795
rect 67281 10693 67315 10727
rect 44557 10625 44591 10659
rect 66361 10625 66395 10659
rect 28365 10557 28399 10591
rect 44189 10557 44223 10591
rect 44337 10557 44371 10591
rect 44465 10557 44499 10591
rect 44741 10557 44775 10591
rect 61853 10557 61887 10591
rect 62129 10557 62163 10591
rect 65349 10557 65383 10591
rect 68753 10557 68787 10591
rect 91017 10557 91051 10591
rect 65257 10489 65291 10523
rect 66361 10489 66395 10523
rect 91293 10489 91327 10523
rect 61669 10421 61703 10455
rect 63233 10421 63267 10455
rect 27261 10217 27295 10251
rect 28089 10217 28123 10251
rect 29929 10217 29963 10251
rect 4905 10149 4939 10183
rect 4353 10081 4387 10115
rect 6653 10081 6687 10115
rect 7297 10081 7331 10115
rect 26137 10081 26171 10115
rect 27997 10081 28031 10115
rect 29929 10081 29963 10115
rect 57437 10217 57471 10251
rect 9413 10013 9447 10047
rect 10885 10013 10919 10047
rect 11161 10013 11195 10047
rect 25881 10013 25915 10047
rect 38117 10013 38151 10047
rect 38393 10013 38427 10047
rect 57529 10217 57563 10251
rect 57529 10081 57563 10115
rect 57713 10081 57747 10115
rect 81173 10081 81207 10115
rect 81725 10081 81759 10115
rect 57989 10013 58023 10047
rect 95893 10013 95927 10047
rect 57437 9945 57471 9979
rect 9781 9877 9815 9911
rect 39681 9877 39715 9911
rect 52469 9877 52503 9911
rect 59553 9877 59587 9911
rect 13001 9605 13035 9639
rect 20361 9605 20395 9639
rect 18889 9537 18923 9571
rect 19349 9537 19383 9571
rect 19441 9537 19475 9571
rect 35541 9537 35575 9571
rect 50905 9537 50939 9571
rect 54309 9537 54343 9571
rect 3249 9469 3283 9503
rect 3433 9469 3467 9503
rect 3617 9469 3651 9503
rect 12449 9469 12483 9503
rect 12725 9469 12759 9503
rect 12817 9469 12851 9503
rect 19165 9469 19199 9503
rect 19533 9469 19567 9503
rect 19717 9469 19751 9503
rect 36001 9469 36035 9503
rect 36277 9469 36311 9503
rect 36369 9469 36403 9503
rect 36645 9469 36679 9503
rect 36829 9469 36863 9503
rect 50629 9469 50663 9503
rect 51089 9469 51123 9503
rect 51365 9469 51399 9503
rect 52285 9469 52319 9503
rect 54033 9469 54067 9503
rect 67373 9469 67407 9503
rect 90741 9469 90775 9503
rect 90833 9469 90867 9503
rect 91017 9469 91051 9503
rect 3709 9401 3743 9435
rect 12633 9401 12667 9435
rect 18981 9333 19015 9367
rect 50629 9333 50663 9367
rect 50813 9333 50847 9367
rect 51273 9333 51307 9367
rect 91201 9333 91235 9367
rect 11437 9129 11471 9163
rect 12265 9129 12299 9163
rect 16681 9129 16715 9163
rect 74457 9129 74491 9163
rect 6009 9061 6043 9095
rect 39773 9061 39807 9095
rect 95525 9061 95559 9095
rect 4721 8993 4755 9027
rect 5089 8993 5123 9027
rect 5457 8993 5491 9027
rect 5641 8993 5675 9027
rect 11621 8993 11655 9027
rect 11804 8993 11838 9027
rect 11989 8993 12023 9027
rect 12173 8993 12207 9027
rect 12449 8993 12483 9027
rect 16497 8993 16531 9027
rect 16773 8993 16807 9027
rect 36921 8993 36955 9027
rect 37104 8993 37138 9027
rect 37473 8993 37507 9027
rect 38393 8993 38427 9027
rect 63049 8993 63083 9027
rect 73813 8993 73847 9027
rect 88809 8993 88843 9027
rect 88993 8993 89027 9027
rect 89361 8993 89395 9027
rect 89453 8993 89487 9027
rect 95157 8993 95191 9027
rect 5181 8925 5215 8959
rect 11897 8925 11931 8959
rect 20821 8925 20855 8959
rect 21097 8925 21131 8959
rect 37197 8925 37231 8959
rect 37289 8925 37323 8959
rect 38117 8925 38151 8959
rect 62773 8925 62807 8959
rect 64153 8925 64187 8959
rect 73960 8925 73994 8959
rect 74181 8925 74215 8959
rect 88441 8925 88475 8959
rect 74089 8857 74123 8891
rect 16313 8789 16347 8823
rect 22201 8789 22235 8823
rect 37565 8789 37599 8823
rect 20453 8585 20487 8619
rect 23673 8585 23707 8619
rect 39497 8585 39531 8619
rect 67281 8585 67315 8619
rect 94145 8585 94179 8619
rect 94605 8585 94639 8619
rect 95157 8585 95191 8619
rect 61117 8517 61151 8551
rect 20085 8449 20119 8483
rect 20177 8449 20211 8483
rect 34345 8449 34379 8483
rect 19809 8381 19843 8415
rect 19992 8381 20026 8415
rect 20361 8381 20395 8415
rect 23029 8381 23063 8415
rect 23122 8381 23156 8415
rect 23305 8381 23339 8415
rect 23535 8381 23569 8415
rect 33701 8381 33735 8415
rect 35449 8381 35483 8415
rect 35725 8381 35759 8415
rect 38853 8381 38887 8415
rect 38946 8381 38980 8415
rect 39221 8381 39255 8415
rect 39359 8381 39393 8415
rect 49249 8381 49283 8415
rect 50709 8381 50743 8415
rect 50997 8381 51031 8415
rect 54309 8381 54343 8415
rect 56609 8381 56643 8415
rect 61117 8381 61151 8415
rect 61301 8381 61335 8415
rect 65993 8381 66027 8415
rect 94467 8517 94501 8551
rect 94697 8449 94731 8483
rect 94789 8449 94823 8483
rect 67465 8381 67499 8415
rect 23397 8313 23431 8347
rect 35265 8313 35299 8347
rect 35633 8313 35667 8347
rect 39129 8313 39163 8347
rect 50537 8313 50571 8347
rect 50905 8313 50939 8347
rect 61853 8313 61887 8347
rect 66361 8313 66395 8347
rect 67281 8313 67315 8347
rect 67833 8313 67867 8347
rect 94329 8313 94363 8347
rect 33333 8041 33367 8075
rect 1409 7905 1443 7939
rect 1777 7905 1811 7939
rect 2053 7905 2087 7939
rect 2145 7905 2179 7939
rect 10425 7905 10459 7939
rect 10793 7905 10827 7939
rect 10977 7905 11011 7939
rect 31953 7905 31987 7939
rect 32229 7905 32263 7939
rect 37289 7905 37323 7939
rect 37657 7905 37691 7939
rect 38025 7905 38059 7939
rect 39129 7905 39163 7939
rect 39313 7905 39347 7939
rect 39405 7905 39439 7939
rect 39549 7905 39583 7939
rect 94513 7905 94547 7939
rect 1869 7837 1903 7871
rect 2697 7837 2731 7871
rect 10057 7837 10091 7871
rect 10517 7837 10551 7871
rect 37565 7837 37599 7871
rect 38117 7837 38151 7871
rect 39698 7837 39732 7871
rect 94789 7837 94823 7871
rect 9689 7769 9723 7803
rect 38485 7769 38519 7803
rect 25053 7497 25087 7531
rect 69581 7497 69615 7531
rect 69949 7497 69983 7531
rect 11897 7429 11931 7463
rect 12265 7429 12299 7463
rect 24961 7429 24995 7463
rect 27169 7429 27203 7463
rect 9597 7361 9631 7395
rect 25421 7361 25455 7395
rect 25513 7361 25547 7395
rect 9137 7293 9171 7327
rect 9505 7293 9539 7327
rect 9873 7293 9907 7327
rect 10057 7293 10091 7327
rect 25237 7293 25271 7327
rect 25605 7293 25639 7327
rect 25789 7293 25823 7327
rect 25973 7293 26007 7327
rect 87061 7361 87095 7395
rect 38577 7293 38611 7327
rect 49238 7293 49272 7327
rect 49433 7293 49467 7327
rect 49617 7293 49651 7327
rect 49893 7293 49927 7327
rect 50031 7293 50065 7327
rect 50537 7293 50571 7327
rect 86877 7293 86911 7327
rect 97917 7293 97951 7327
rect 10425 7225 10459 7259
rect 27169 7225 27203 7259
rect 4905 6817 4939 6851
rect 5273 6817 5307 6851
rect 5641 6817 5675 6851
rect 43361 6817 43395 6851
rect 62221 6817 62255 6851
rect 63601 6817 63635 6851
rect 72433 6817 72467 6851
rect 72617 6817 72651 6851
rect 72801 6817 72835 6851
rect 72893 6817 72927 6851
rect 97549 6817 97583 6851
rect 4997 6749 5031 6783
rect 5457 6749 5491 6783
rect 61945 6749 61979 6783
rect 3525 6613 3559 6647
rect 3709 6613 3743 6647
rect 3985 6613 4019 6647
rect 4169 6613 4203 6647
rect 4445 6613 4479 6647
rect 5825 6613 5859 6647
rect 6009 6613 6043 6647
rect 6193 6613 6227 6647
rect 6377 6613 6411 6647
rect 6561 6613 6595 6647
rect 82093 6409 82127 6443
rect 96077 6409 96111 6443
rect 96261 6409 96295 6443
rect 15853 6341 15887 6375
rect 21097 6341 21131 6375
rect 21235 6341 21269 6375
rect 51457 6341 51491 6375
rect 15485 6273 15519 6307
rect 86601 6273 86635 6307
rect 3341 6205 3375 6239
rect 4353 6205 4387 6239
rect 15117 6205 15151 6239
rect 15301 6205 15335 6239
rect 15393 6205 15427 6239
rect 15669 6205 15703 6239
rect 21034 6205 21068 6239
rect 33149 6205 33183 6239
rect 34437 6205 34471 6239
rect 51273 6205 51307 6239
rect 52745 6205 52779 6239
rect 53014 6205 53048 6239
rect 81541 6205 81575 6239
rect 81909 6205 81943 6239
rect 85957 6205 85991 6239
rect 96997 6205 97031 6239
rect 97641 6205 97675 6239
rect 15025 6137 15059 6171
rect 21373 6137 21407 6171
rect 33701 6137 33735 6171
rect 81725 6137 81759 6171
rect 81817 6137 81851 6171
rect 20545 6069 20579 6103
rect 20729 6069 20763 6103
rect 8309 5865 8343 5899
rect 73905 5865 73939 5899
rect 95893 5865 95927 5899
rect 7389 5797 7423 5831
rect 2421 5729 2455 5763
rect 3065 5729 3099 5763
rect 4445 5729 4479 5763
rect 7021 5729 7055 5763
rect 7665 5729 7699 5763
rect 7848 5729 7882 5763
rect 8217 5729 8251 5763
rect 8585 5729 8619 5763
rect 26525 5729 26559 5763
rect 74089 5729 74123 5763
rect 95249 5729 95283 5763
rect 95432 5729 95466 5763
rect 95525 5729 95559 5763
rect 95801 5729 95835 5763
rect 96445 5729 96479 5763
rect 97549 5729 97583 5763
rect 7941 5661 7975 5695
rect 8033 5661 8067 5695
rect 26249 5661 26283 5695
rect 95617 5661 95651 5695
rect 5089 5525 5123 5559
rect 7389 5525 7423 5559
rect 7573 5525 7607 5559
rect 27629 5525 27663 5559
rect 95065 5525 95099 5559
rect 6469 5321 6503 5355
rect 24317 5321 24351 5355
rect 65257 5321 65291 5355
rect 79701 5321 79735 5355
rect 6285 5253 6319 5287
rect 2421 5185 2455 5219
rect 2697 5185 2731 5219
rect 2881 5185 2915 5219
rect 3341 5117 3375 5151
rect 5641 5117 5675 5151
rect 34345 5253 34379 5287
rect 38485 5253 38519 5287
rect 8585 5185 8619 5219
rect 12541 5185 12575 5219
rect 23213 5185 23247 5219
rect 6469 5117 6503 5151
rect 6837 5117 6871 5151
rect 8033 5117 8067 5151
rect 9137 5117 9171 5151
rect 22937 5117 22971 5151
rect 25053 5117 25087 5151
rect 25697 5117 25731 5151
rect 26341 5117 26375 5151
rect 27813 5117 27847 5151
rect 33793 5117 33827 5151
rect 34161 5117 34195 5151
rect 36369 5117 36403 5151
rect 36645 5117 36679 5151
rect 36829 5117 36863 5151
rect 36921 5117 36955 5151
rect 1869 5049 1903 5083
rect 4353 5049 4387 5083
rect 6285 5049 6319 5083
rect 7021 5049 7055 5083
rect 33977 5049 34011 5083
rect 34069 5049 34103 5083
rect 45293 5185 45327 5219
rect 82737 5185 82771 5219
rect 91385 5185 91419 5219
rect 38761 5117 38795 5151
rect 39221 5117 39255 5151
rect 44925 5117 44959 5151
rect 64705 5117 64739 5151
rect 64889 5117 64923 5151
rect 65073 5117 65107 5151
rect 76941 5117 76975 5151
rect 77585 5117 77619 5151
rect 79701 5117 79735 5151
rect 82093 5117 82127 5151
rect 82461 5117 82495 5151
rect 85865 5117 85899 5151
rect 87337 5117 87371 5151
rect 87613 5117 87647 5151
rect 88073 5117 88107 5151
rect 88717 5117 88751 5151
rect 90741 5117 90775 5151
rect 90925 5117 90959 5151
rect 91109 5117 91143 5151
rect 91477 5117 91511 5151
rect 92949 5117 92983 5151
rect 94237 5117 94271 5151
rect 94881 5117 94915 5151
rect 95985 5117 96019 5151
rect 97181 5117 97215 5151
rect 97825 5117 97859 5151
rect 64981 5049 65015 5083
rect 82277 5049 82311 5083
rect 85957 5049 85991 5083
rect 1961 4981 1995 5015
rect 3433 4981 3467 5015
rect 4445 4981 4479 5015
rect 5733 4981 5767 5015
rect 6745 4981 6779 5015
rect 36461 4981 36495 5015
rect 38485 4981 38519 5015
rect 90097 4981 90131 5015
rect 90373 4981 90407 5015
rect 90557 4981 90591 5015
rect 91937 4981 91971 5015
rect 92213 4981 92247 5015
rect 92397 4981 92431 5015
rect 92581 4981 92615 5015
rect 92765 4981 92799 5015
rect 1961 4777 1995 4811
rect 2513 4777 2547 4811
rect 6837 4777 6871 4811
rect 7021 4777 7055 4811
rect 7573 4777 7607 4811
rect 32873 4777 32907 4811
rect 53297 4777 53331 4811
rect 53941 4777 53975 4811
rect 54125 4777 54159 4811
rect 2881 4709 2915 4743
rect 6653 4709 6687 4743
rect 7297 4709 7331 4743
rect 7665 4709 7699 4743
rect 7941 4709 7975 4743
rect 26985 4709 27019 4743
rect 39037 4709 39071 4743
rect 1869 4641 1903 4675
rect 3985 4641 4019 4675
rect 4169 4641 4203 4675
rect 4353 4641 4387 4675
rect 4537 4641 4571 4675
rect 4721 4641 4755 4675
rect 4905 4641 4939 4675
rect 5273 4641 5307 4675
rect 9505 4641 9539 4675
rect 10609 4641 10643 4675
rect 11253 4641 11287 4675
rect 11897 4641 11931 4675
rect 12541 4641 12575 4675
rect 14749 4641 14783 4675
rect 15393 4641 15427 4675
rect 16129 4641 16163 4675
rect 17325 4641 17359 4675
rect 17969 4641 18003 4675
rect 18613 4641 18647 4675
rect 19993 4641 20027 4675
rect 21005 4641 21039 4675
rect 22017 4641 22051 4675
rect 22661 4641 22695 4675
rect 23305 4641 23339 4675
rect 25697 4641 25731 4675
rect 26065 4641 26099 4675
rect 26341 4641 26375 4675
rect 26433 4641 26467 4675
rect 27537 4641 27571 4675
rect 29101 4641 29135 4675
rect 33149 4641 33183 4675
rect 34253 4641 34287 4675
rect 36093 4641 36127 4675
rect 36737 4641 36771 4675
rect 37289 4641 37323 4675
rect 37657 4641 37691 4675
rect 39497 4641 39531 4675
rect 40969 4641 41003 4675
rect 41613 4641 41647 4675
rect 44005 4641 44039 4675
rect 44649 4641 44683 4675
rect 46213 4641 46247 4675
rect 47041 4641 47075 4675
rect 47685 4641 47719 4675
rect 52561 4641 52595 4675
rect 53481 4641 53515 4675
rect 53665 4641 53699 4675
rect 53849 4641 53883 4675
rect 54125 4641 54159 4675
rect 54217 4777 54251 4811
rect 4997 4573 5031 4607
rect 26157 4573 26191 4607
rect 37381 4573 37415 4607
rect 65625 4709 65659 4743
rect 78229 4709 78263 4743
rect 54309 4641 54343 4675
rect 61945 4641 61979 4675
rect 62128 4641 62162 4675
rect 62313 4641 62347 4675
rect 62497 4641 62531 4675
rect 64245 4641 64279 4675
rect 66085 4641 66119 4675
rect 68385 4641 68419 4675
rect 70777 4641 70811 4675
rect 73813 4641 73847 4675
rect 76297 4641 76331 4675
rect 77953 4641 77987 4675
rect 78137 4641 78171 4675
rect 78689 4641 78723 4675
rect 79333 4641 79367 4675
rect 79977 4641 80011 4675
rect 80621 4641 80655 4675
rect 81265 4641 81299 4675
rect 82921 4641 82955 4675
rect 83565 4641 83599 4675
rect 85405 4641 85439 4675
rect 86049 4641 86083 4675
rect 88165 4641 88199 4675
rect 88809 4641 88843 4675
rect 89453 4641 89487 4675
rect 90097 4641 90131 4675
rect 90741 4641 90775 4675
rect 91385 4641 91419 4675
rect 92029 4641 92063 4675
rect 93409 4641 93443 4675
rect 94053 4641 94087 4675
rect 94697 4641 94731 4675
rect 95341 4641 95375 4675
rect 95985 4641 96019 4675
rect 96629 4641 96663 4675
rect 97273 4641 97307 4675
rect 62221 4573 62255 4607
rect 63509 4573 63543 4607
rect 63969 4573 64003 4607
rect 2697 4505 2731 4539
rect 7113 4505 7147 4539
rect 8125 4505 8159 4539
rect 54217 4505 54251 4539
rect 77769 4505 77803 4539
rect 28641 4437 28675 4471
rect 42809 4437 42843 4471
rect 62589 4437 62623 4471
rect 87061 4437 87095 4471
rect 3801 4165 3835 4199
rect 19993 4165 20027 4199
rect 86877 4165 86911 4199
rect 2973 4097 3007 4131
rect 34989 4097 35023 4131
rect 88165 4097 88199 4131
rect 91845 4097 91879 4131
rect 92305 4097 92339 4131
rect 96997 4097 97031 4131
rect 2697 4029 2731 4063
rect 3617 4029 3651 4063
rect 4721 4029 4755 4063
rect 6837 4029 6871 4063
rect 7757 4029 7791 4063
rect 9413 4029 9447 4063
rect 10057 4029 10091 4063
rect 10701 4029 10735 4063
rect 12357 4029 12391 4063
rect 12909 4029 12943 4063
rect 13185 4029 13219 4063
rect 13645 4029 13679 4063
rect 14289 4029 14323 4063
rect 16037 4029 16071 4063
rect 17325 4029 17359 4063
rect 18429 4029 18463 4063
rect 20453 4029 20487 4063
rect 21097 4029 21131 4063
rect 23029 4029 23063 4063
rect 23489 4029 23523 4063
rect 24409 4029 24443 4063
rect 25053 4029 25087 4063
rect 25605 4029 25639 4063
rect 25881 4029 25915 4063
rect 26341 4029 26375 4063
rect 27813 4029 27847 4063
rect 28457 4029 28491 4063
rect 29101 4029 29135 4063
rect 29745 4029 29779 4063
rect 31217 4029 31251 4063
rect 33057 4029 33091 4063
rect 33701 4029 33735 4063
rect 34437 4029 34471 4063
rect 35541 4029 35575 4063
rect 36185 4029 36219 4063
rect 36829 4029 36863 4063
rect 38669 4029 38703 4063
rect 39313 4029 39347 4063
rect 39957 4029 39991 4063
rect 40601 4029 40635 4063
rect 41245 4029 41279 4063
rect 41889 4029 41923 4063
rect 43545 4029 43579 4063
rect 44189 4029 44223 4063
rect 45385 4029 45419 4063
rect 46029 4029 46063 4063
rect 46673 4029 46707 4063
rect 47317 4029 47351 4063
rect 48789 4029 48823 4063
rect 49433 4029 49467 4063
rect 50077 4029 50111 4063
rect 50721 4029 50755 4063
rect 51365 4029 51399 4063
rect 52009 4029 52043 4063
rect 52653 4029 52687 4063
rect 54033 4029 54067 4063
rect 54677 4029 54711 4063
rect 55321 4029 55355 4063
rect 55965 4029 55999 4063
rect 56609 4029 56643 4063
rect 57253 4029 57287 4063
rect 57897 4029 57931 4063
rect 59277 4029 59311 4063
rect 59921 4029 59955 4063
rect 60565 4029 60599 4063
rect 61209 4029 61243 4063
rect 61845 4029 61879 4063
rect 62497 4029 62531 4063
rect 63133 4029 63167 4063
rect 64521 4029 64555 4063
rect 65165 4029 65199 4063
rect 65809 4029 65843 4063
rect 66453 4029 66487 4063
rect 67097 4029 67131 4063
rect 67741 4029 67775 4063
rect 68385 4029 68419 4063
rect 69765 4029 69799 4063
rect 70409 4029 70443 4063
rect 71053 4029 71087 4063
rect 71697 4029 71731 4063
rect 72341 4029 72375 4063
rect 72985 4029 73019 4063
rect 73629 4029 73663 4063
rect 75009 4029 75043 4063
rect 75653 4029 75687 4063
rect 76297 4029 76331 4063
rect 77125 4029 77159 4063
rect 78321 4029 78355 4063
rect 78965 4029 78999 4063
rect 80805 4029 80839 4063
rect 81449 4029 81483 4063
rect 82093 4029 82127 4063
rect 82737 4029 82771 4063
rect 83657 4029 83691 4063
rect 84301 4029 84335 4063
rect 85497 4029 85531 4063
rect 87889 4029 87923 4063
rect 91201 4029 91235 4063
rect 91385 4029 91419 4063
rect 91569 4029 91603 4063
rect 91937 4029 91971 4063
rect 93041 4029 93075 4063
rect 93685 4029 93719 4063
rect 94329 4029 94363 4063
rect 95985 4029 96019 4063
rect 97181 4029 97215 4063
rect 97733 4029 97767 4063
rect 97917 4029 97951 4063
rect 1869 3961 1903 3995
rect 2237 3961 2271 3995
rect 4353 3961 4387 3995
rect 4997 3961 5031 3995
rect 5733 3961 5767 3995
rect 8677 3961 8711 3995
rect 15393 3961 15427 3995
rect 19165 3961 19199 3995
rect 91109 3961 91143 3995
rect 97365 3961 97399 3995
rect 4445 3893 4479 3927
rect 5825 3893 5859 3927
rect 7021 3893 7055 3927
rect 7941 3893 7975 3927
rect 8769 3893 8803 3927
rect 9505 3893 9539 3927
rect 12449 3893 12483 3927
rect 15485 3893 15519 3927
rect 18521 3893 18555 3927
rect 19257 3893 19291 3927
rect 23489 3893 23523 3927
rect 89269 3893 89303 3927
rect 98009 3893 98043 3927
rect 11897 3689 11931 3723
rect 40417 3689 40451 3723
rect 81449 3689 81483 3723
rect 3065 3621 3099 3655
rect 4721 3621 4755 3655
rect 5549 3621 5583 3655
rect 6285 3621 6319 3655
rect 8125 3621 8159 3655
rect 11069 3621 11103 3655
rect 13277 3621 13311 3655
rect 14841 3621 14875 3655
rect 15577 3621 15611 3655
rect 17894 3621 17928 3655
rect 20821 3621 20855 3655
rect 21557 3621 21591 3655
rect 37381 3621 37415 3655
rect 1869 3553 1903 3587
rect 2789 3553 2823 3587
rect 4353 3553 4387 3587
rect 6929 3553 6963 3587
rect 7849 3553 7883 3587
rect 9597 3553 9631 3587
rect 10333 3553 10367 3587
rect 11805 3553 11839 3587
rect 12541 3553 12575 3587
rect 16313 3553 16347 3587
rect 17141 3553 17175 3587
rect 18521 3553 18555 3587
rect 20085 3553 20119 3587
rect 21005 3553 21039 3587
rect 22201 3553 22235 3587
rect 22845 3553 22879 3587
rect 24041 3553 24075 3587
rect 25237 3553 25271 3587
rect 25881 3553 25915 3587
rect 26801 3553 26835 3587
rect 27721 3553 27755 3587
rect 28917 3553 28951 3587
rect 30481 3553 30515 3587
rect 31125 3553 31159 3587
rect 31953 3553 31987 3587
rect 32597 3553 32631 3587
rect 33241 3553 33275 3587
rect 34437 3553 34471 3587
rect 35725 3553 35759 3587
rect 36369 3553 36403 3587
rect 37749 3553 37783 3587
rect 38945 3553 38979 3587
rect 39589 3553 39623 3587
rect 2145 3485 2179 3519
rect 7113 3485 7147 3519
rect 16865 3485 16899 3519
rect 81725 3621 81759 3655
rect 96629 3621 96663 3655
rect 96813 3621 96847 3655
rect 40969 3553 41003 3587
rect 41705 3553 41739 3587
rect 42349 3553 42383 3587
rect 42993 3553 43027 3587
rect 43637 3553 43671 3587
rect 44833 3553 44867 3587
rect 47225 3553 47259 3587
rect 47869 3553 47903 3587
rect 48513 3553 48547 3587
rect 49157 3553 49191 3587
rect 49793 3553 49827 3587
rect 51457 3553 51491 3587
rect 52101 3553 52135 3587
rect 52745 3553 52779 3587
rect 53389 3553 53423 3587
rect 54033 3553 54067 3587
rect 54677 3553 54711 3587
rect 55321 3553 55355 3587
rect 56701 3553 56735 3587
rect 57345 3553 57379 3587
rect 58173 3553 58207 3587
rect 58817 3553 58851 3587
rect 59461 3553 59495 3587
rect 60657 3553 60691 3587
rect 61945 3553 61979 3587
rect 62589 3553 62623 3587
rect 63233 3553 63267 3587
rect 63877 3553 63911 3587
rect 64521 3553 64555 3587
rect 65165 3553 65199 3587
rect 65809 3553 65843 3587
rect 67189 3553 67223 3587
rect 67925 3553 67959 3587
rect 68569 3553 68603 3587
rect 69213 3553 69247 3587
rect 69857 3553 69891 3587
rect 70501 3553 70535 3587
rect 71145 3553 71179 3587
rect 72433 3553 72467 3587
rect 73077 3553 73111 3587
rect 74089 3553 74123 3587
rect 74733 3553 74767 3587
rect 75929 3553 75963 3587
rect 76573 3553 76607 3587
rect 78321 3553 78355 3587
rect 79333 3553 79367 3587
rect 79885 3553 79919 3587
rect 80529 3553 80563 3587
rect 83013 3553 83047 3587
rect 84301 3553 84335 3587
rect 84945 3553 84979 3587
rect 85589 3553 85623 3587
rect 86233 3553 86267 3587
rect 86877 3553 86911 3587
rect 88165 3553 88199 3587
rect 88809 3553 88843 3587
rect 89453 3553 89487 3587
rect 90097 3553 90131 3587
rect 90741 3553 90775 3587
rect 91385 3553 91419 3587
rect 92029 3553 92063 3587
rect 93409 3553 93443 3587
rect 94053 3553 94087 3587
rect 94881 3553 94915 3587
rect 95157 3553 95191 3587
rect 95709 3553 95743 3587
rect 97549 3553 97583 3587
rect 15761 3417 15795 3451
rect 16957 3417 16991 3451
rect 17693 3417 17727 3451
rect 21741 3417 21775 3451
rect 40417 3417 40451 3451
rect 78965 3417 78999 3451
rect 79149 3417 79183 3451
rect 81541 3417 81575 3451
rect 83841 3417 83875 3451
rect 94973 3417 95007 3451
rect 96997 3417 97031 3451
rect 9689 3349 9723 3383
rect 10425 3349 10459 3383
rect 11161 3349 11195 3383
rect 12633 3349 12667 3383
rect 13369 3349 13403 3383
rect 14933 3349 14967 3383
rect 16405 3349 16439 3383
rect 17601 3349 17635 3383
rect 18613 3349 18647 3383
rect 20177 3349 20211 3383
rect 26893 3349 26927 3383
rect 46765 3349 46799 3383
rect 77861 3349 77895 3383
rect 97641 3349 97675 3383
rect 4261 3145 4295 3179
rect 14381 3145 14415 3179
rect 15945 3145 15979 3179
rect 20269 3145 20303 3179
rect 21005 3145 21039 3179
rect 38117 3145 38151 3179
rect 74825 3145 74859 3179
rect 76389 3145 76423 3179
rect 76481 3145 76515 3179
rect 78505 3145 78539 3179
rect 80713 3145 80747 3179
rect 80805 3145 80839 3179
rect 81541 3145 81575 3179
rect 85681 3145 85715 3179
rect 89085 3145 89119 3179
rect 90465 3145 90499 3179
rect 90557 3145 90591 3179
rect 94421 3145 94455 3179
rect 95801 3145 95835 3179
rect 97273 3145 97307 3179
rect 5089 3077 5123 3111
rect 22017 3077 22051 3111
rect 66821 3077 66855 3111
rect 69489 3077 69523 3111
rect 69581 3077 69615 3111
rect 2145 3009 2179 3043
rect 3341 3009 3375 3043
rect 7205 3009 7239 3043
rect 10885 3009 10919 3043
rect 13553 3009 13587 3043
rect 17509 3009 17543 3043
rect 1593 2941 1627 2975
rect 2789 2941 2823 2975
rect 3985 2941 4019 2975
rect 5733 2941 5767 2975
rect 7757 2941 7791 2975
rect 8033 2941 8067 2975
rect 10333 2941 10367 2975
rect 12081 2941 12115 2975
rect 13277 2941 13311 2975
rect 14197 2941 14231 2975
rect 15025 2941 15059 2975
rect 15761 2941 15795 2975
rect 17325 2941 17359 2975
rect 18245 2941 18279 2975
rect 19165 2941 19199 2975
rect 20085 2941 20119 2975
rect 35541 3009 35575 3043
rect 46949 3009 46983 3043
rect 55229 3009 55263 3043
rect 71605 3009 71639 3043
rect 23305 2941 23339 2975
rect 23949 2941 23983 2975
rect 25053 2941 25087 2975
rect 25605 2941 25639 2975
rect 27629 2941 27663 2975
rect 27997 2941 28031 2975
rect 28365 2941 28399 2975
rect 28733 2941 28767 2975
rect 29193 2941 29227 2975
rect 29837 2941 29871 2975
rect 30481 2941 30515 2975
rect 31125 2941 31159 2975
rect 31769 2941 31803 2975
rect 33057 2941 33091 2975
rect 33701 2941 33735 2975
rect 34345 2941 34379 2975
rect 35357 2941 35391 2975
rect 36369 2941 36403 2975
rect 37013 2941 37047 2975
rect 39037 2941 39071 2975
rect 40233 2941 40267 2975
rect 42073 2941 42107 2975
rect 44281 2941 44315 2975
rect 44925 2941 44959 2975
rect 45477 2941 45511 2975
rect 45753 2941 45787 2975
rect 46397 2941 46431 2975
rect 47041 2941 47075 2975
rect 47225 2941 47259 2975
rect 48881 2941 48915 2975
rect 49433 2941 49467 2975
rect 49709 2941 49743 2975
rect 50261 2941 50295 2975
rect 51825 2941 51859 2975
rect 52469 2941 52503 2975
rect 54125 2941 54159 2975
rect 55505 2941 55539 2975
rect 56701 2941 56735 2975
rect 57345 2941 57379 2975
rect 57989 2941 58023 2975
rect 59369 2941 59403 2975
rect 60013 2941 60047 2975
rect 60657 2941 60691 2975
rect 62773 2941 62807 2975
rect 63601 2941 63635 2975
rect 65257 2941 65291 2975
rect 65901 2941 65935 2975
rect 67097 2941 67131 2975
rect 67649 2941 67683 2975
rect 68293 2941 68327 2975
rect 69489 2941 69523 2975
rect 69949 2941 69983 2975
rect 70501 2941 70535 2975
rect 70777 2941 70811 2975
rect 71329 2941 71363 2975
rect 71512 2941 71546 2975
rect 71697 2941 71731 2975
rect 71881 2941 71915 2975
rect 73261 2941 73295 2975
rect 73905 2941 73939 2975
rect 75193 2941 75227 2975
rect 75745 2941 75779 2975
rect 76389 2941 76423 2975
rect 76849 2941 76883 2975
rect 78045 2941 78079 2975
rect 78689 2941 78723 2975
rect 78873 2941 78907 2975
rect 80161 2941 80195 2975
rect 80437 2941 80471 2975
rect 4905 2873 4939 2907
rect 6929 2873 6963 2907
rect 9137 2873 9171 2907
rect 12357 2873 12391 2907
rect 18521 2873 18555 2907
rect 19441 2873 19475 2907
rect 20913 2873 20947 2907
rect 22017 2873 22051 2907
rect 22661 2873 22695 2907
rect 26341 2873 26375 2907
rect 27813 2873 27847 2907
rect 38301 2873 38335 2907
rect 38485 2873 38519 2907
rect 41429 2873 41463 2907
rect 43637 2873 43671 2907
rect 45569 2873 45603 2907
rect 49525 2873 49559 2907
rect 51181 2873 51215 2907
rect 55321 2873 55355 2907
rect 61577 2873 61611 2907
rect 64521 2873 64555 2907
rect 64705 2873 64739 2907
rect 66913 2873 66947 2907
rect 69765 2873 69799 2907
rect 70593 2873 70627 2907
rect 72617 2873 72651 2907
rect 75009 2873 75043 2907
rect 76665 2873 76699 2907
rect 80253 2873 80287 2907
rect 96721 3009 96755 3043
rect 81725 2941 81759 2975
rect 81909 2941 81943 2975
rect 82553 2941 82587 2975
rect 83197 2941 83231 2975
rect 83841 2941 83875 2975
rect 86601 2941 86635 2975
rect 87705 2941 87739 2975
rect 87981 2941 88015 2975
rect 90465 2941 90499 2975
rect 90925 2941 90959 2975
rect 91569 2941 91603 2975
rect 92305 2941 92339 2975
rect 93961 2941 93995 2975
rect 94605 2941 94639 2975
rect 94789 2941 94823 2975
rect 97457 2941 97491 2975
rect 97641 2941 97675 2975
rect 80989 2873 81023 2907
rect 81173 2873 81207 2907
rect 85865 2873 85899 2907
rect 86049 2873 86083 2907
rect 90741 2873 90775 2907
rect 93133 2873 93167 2907
rect 93317 2873 93351 2907
rect 95985 2873 96019 2907
rect 96169 2873 96203 2907
rect 96629 2873 96663 2907
rect 96905 2873 96939 2907
rect 9229 2805 9263 2839
rect 15117 2805 15151 2839
rect 22753 2805 22787 2839
rect 25697 2805 25731 2839
rect 26433 2805 26467 2839
rect 36461 2805 36495 2839
rect 40325 2805 40359 2839
rect 41521 2805 41555 2839
rect 43729 2805 43763 2839
rect 46489 2805 46523 2839
rect 48973 2805 49007 2839
rect 51273 2805 51307 2839
rect 54217 2805 54251 2839
rect 56793 2805 56827 2839
rect 59461 2805 59495 2839
rect 61669 2805 61703 2839
rect 62865 2805 62899 2839
rect 64429 2805 64463 2839
rect 71973 2805 72007 2839
rect 72709 2805 72743 2839
rect 78137 2805 78171 2839
rect 80713 2805 80747 2839
rect 82645 2805 82679 2839
rect 91661 2805 91695 2839
rect 92397 2805 92431 2839
rect 92949 2805 92983 2839
rect 94053 2805 94087 2839
rect 8401 2601 8435 2635
rect 11069 2601 11103 2635
rect 15301 2601 15335 2635
rect 36369 2601 36403 2635
rect 37933 2601 37967 2635
rect 41797 2601 41831 2635
rect 43269 2601 43303 2635
rect 44833 2601 44867 2635
rect 47869 2601 47903 2635
rect 48329 2601 48363 2635
rect 49893 2601 49927 2635
rect 53205 2601 53239 2635
rect 56609 2601 56643 2635
rect 57437 2601 57471 2635
rect 61117 2601 61151 2635
rect 61577 2601 61611 2635
rect 64613 2601 64647 2635
rect 66729 2601 66763 2635
rect 67005 2601 67039 2635
rect 68109 2601 68143 2635
rect 68845 2601 68879 2635
rect 74181 2601 74215 2635
rect 77953 2601 77987 2635
rect 79517 2601 79551 2635
rect 80253 2601 80287 2635
rect 85773 2601 85807 2635
rect 89453 2601 89487 2635
rect 90189 2601 90223 2635
rect 90925 2601 90959 2635
rect 92121 2601 92155 2635
rect 94789 2601 94823 2635
rect 7389 2533 7423 2567
rect 10149 2533 10183 2567
rect 13461 2533 13495 2567
rect 17877 2533 17911 2567
rect 18797 2533 18831 2567
rect 20545 2533 20579 2567
rect 21649 2533 21683 2567
rect 22845 2533 22879 2567
rect 23121 2533 23155 2567
rect 23765 2533 23799 2567
rect 25421 2533 25455 2567
rect 25789 2533 25823 2567
rect 27077 2533 27111 2567
rect 28181 2533 28215 2567
rect 28457 2533 28491 2567
rect 31033 2533 31067 2567
rect 32505 2533 32539 2567
rect 33701 2533 33735 2567
rect 34437 2533 34471 2567
rect 35173 2533 35207 2567
rect 36093 2533 36127 2567
rect 37841 2533 37875 2567
rect 38853 2533 38887 2567
rect 39129 2533 39163 2567
rect 39589 2533 39623 2567
rect 39865 2533 39899 2567
rect 40325 2533 40359 2567
rect 40601 2533 40635 2567
rect 40785 2533 40819 2567
rect 42441 2533 42475 2567
rect 43177 2533 43211 2567
rect 44189 2533 44223 2567
rect 44465 2533 44499 2567
rect 45201 2533 45235 2567
rect 45845 2533 45879 2567
rect 47777 2533 47811 2567
rect 48605 2533 48639 2567
rect 48789 2533 48823 2567
rect 52377 2533 52411 2567
rect 53113 2533 53147 2567
rect 53849 2533 53883 2567
rect 55045 2533 55079 2567
rect 55781 2533 55815 2567
rect 55965 2533 55999 2567
rect 56517 2533 56551 2567
rect 57805 2533 57839 2567
rect 58357 2533 58391 2567
rect 59185 2533 59219 2567
rect 60197 2533 60231 2567
rect 60473 2533 60507 2567
rect 62865 2533 62899 2567
rect 63141 2533 63175 2567
rect 63785 2533 63819 2567
rect 65717 2533 65751 2567
rect 66269 2533 66303 2567
rect 66545 2533 66579 2567
rect 67281 2533 67315 2567
rect 67465 2533 67499 2567
rect 68477 2533 68511 2567
rect 69213 2533 69247 2567
rect 69857 2533 69891 2567
rect 71053 2533 71087 2567
rect 71973 2533 72007 2567
rect 73721 2533 73755 2567
rect 74549 2533 74583 2567
rect 75009 2533 75043 2567
rect 75285 2533 75319 2567
rect 77861 2533 77895 2567
rect 79885 2533 79919 2567
rect 80621 2533 80655 2567
rect 82001 2533 82035 2567
rect 82185 2533 82219 2567
rect 82737 2533 82771 2567
rect 83013 2533 83047 2567
rect 87061 2533 87095 2567
rect 87797 2533 87831 2567
rect 89637 2533 89671 2567
rect 89821 2533 89855 2567
rect 90557 2533 90591 2567
rect 91293 2533 91327 2567
rect 92489 2533 92523 2567
rect 93852 2533 93886 2567
rect 95157 2533 95191 2567
rect 96721 2533 96755 2567
rect 1777 2465 1811 2499
rect 4353 2465 4387 2499
rect 5549 2465 5583 2499
rect 7021 2465 7055 2499
rect 8309 2465 8343 2499
rect 9689 2465 9723 2499
rect 10885 2465 10919 2499
rect 12357 2465 12391 2499
rect 13185 2465 13219 2499
rect 15025 2465 15059 2499
rect 15853 2465 15887 2499
rect 17601 2465 17635 2499
rect 18521 2465 18555 2499
rect 20269 2465 20303 2499
rect 21281 2465 21315 2499
rect 24501 2465 24535 2499
rect 26249 2465 26283 2499
rect 26525 2465 26559 2499
rect 26893 2465 26927 2499
rect 27261 2465 27295 2499
rect 29101 2465 29135 2499
rect 29837 2465 29871 2499
rect 31769 2465 31803 2499
rect 36461 2465 36495 2499
rect 36921 2465 36955 2499
rect 37197 2465 37231 2499
rect 41705 2465 41739 2499
rect 46029 2465 46063 2499
rect 47041 2465 47075 2499
rect 50077 2465 50111 2499
rect 50261 2465 50295 2499
rect 50353 2465 50387 2499
rect 50905 2465 50939 2499
rect 58541 2465 58575 2499
rect 60933 2465 60967 2499
rect 61209 2465 61243 2499
rect 61945 2465 61979 2499
rect 62957 2465 62991 2499
rect 64521 2465 64555 2499
rect 67097 2465 67131 2499
rect 71789 2465 71823 2499
rect 72617 2465 72651 2499
rect 75101 2465 75135 2499
rect 76389 2465 76423 2499
rect 77125 2465 77159 2499
rect 78689 2465 78723 2499
rect 79149 2465 79183 2499
rect 80437 2465 80471 2499
rect 84393 2465 84427 2499
rect 84669 2465 84703 2499
rect 88441 2465 88475 2499
rect 88625 2465 88659 2499
rect 90373 2465 90407 2499
rect 92305 2465 92339 2499
rect 93133 2465 93167 2499
rect 94973 2465 95007 2499
rect 95801 2465 95835 2499
rect 96537 2465 96571 2499
rect 97917 2465 97951 2499
rect 2605 2397 2639 2431
rect 4905 2397 4939 2431
rect 16129 2397 16163 2431
rect 25605 2397 25639 2431
rect 32689 2397 32723 2431
rect 39681 2397 39715 2431
rect 44281 2397 44315 2431
rect 48421 2397 48455 2431
rect 52561 2397 52595 2431
rect 59369 2397 59403 2431
rect 73905 2397 73939 2431
rect 77309 2397 77343 2431
rect 22937 2329 22971 2363
rect 24685 2329 24719 2363
rect 26341 2329 26375 2363
rect 28273 2329 28307 2363
rect 30021 2329 30055 2363
rect 31953 2329 31987 2363
rect 34621 2329 34655 2363
rect 37013 2329 37047 2363
rect 38945 2329 38979 2363
rect 42625 2329 42659 2363
rect 47225 2329 47259 2363
rect 54033 2329 54067 2363
rect 60289 2329 60323 2363
rect 61761 2329 61795 2363
rect 66361 2329 66395 2363
rect 68293 2329 68327 2363
rect 70041 2329 70075 2363
rect 71237 2329 71271 2363
rect 74365 2329 74399 2363
rect 79701 2397 79735 2431
rect 87981 2397 88015 2431
rect 96261 2397 96295 2431
rect 78965 2329 78999 2363
rect 82829 2329 82863 2363
rect 91109 2329 91143 2363
rect 95985 2329 96019 2363
rect 98101 2329 98135 2363
rect 5825 2261 5859 2295
rect 12633 2261 12667 2295
rect 23857 2261 23891 2295
rect 29193 2261 29227 2295
rect 31125 2261 31159 2295
rect 33793 2261 33827 2295
rect 35265 2261 35299 2295
rect 36645 2261 36679 2295
rect 40509 2261 40543 2295
rect 45109 2261 45143 2295
rect 50997 2261 51031 2295
rect 55137 2261 55171 2295
rect 57713 2261 57747 2295
rect 58173 2261 58207 2295
rect 63877 2261 63911 2295
rect 65809 2261 65843 2295
rect 69121 2261 69155 2295
rect 72249 2261 72283 2295
rect 72525 2261 72559 2295
rect 76481 2261 76515 2295
rect 78689 2261 78723 2295
rect 78781 2261 78815 2295
rect 82277 2261 82311 2295
rect 87153 2261 87187 2295
rect 88349 2261 88383 2295
rect 88809 2261 88843 2295
rect 93225 2261 93259 2295
rect 93961 2261 93995 2295
rect 51549 2057 51583 2091
rect 49433 1241 49467 1275
rect 40601 1105 40635 1139
rect 31033 901 31067 935
rect 40693 1105 40727 1139
rect 40693 901 40727 935
rect 40785 901 40819 935
rect 46121 561 46155 595
rect 45017 493 45051 527
rect 44741 425 44775 459
rect 51549 1173 51583 1207
rect 58173 1309 58207 1343
rect 58173 1037 58207 1071
rect 49433 425 49467 459
rect 46121 85 46155 119
rect 31033 17 31067 51
<< metal1 >>
rect 37458 39584 37464 39636
rect 37516 39624 37522 39636
rect 80149 39627 80207 39633
rect 80149 39624 80161 39627
rect 37516 39596 80161 39624
rect 37516 39584 37522 39596
rect 80149 39593 80161 39596
rect 80195 39593 80207 39627
rect 80149 39587 80207 39593
rect 40770 39380 40776 39432
rect 40828 39420 40834 39432
rect 55490 39420 55496 39432
rect 40828 39392 55496 39420
rect 40828 39380 40834 39392
rect 55490 39380 55496 39392
rect 55548 39380 55554 39432
rect 31389 39355 31447 39361
rect 31389 39321 31401 39355
rect 31435 39352 31447 39355
rect 44726 39352 44732 39364
rect 31435 39324 44732 39352
rect 31435 39321 31447 39324
rect 31389 39315 31447 39321
rect 44726 39312 44732 39324
rect 44784 39312 44790 39364
rect 46474 39312 46480 39364
rect 46532 39352 46538 39364
rect 61102 39352 61108 39364
rect 46532 39324 61108 39352
rect 46532 39312 46538 39324
rect 61102 39312 61108 39324
rect 61160 39312 61166 39364
rect 21910 39244 21916 39296
rect 21968 39284 21974 39296
rect 89438 39284 89444 39296
rect 21968 39256 89444 39284
rect 21968 39244 21974 39256
rect 89438 39244 89444 39256
rect 89496 39244 89502 39296
rect 13722 39176 13728 39228
rect 13780 39216 13786 39228
rect 40037 39219 40095 39225
rect 40037 39216 40049 39219
rect 13780 39188 40049 39216
rect 13780 39176 13786 39188
rect 40037 39185 40049 39188
rect 40083 39185 40095 39219
rect 40037 39179 40095 39185
rect 41966 39176 41972 39228
rect 42024 39216 42030 39228
rect 63773 39219 63831 39225
rect 63773 39216 63785 39219
rect 42024 39188 63785 39216
rect 42024 39176 42030 39188
rect 63773 39185 63785 39188
rect 63819 39185 63831 39219
rect 63773 39179 63831 39185
rect 30098 39108 30104 39160
rect 30156 39148 30162 39160
rect 52365 39151 52423 39157
rect 52365 39148 52377 39151
rect 30156 39120 52377 39148
rect 30156 39108 30162 39120
rect 52365 39117 52377 39120
rect 52411 39117 52423 39151
rect 52365 39111 52423 39117
rect 54205 39151 54263 39157
rect 54205 39117 54217 39151
rect 54251 39148 54263 39151
rect 59446 39148 59452 39160
rect 54251 39120 59452 39148
rect 54251 39117 54263 39120
rect 54205 39111 54263 39117
rect 59446 39108 59452 39120
rect 59504 39108 59510 39160
rect 32858 39040 32864 39092
rect 32916 39080 32922 39092
rect 89901 39083 89959 39089
rect 89901 39080 89913 39083
rect 32916 39052 89913 39080
rect 32916 39040 32922 39052
rect 89901 39049 89913 39052
rect 89947 39049 89959 39083
rect 89901 39043 89959 39049
rect 25682 38972 25688 39024
rect 25740 39012 25746 39024
rect 84381 39015 84439 39021
rect 84381 39012 84393 39015
rect 25740 38984 84393 39012
rect 25740 38972 25746 38984
rect 84381 38981 84393 38984
rect 84427 38981 84439 39015
rect 84381 38975 84439 38981
rect 23934 38904 23940 38956
rect 23992 38944 23998 38956
rect 42337 38947 42395 38953
rect 42337 38944 42349 38947
rect 23992 38916 42349 38944
rect 23992 38904 23998 38916
rect 42337 38913 42349 38916
rect 42383 38913 42395 38947
rect 48682 38944 48688 38956
rect 42337 38907 42395 38913
rect 48424 38916 48688 38944
rect 10778 38836 10784 38888
rect 10836 38876 10842 38888
rect 38470 38876 38476 38888
rect 10836 38848 38476 38876
rect 10836 38836 10842 38848
rect 38470 38836 38476 38848
rect 38528 38836 38534 38888
rect 41693 38879 41751 38885
rect 41693 38845 41705 38879
rect 41739 38876 41751 38879
rect 48424 38876 48452 38916
rect 48682 38904 48688 38916
rect 48740 38904 48746 38956
rect 50062 38904 50068 38956
rect 50120 38944 50126 38956
rect 74261 38947 74319 38953
rect 74261 38944 74273 38947
rect 50120 38916 74273 38944
rect 50120 38904 50126 38916
rect 74261 38913 74273 38916
rect 74307 38913 74319 38947
rect 74261 38907 74319 38913
rect 41739 38848 48452 38876
rect 48501 38879 48559 38885
rect 41739 38845 41751 38848
rect 41693 38839 41751 38845
rect 48501 38845 48513 38879
rect 48547 38876 48559 38879
rect 76282 38876 76288 38888
rect 48547 38848 76288 38876
rect 48547 38845 48559 38848
rect 48501 38839 48559 38845
rect 76282 38836 76288 38848
rect 76340 38836 76346 38888
rect 19978 38768 19984 38820
rect 20036 38808 20042 38820
rect 87141 38811 87199 38817
rect 87141 38808 87153 38811
rect 20036 38780 87153 38808
rect 20036 38768 20042 38780
rect 87141 38777 87153 38780
rect 87187 38777 87199 38811
rect 87141 38771 87199 38777
rect 13906 38700 13912 38752
rect 13964 38740 13970 38752
rect 90450 38740 90456 38752
rect 13964 38712 90456 38740
rect 13964 38700 13970 38712
rect 90450 38700 90456 38712
rect 90508 38700 90514 38752
rect 5721 38675 5779 38681
rect 5721 38641 5733 38675
rect 5767 38672 5779 38675
rect 93118 38672 93124 38684
rect 5767 38644 93124 38672
rect 5767 38641 5779 38644
rect 5721 38635 5779 38641
rect 93118 38632 93124 38644
rect 93176 38632 93182 38684
rect 27982 38564 27988 38616
rect 28040 38604 28046 38616
rect 36449 38607 36507 38613
rect 36449 38604 36461 38607
rect 28040 38576 36461 38604
rect 28040 38564 28046 38576
rect 36449 38573 36461 38576
rect 36495 38573 36507 38607
rect 36449 38567 36507 38573
rect 36630 38564 36636 38616
rect 36688 38604 36694 38616
rect 68830 38604 68836 38616
rect 36688 38576 68836 38604
rect 36688 38564 36694 38576
rect 68830 38564 68836 38576
rect 68888 38564 68894 38616
rect 23290 38496 23296 38548
rect 23348 38536 23354 38548
rect 54205 38539 54263 38545
rect 54205 38536 54217 38539
rect 23348 38508 54217 38536
rect 23348 38496 23354 38508
rect 54205 38505 54217 38508
rect 54251 38505 54263 38539
rect 54205 38499 54263 38505
rect 54294 38496 54300 38548
rect 54352 38536 54358 38548
rect 56137 38539 56195 38545
rect 56137 38536 56149 38539
rect 54352 38508 56149 38536
rect 54352 38496 54358 38508
rect 56137 38505 56149 38508
rect 56183 38505 56195 38539
rect 56137 38499 56195 38505
rect 18690 38428 18696 38480
rect 18748 38468 18754 38480
rect 74810 38468 74816 38480
rect 18748 38440 74816 38468
rect 18748 38428 18754 38440
rect 74810 38428 74816 38440
rect 74868 38428 74874 38480
rect 16482 38360 16488 38412
rect 16540 38400 16546 38412
rect 75730 38400 75736 38412
rect 16540 38372 75736 38400
rect 16540 38360 16546 38372
rect 75730 38360 75736 38372
rect 75788 38360 75794 38412
rect 88978 38360 88984 38412
rect 89036 38400 89042 38412
rect 89622 38400 89628 38412
rect 89036 38372 89628 38400
rect 89036 38360 89042 38372
rect 89622 38360 89628 38372
rect 89680 38360 89686 38412
rect 26513 38335 26571 38341
rect 26513 38301 26525 38335
rect 26559 38332 26571 38335
rect 32582 38332 32588 38344
rect 26559 38304 32588 38332
rect 26559 38301 26571 38304
rect 26513 38295 26571 38301
rect 32582 38292 32588 38304
rect 32640 38292 32646 38344
rect 36449 38335 36507 38341
rect 36449 38301 36461 38335
rect 36495 38332 36507 38335
rect 90910 38332 90916 38344
rect 36495 38304 90916 38332
rect 36495 38301 36507 38304
rect 36449 38295 36507 38301
rect 90910 38292 90916 38304
rect 90968 38292 90974 38344
rect 17494 38224 17500 38276
rect 17552 38264 17558 38276
rect 81986 38264 81992 38276
rect 17552 38236 81992 38264
rect 17552 38224 17558 38236
rect 81986 38224 81992 38236
rect 82044 38224 82050 38276
rect 15378 38156 15384 38208
rect 15436 38196 15442 38208
rect 86218 38196 86224 38208
rect 15436 38168 86224 38196
rect 15436 38156 15442 38168
rect 86218 38156 86224 38168
rect 86276 38156 86282 38208
rect 4338 38088 4344 38140
rect 4396 38128 4402 38140
rect 16850 38128 16856 38140
rect 4396 38100 16856 38128
rect 4396 38088 4402 38100
rect 16850 38088 16856 38100
rect 16908 38088 16914 38140
rect 17954 38128 17960 38140
rect 16960 38100 17960 38128
rect 10410 38020 10416 38072
rect 10468 38060 10474 38072
rect 16960 38060 16988 38100
rect 17954 38088 17960 38100
rect 18012 38088 18018 38140
rect 19242 38088 19248 38140
rect 19300 38128 19306 38140
rect 93578 38128 93584 38140
rect 19300 38100 93584 38128
rect 19300 38088 19306 38100
rect 93578 38088 93584 38100
rect 93636 38088 93642 38140
rect 10468 38032 16988 38060
rect 17221 38063 17279 38069
rect 10468 38020 10474 38032
rect 17221 38029 17233 38063
rect 17267 38060 17279 38063
rect 24946 38060 24952 38072
rect 17267 38032 24952 38060
rect 17267 38029 17279 38032
rect 17221 38023 17279 38029
rect 24946 38020 24952 38032
rect 25004 38020 25010 38072
rect 26142 38020 26148 38072
rect 26200 38060 26206 38072
rect 30558 38060 30564 38072
rect 26200 38032 30564 38060
rect 26200 38020 26206 38032
rect 30558 38020 30564 38032
rect 30616 38020 30622 38072
rect 31570 38020 31576 38072
rect 31628 38060 31634 38072
rect 47854 38060 47860 38072
rect 31628 38032 47860 38060
rect 31628 38020 31634 38032
rect 47854 38020 47860 38032
rect 47912 38020 47918 38072
rect 47949 38063 48007 38069
rect 47949 38029 47961 38063
rect 47995 38060 48007 38063
rect 57790 38060 57796 38072
rect 47995 38032 57796 38060
rect 47995 38029 48007 38032
rect 47949 38023 48007 38029
rect 57790 38020 57796 38032
rect 57848 38020 57854 38072
rect 57885 38063 57943 38069
rect 57885 38029 57897 38063
rect 57931 38060 57943 38063
rect 71498 38060 71504 38072
rect 57931 38032 71504 38060
rect 57931 38029 57943 38032
rect 57885 38023 57943 38029
rect 71498 38020 71504 38032
rect 71556 38020 71562 38072
rect 15102 37952 15108 38004
rect 15160 37992 15166 38004
rect 42242 37992 42248 38004
rect 15160 37964 42248 37992
rect 15160 37952 15166 37964
rect 42242 37952 42248 37964
rect 42300 37952 42306 38004
rect 45278 37952 45284 38004
rect 45336 37992 45342 38004
rect 45336 37964 46336 37992
rect 45336 37952 45342 37964
rect 11054 37884 11060 37936
rect 11112 37924 11118 37936
rect 11112 37896 37504 37924
rect 11112 37884 11118 37896
rect 3326 37816 3332 37868
rect 3384 37856 3390 37868
rect 37366 37856 37372 37868
rect 3384 37828 37372 37856
rect 3384 37816 3390 37828
rect 37366 37816 37372 37828
rect 37424 37816 37430 37868
rect 37476 37856 37504 37896
rect 39114 37884 39120 37936
rect 39172 37924 39178 37936
rect 46308 37924 46336 37964
rect 50706 37952 50712 38004
rect 50764 37992 50770 38004
rect 70394 37992 70400 38004
rect 50764 37964 70400 37992
rect 50764 37952 50770 37964
rect 70394 37952 70400 37964
rect 70452 37952 70458 38004
rect 86034 37924 86040 37936
rect 39172 37896 46244 37924
rect 46308 37896 86040 37924
rect 39172 37884 39178 37896
rect 40310 37856 40316 37868
rect 37476 37828 40316 37856
rect 40310 37816 40316 37828
rect 40368 37816 40374 37868
rect 7006 37748 7012 37800
rect 7064 37788 7070 37800
rect 13814 37788 13820 37800
rect 7064 37760 13820 37788
rect 7064 37748 7070 37760
rect 13814 37748 13820 37760
rect 13872 37748 13878 37800
rect 14918 37748 14924 37800
rect 14976 37788 14982 37800
rect 34698 37788 34704 37800
rect 14976 37760 34704 37788
rect 14976 37748 14982 37760
rect 34698 37748 34704 37760
rect 34756 37748 34762 37800
rect 37090 37748 37096 37800
rect 37148 37788 37154 37800
rect 41690 37788 41696 37800
rect 37148 37760 41414 37788
rect 41651 37760 41696 37788
rect 37148 37748 37154 37760
rect 5718 37720 5724 37732
rect 5679 37692 5724 37720
rect 5718 37680 5724 37692
rect 5776 37680 5782 37732
rect 12342 37680 12348 37732
rect 12400 37720 12406 37732
rect 17221 37723 17279 37729
rect 17221 37720 17233 37723
rect 12400 37692 17233 37720
rect 12400 37680 12406 37692
rect 17221 37689 17233 37692
rect 17267 37689 17279 37723
rect 17221 37683 17279 37689
rect 17678 37680 17684 37732
rect 17736 37720 17742 37732
rect 25498 37720 25504 37732
rect 17736 37692 25504 37720
rect 17736 37680 17742 37692
rect 25498 37680 25504 37692
rect 25556 37680 25562 37732
rect 26510 37720 26516 37732
rect 26471 37692 26516 37720
rect 26510 37680 26516 37692
rect 26568 37680 26574 37732
rect 27062 37680 27068 37732
rect 27120 37720 27126 37732
rect 31202 37720 31208 37732
rect 27120 37692 31208 37720
rect 27120 37680 27126 37692
rect 31202 37680 31208 37692
rect 31260 37680 31266 37732
rect 31386 37720 31392 37732
rect 31347 37692 31392 37720
rect 31386 37680 31392 37692
rect 31444 37680 31450 37732
rect 40034 37720 40040 37732
rect 39995 37692 40040 37720
rect 40034 37680 40040 37692
rect 40092 37680 40098 37732
rect 41386 37720 41414 37760
rect 41690 37748 41696 37760
rect 41748 37748 41754 37800
rect 42334 37788 42340 37800
rect 42295 37760 42340 37788
rect 42334 37748 42340 37760
rect 42392 37748 42398 37800
rect 46216 37788 46244 37896
rect 86034 37884 86040 37896
rect 86092 37884 86098 37936
rect 48406 37816 48412 37868
rect 48464 37856 48470 37868
rect 56042 37856 56048 37868
rect 48464 37828 56048 37856
rect 48464 37816 48470 37828
rect 56042 37816 56048 37828
rect 56100 37816 56106 37868
rect 56137 37859 56195 37865
rect 56137 37825 56149 37859
rect 56183 37856 56195 37859
rect 66438 37856 66444 37868
rect 56183 37828 66444 37856
rect 56183 37825 56195 37828
rect 56137 37819 56195 37825
rect 66438 37816 66444 37828
rect 66496 37816 66502 37868
rect 66530 37788 66536 37800
rect 46216 37760 66536 37788
rect 66530 37748 66536 37760
rect 66588 37748 66594 37800
rect 75362 37748 75368 37800
rect 75420 37788 75426 37800
rect 96062 37788 96068 37800
rect 75420 37760 96068 37788
rect 75420 37748 75426 37760
rect 96062 37748 96068 37760
rect 96120 37748 96126 37800
rect 70118 37720 70124 37732
rect 41386 37692 70124 37720
rect 70118 37680 70124 37692
rect 70176 37680 70182 37732
rect 74258 37720 74264 37732
rect 74219 37692 74264 37720
rect 74258 37680 74264 37692
rect 74316 37680 74322 37732
rect 75454 37680 75460 37732
rect 75512 37720 75518 37732
rect 79042 37720 79048 37732
rect 75512 37692 79048 37720
rect 75512 37680 75518 37692
rect 79042 37680 79048 37692
rect 79100 37680 79106 37732
rect 81802 37680 81808 37732
rect 81860 37720 81866 37732
rect 81860 37692 85344 37720
rect 81860 37680 81866 37692
rect 4706 37612 4712 37664
rect 4764 37652 4770 37664
rect 8386 37652 8392 37664
rect 4764 37624 8392 37652
rect 4764 37612 4770 37624
rect 8386 37612 8392 37624
rect 8444 37612 8450 37664
rect 8478 37612 8484 37664
rect 8536 37652 8542 37664
rect 15930 37652 15936 37664
rect 8536 37624 15936 37652
rect 8536 37612 8542 37624
rect 15930 37612 15936 37624
rect 15988 37612 15994 37664
rect 23014 37612 23020 37664
rect 23072 37652 23078 37664
rect 36170 37652 36176 37664
rect 23072 37624 36176 37652
rect 23072 37612 23078 37624
rect 36170 37612 36176 37624
rect 36228 37612 36234 37664
rect 38930 37612 38936 37664
rect 38988 37652 38994 37664
rect 42518 37652 42524 37664
rect 38988 37624 42524 37652
rect 38988 37612 38994 37624
rect 42518 37612 42524 37624
rect 42576 37612 42582 37664
rect 43070 37612 43076 37664
rect 43128 37652 43134 37664
rect 47949 37655 48007 37661
rect 47949 37652 47961 37655
rect 43128 37624 47961 37652
rect 43128 37612 43134 37624
rect 47949 37621 47961 37624
rect 47995 37621 48007 37655
rect 48498 37652 48504 37664
rect 48459 37624 48504 37652
rect 47949 37615 48007 37621
rect 48498 37612 48504 37624
rect 48556 37612 48562 37664
rect 52362 37652 52368 37664
rect 52323 37624 52368 37652
rect 52362 37612 52368 37624
rect 52420 37612 52426 37664
rect 54938 37612 54944 37664
rect 54996 37652 55002 37664
rect 57885 37655 57943 37661
rect 57885 37652 57897 37655
rect 54996 37624 57897 37652
rect 54996 37612 55002 37624
rect 57885 37621 57897 37624
rect 57931 37621 57943 37655
rect 63770 37652 63776 37664
rect 63731 37624 63776 37652
rect 57885 37615 57943 37621
rect 63770 37612 63776 37624
rect 63828 37612 63834 37664
rect 64874 37612 64880 37664
rect 64932 37652 64938 37664
rect 76926 37652 76932 37664
rect 64932 37624 76932 37652
rect 64932 37612 64938 37624
rect 76926 37612 76932 37624
rect 76984 37612 76990 37664
rect 80149 37655 80207 37661
rect 80149 37621 80161 37655
rect 80195 37652 80207 37655
rect 80238 37652 80244 37664
rect 80195 37624 80244 37652
rect 80195 37621 80207 37624
rect 80149 37615 80207 37621
rect 80238 37612 80244 37624
rect 80296 37612 80302 37664
rect 84381 37655 84439 37661
rect 84381 37621 84393 37655
rect 84427 37652 84439 37655
rect 85206 37652 85212 37664
rect 84427 37624 85212 37652
rect 84427 37621 84439 37624
rect 84381 37615 84439 37621
rect 85206 37612 85212 37624
rect 85264 37612 85270 37664
rect 85316 37652 85344 37692
rect 86954 37680 86960 37732
rect 87012 37720 87018 37732
rect 97626 37720 97632 37732
rect 87012 37692 97632 37720
rect 87012 37680 87018 37692
rect 97626 37680 97632 37692
rect 97684 37680 97690 37732
rect 87046 37652 87052 37664
rect 85316 37624 87052 37652
rect 87046 37612 87052 37624
rect 87104 37612 87110 37664
rect 87141 37655 87199 37661
rect 87141 37621 87153 37655
rect 87187 37652 87199 37655
rect 87874 37652 87880 37664
rect 87187 37624 87880 37652
rect 87187 37621 87199 37624
rect 87141 37615 87199 37621
rect 87874 37612 87880 37624
rect 87932 37612 87938 37664
rect 89901 37655 89959 37661
rect 89901 37621 89913 37655
rect 89947 37652 89959 37655
rect 90542 37652 90548 37664
rect 89947 37624 90548 37652
rect 89947 37621 89959 37624
rect 89901 37615 89959 37621
rect 90542 37612 90548 37624
rect 90600 37612 90606 37664
rect 1104 37562 98808 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 50326 37562
rect 50378 37510 50390 37562
rect 50442 37510 50454 37562
rect 50506 37510 50518 37562
rect 50570 37510 81046 37562
rect 81098 37510 81110 37562
rect 81162 37510 81174 37562
rect 81226 37510 81238 37562
rect 81290 37510 98808 37562
rect 1104 37488 98808 37510
rect 1394 37408 1400 37460
rect 1452 37448 1458 37460
rect 4433 37451 4491 37457
rect 4433 37448 4445 37451
rect 1452 37420 4445 37448
rect 1452 37408 1458 37420
rect 4433 37417 4445 37420
rect 4479 37417 4491 37451
rect 4433 37411 4491 37417
rect 6454 37408 6460 37460
rect 6512 37448 6518 37460
rect 7837 37451 7895 37457
rect 7837 37448 7849 37451
rect 6512 37420 7849 37448
rect 6512 37408 6518 37420
rect 7837 37417 7849 37420
rect 7883 37417 7895 37451
rect 7837 37411 7895 37417
rect 8386 37408 8392 37460
rect 8444 37448 8450 37460
rect 8573 37451 8631 37457
rect 8573 37448 8585 37451
rect 8444 37420 8585 37448
rect 8444 37408 8450 37420
rect 8573 37417 8585 37420
rect 8619 37417 8631 37451
rect 8573 37411 8631 37417
rect 9493 37451 9551 37457
rect 9493 37417 9505 37451
rect 9539 37448 9551 37451
rect 10778 37448 10784 37460
rect 9539 37420 10784 37448
rect 9539 37417 9551 37420
rect 9493 37411 9551 37417
rect 382 37340 388 37392
rect 440 37380 446 37392
rect 1857 37383 1915 37389
rect 1857 37380 1869 37383
rect 440 37352 1869 37380
rect 440 37340 446 37352
rect 1857 37349 1869 37352
rect 1903 37349 1915 37383
rect 1857 37343 1915 37349
rect 3878 37340 3884 37392
rect 3936 37380 3942 37392
rect 7006 37380 7012 37392
rect 3936 37352 6914 37380
rect 6967 37352 7012 37380
rect 3936 37340 3942 37352
rect 2958 37312 2964 37324
rect 2919 37284 2964 37312
rect 2958 37272 2964 37284
rect 3016 37272 3022 37324
rect 4338 37312 4344 37324
rect 4299 37284 4344 37312
rect 4338 37272 4344 37284
rect 4396 37272 4402 37324
rect 5353 37315 5411 37321
rect 5353 37281 5365 37315
rect 5399 37312 5411 37315
rect 5442 37312 5448 37324
rect 5399 37284 5448 37312
rect 5399 37281 5411 37284
rect 5353 37275 5411 37281
rect 5442 37272 5448 37284
rect 5500 37272 5506 37324
rect 5718 37312 5724 37324
rect 5679 37284 5724 37312
rect 5718 37272 5724 37284
rect 5776 37272 5782 37324
rect 6886 37312 6914 37352
rect 7006 37340 7012 37352
rect 7064 37340 7070 37392
rect 8478 37380 8484 37392
rect 8439 37352 8484 37380
rect 8478 37340 8484 37352
rect 8536 37340 8542 37392
rect 9122 37340 9128 37392
rect 9180 37380 9186 37392
rect 9784 37389 9812 37420
rect 10778 37408 10784 37420
rect 10836 37408 10842 37460
rect 11054 37448 11060 37460
rect 11015 37420 11060 37448
rect 11054 37408 11060 37420
rect 11112 37408 11118 37460
rect 11698 37408 11704 37460
rect 11756 37448 11762 37460
rect 12437 37451 12495 37457
rect 12437 37448 12449 37451
rect 11756 37420 12449 37448
rect 11756 37408 11762 37420
rect 12437 37417 12449 37420
rect 12483 37417 12495 37451
rect 12437 37411 12495 37417
rect 14829 37451 14887 37457
rect 14829 37417 14841 37451
rect 14875 37448 14887 37451
rect 16482 37448 16488 37460
rect 14875 37420 15148 37448
rect 16443 37420 16488 37448
rect 14875 37417 14887 37420
rect 14829 37411 14887 37417
rect 15120 37392 15148 37420
rect 16482 37408 16488 37420
rect 16540 37408 16546 37460
rect 17034 37408 17040 37460
rect 17092 37448 17098 37460
rect 17773 37451 17831 37457
rect 17773 37448 17785 37451
rect 17092 37420 17785 37448
rect 17092 37408 17098 37420
rect 17773 37417 17785 37420
rect 17819 37417 17831 37451
rect 17773 37411 17831 37417
rect 17954 37408 17960 37460
rect 18012 37448 18018 37460
rect 21545 37451 21603 37457
rect 21545 37448 21557 37451
rect 18012 37420 21557 37448
rect 18012 37408 18018 37420
rect 21545 37417 21557 37420
rect 21591 37417 21603 37451
rect 21545 37411 21603 37417
rect 22278 37408 22284 37460
rect 22336 37448 22342 37460
rect 23109 37451 23167 37457
rect 23109 37448 23121 37451
rect 22336 37420 23121 37448
rect 22336 37408 22342 37420
rect 23109 37417 23121 37420
rect 23155 37417 23167 37451
rect 23109 37411 23167 37417
rect 23198 37408 23204 37460
rect 23256 37448 23262 37460
rect 23256 37420 24716 37448
rect 23256 37408 23262 37420
rect 9585 37383 9643 37389
rect 9585 37380 9597 37383
rect 9180 37352 9597 37380
rect 9180 37340 9186 37352
rect 9585 37349 9597 37352
rect 9631 37349 9643 37383
rect 9585 37343 9643 37349
rect 9769 37383 9827 37389
rect 9769 37349 9781 37383
rect 9815 37380 9827 37383
rect 11146 37380 11152 37392
rect 9815 37352 9849 37380
rect 10796 37352 11152 37380
rect 9815 37349 9827 37352
rect 9769 37343 9827 37349
rect 7193 37315 7251 37321
rect 7193 37312 7205 37315
rect 5828 37284 6040 37312
rect 6886 37284 7205 37312
rect 2314 37204 2320 37256
rect 2372 37244 2378 37256
rect 5828 37244 5856 37284
rect 2372 37216 5856 37244
rect 6012 37244 6040 37284
rect 7193 37281 7205 37284
rect 7239 37281 7251 37315
rect 7193 37275 7251 37281
rect 7745 37315 7803 37321
rect 7745 37281 7757 37315
rect 7791 37312 7803 37315
rect 10796 37312 10824 37352
rect 11146 37340 11152 37352
rect 11204 37340 11210 37392
rect 12342 37380 12348 37392
rect 12303 37352 12348 37380
rect 12342 37340 12348 37352
rect 12400 37340 12406 37392
rect 13817 37383 13875 37389
rect 13817 37349 13829 37383
rect 13863 37380 13875 37383
rect 13906 37380 13912 37392
rect 13863 37352 13912 37380
rect 13863 37349 13875 37352
rect 13817 37343 13875 37349
rect 13906 37340 13912 37352
rect 13964 37340 13970 37392
rect 14366 37340 14372 37392
rect 14424 37380 14430 37392
rect 14921 37383 14979 37389
rect 14921 37380 14933 37383
rect 14424 37352 14933 37380
rect 14424 37340 14430 37352
rect 14921 37349 14933 37352
rect 14967 37349 14979 37383
rect 15102 37380 15108 37392
rect 15063 37352 15108 37380
rect 14921 37343 14979 37349
rect 15102 37340 15108 37352
rect 15160 37340 15166 37392
rect 16114 37340 16120 37392
rect 16172 37380 16178 37392
rect 16209 37383 16267 37389
rect 16209 37380 16221 37383
rect 16172 37352 16221 37380
rect 16172 37340 16178 37352
rect 16209 37349 16221 37352
rect 16255 37349 16267 37383
rect 17678 37380 17684 37392
rect 17639 37352 17684 37380
rect 16209 37343 16267 37349
rect 17678 37340 17684 37352
rect 17736 37340 17742 37392
rect 18782 37340 18788 37392
rect 18840 37380 18846 37392
rect 18877 37383 18935 37389
rect 18877 37380 18889 37383
rect 18840 37352 18889 37380
rect 18840 37340 18846 37352
rect 18877 37349 18889 37352
rect 18923 37349 18935 37383
rect 19242 37380 19248 37392
rect 19203 37352 19248 37380
rect 18877 37343 18935 37349
rect 19242 37340 19248 37352
rect 19300 37340 19306 37392
rect 19886 37340 19892 37392
rect 19944 37380 19950 37392
rect 20533 37383 20591 37389
rect 20533 37380 20545 37383
rect 19944 37352 20545 37380
rect 19944 37340 19950 37352
rect 20533 37349 20545 37352
rect 20579 37349 20591 37383
rect 20533 37343 20591 37349
rect 21358 37340 21364 37392
rect 21416 37380 21422 37392
rect 21453 37383 21511 37389
rect 21453 37380 21465 37383
rect 21416 37352 21465 37380
rect 21416 37340 21422 37352
rect 21453 37349 21465 37352
rect 21499 37349 21511 37383
rect 23014 37380 23020 37392
rect 22975 37352 23020 37380
rect 21453 37343 21511 37349
rect 23014 37340 23020 37352
rect 23072 37340 23078 37392
rect 24026 37380 24032 37392
rect 23860 37352 24032 37380
rect 7791 37284 10824 37312
rect 10873 37315 10931 37321
rect 7791 37281 7803 37284
rect 7745 37275 7803 37281
rect 10873 37281 10885 37315
rect 10919 37312 10931 37315
rect 10962 37312 10968 37324
rect 10919 37284 10968 37312
rect 10919 37281 10931 37284
rect 10873 37275 10931 37281
rect 10962 37272 10968 37284
rect 11020 37272 11026 37324
rect 13538 37312 13544 37324
rect 13499 37284 13544 37312
rect 13538 37272 13544 37284
rect 13596 37272 13602 37324
rect 20349 37315 20407 37321
rect 13648 37284 13860 37312
rect 13648 37244 13676 37284
rect 6012 37216 13676 37244
rect 13832 37244 13860 37284
rect 20349 37281 20361 37315
rect 20395 37312 20407 37315
rect 20806 37312 20812 37324
rect 20395 37284 20812 37312
rect 20395 37281 20407 37284
rect 20349 37275 20407 37281
rect 20806 37272 20812 37284
rect 20864 37272 20870 37324
rect 23860 37321 23888 37352
rect 24026 37340 24032 37352
rect 24084 37340 24090 37392
rect 24688 37380 24716 37420
rect 24854 37408 24860 37460
rect 24912 37448 24918 37460
rect 25777 37451 25835 37457
rect 25777 37448 25789 37451
rect 24912 37420 25789 37448
rect 24912 37408 24918 37420
rect 25777 37417 25789 37420
rect 25823 37417 25835 37451
rect 25777 37411 25835 37417
rect 25866 37408 25872 37460
rect 25924 37448 25930 37460
rect 27249 37451 27307 37457
rect 27249 37448 27261 37451
rect 25924 37420 27261 37448
rect 25924 37408 25930 37420
rect 27249 37417 27261 37420
rect 27295 37417 27307 37451
rect 27249 37411 27307 37417
rect 28442 37408 28448 37460
rect 28500 37448 28506 37460
rect 29181 37451 29239 37457
rect 29181 37448 29193 37451
rect 28500 37420 29193 37448
rect 28500 37408 28506 37420
rect 29181 37417 29193 37420
rect 29227 37417 29239 37451
rect 29181 37411 29239 37417
rect 30190 37408 30196 37460
rect 30248 37448 30254 37460
rect 31113 37451 31171 37457
rect 31113 37448 31125 37451
rect 30248 37420 31125 37448
rect 30248 37408 30254 37420
rect 31113 37417 31125 37420
rect 31159 37417 31171 37451
rect 31113 37411 31171 37417
rect 31202 37408 31208 37460
rect 31260 37448 31266 37460
rect 32125 37451 32183 37457
rect 32125 37448 32137 37451
rect 31260 37420 32137 37448
rect 31260 37408 31266 37420
rect 32125 37417 32137 37420
rect 32171 37417 32183 37451
rect 32125 37411 32183 37417
rect 32766 37408 32772 37460
rect 32824 37448 32830 37460
rect 33781 37451 33839 37457
rect 33781 37448 33793 37451
rect 32824 37420 33793 37448
rect 32824 37408 32830 37420
rect 33781 37417 33793 37420
rect 33827 37417 33839 37451
rect 34698 37448 34704 37460
rect 34659 37420 34704 37448
rect 33781 37411 33839 37417
rect 34698 37408 34704 37420
rect 34756 37408 34762 37460
rect 35434 37408 35440 37460
rect 35492 37448 35498 37460
rect 36449 37451 36507 37457
rect 36449 37448 36461 37451
rect 35492 37420 36461 37448
rect 35492 37408 35498 37420
rect 36449 37417 36461 37420
rect 36495 37417 36507 37451
rect 37366 37448 37372 37460
rect 37327 37420 37372 37448
rect 36449 37411 36507 37417
rect 37366 37408 37372 37420
rect 37424 37408 37430 37460
rect 38102 37408 38108 37460
rect 38160 37448 38166 37460
rect 39117 37451 39175 37457
rect 39117 37448 39129 37451
rect 38160 37420 39129 37448
rect 38160 37408 38166 37420
rect 39117 37417 39129 37420
rect 39163 37417 39175 37451
rect 40034 37448 40040 37460
rect 39995 37420 40040 37448
rect 39117 37411 39175 37417
rect 40034 37408 40040 37420
rect 40092 37408 40098 37460
rect 40678 37408 40684 37460
rect 40736 37448 40742 37460
rect 41785 37451 41843 37457
rect 41785 37448 41797 37451
rect 40736 37420 41797 37448
rect 40736 37408 40742 37420
rect 41785 37417 41797 37420
rect 41831 37417 41843 37451
rect 42518 37448 42524 37460
rect 42479 37420 42524 37448
rect 41785 37411 41843 37417
rect 42518 37408 42524 37420
rect 42576 37408 42582 37460
rect 44453 37451 44511 37457
rect 44453 37448 44465 37451
rect 43088 37420 44465 37448
rect 26329 37383 26387 37389
rect 26329 37380 26341 37383
rect 24688 37352 26341 37380
rect 26329 37349 26341 37352
rect 26375 37349 26387 37383
rect 26510 37380 26516 37392
rect 26471 37352 26516 37380
rect 26329 37343 26387 37349
rect 26510 37340 26516 37352
rect 26568 37340 26574 37392
rect 27522 37340 27528 37392
rect 27580 37380 27586 37392
rect 28537 37383 28595 37389
rect 28537 37380 28549 37383
rect 27580 37352 28549 37380
rect 27580 37340 27586 37352
rect 28537 37349 28549 37352
rect 28583 37349 28595 37383
rect 28537 37343 28595 37349
rect 30009 37383 30067 37389
rect 30009 37349 30021 37383
rect 30055 37380 30067 37383
rect 30926 37380 30932 37392
rect 30055 37352 30932 37380
rect 30055 37349 30067 37352
rect 30009 37343 30067 37349
rect 30926 37340 30932 37352
rect 30984 37340 30990 37392
rect 31021 37383 31079 37389
rect 31021 37349 31033 37383
rect 31067 37380 31079 37383
rect 31386 37380 31392 37392
rect 31067 37352 31392 37380
rect 31067 37349 31079 37352
rect 31021 37343 31079 37349
rect 31386 37340 31392 37352
rect 31444 37340 31450 37392
rect 31938 37340 31944 37392
rect 31996 37380 32002 37392
rect 32033 37383 32091 37389
rect 32033 37380 32045 37383
rect 31996 37352 32045 37380
rect 31996 37340 32002 37352
rect 32033 37349 32045 37352
rect 32079 37349 32091 37383
rect 32033 37343 32091 37349
rect 34514 37340 34520 37392
rect 34572 37380 34578 37392
rect 34609 37383 34667 37389
rect 34609 37380 34621 37383
rect 34572 37352 34621 37380
rect 34572 37340 34578 37352
rect 34609 37349 34621 37352
rect 34655 37349 34667 37383
rect 34609 37343 34667 37349
rect 36357 37383 36415 37389
rect 36357 37349 36369 37383
rect 36403 37380 36415 37383
rect 41322 37380 41328 37392
rect 36403 37352 41328 37380
rect 36403 37349 36415 37352
rect 36357 37343 36415 37349
rect 41322 37340 41328 37352
rect 41380 37340 41386 37392
rect 41598 37340 41604 37392
rect 41656 37380 41662 37392
rect 43088 37380 43116 37420
rect 44453 37417 44465 37420
rect 44499 37417 44511 37451
rect 45278 37448 45284 37460
rect 45239 37420 45284 37448
rect 44453 37411 44511 37417
rect 45278 37408 45284 37420
rect 45336 37408 45342 37460
rect 45922 37408 45928 37460
rect 45980 37448 45986 37460
rect 47121 37451 47179 37457
rect 47121 37448 47133 37451
rect 45980 37420 47133 37448
rect 45980 37408 45986 37420
rect 47121 37417 47133 37420
rect 47167 37417 47179 37451
rect 47854 37448 47860 37460
rect 47815 37420 47860 37448
rect 47121 37411 47179 37417
rect 47854 37408 47860 37420
rect 47912 37408 47918 37460
rect 48590 37448 48596 37460
rect 48551 37420 48596 37448
rect 48590 37408 48596 37420
rect 48648 37408 48654 37460
rect 50525 37451 50583 37457
rect 50525 37417 50537 37451
rect 50571 37448 50583 37451
rect 50706 37448 50712 37460
rect 50571 37420 50712 37448
rect 50571 37417 50583 37420
rect 50525 37411 50583 37417
rect 50706 37408 50712 37420
rect 50764 37408 50770 37460
rect 51258 37448 51264 37460
rect 51219 37420 51264 37448
rect 51258 37408 51264 37420
rect 51316 37408 51322 37460
rect 52086 37408 52092 37460
rect 52144 37448 52150 37460
rect 55861 37451 55919 37457
rect 55861 37448 55873 37451
rect 52144 37420 55873 37448
rect 52144 37408 52150 37420
rect 55861 37417 55873 37420
rect 55907 37417 55919 37451
rect 55861 37411 55919 37417
rect 56502 37408 56508 37460
rect 56560 37448 56566 37460
rect 56597 37451 56655 37457
rect 56597 37448 56609 37451
rect 56560 37420 56609 37448
rect 56560 37408 56566 37420
rect 56597 37417 56609 37420
rect 56643 37417 56655 37451
rect 57790 37448 57796 37460
rect 57751 37420 57796 37448
rect 56597 37411 56655 37417
rect 57790 37408 57796 37420
rect 57848 37408 57854 37460
rect 59078 37408 59084 37460
rect 59136 37448 59142 37460
rect 61749 37451 61807 37457
rect 61749 37448 61761 37451
rect 59136 37420 61761 37448
rect 59136 37408 59142 37420
rect 61749 37417 61761 37420
rect 61795 37417 61807 37451
rect 61749 37411 61807 37417
rect 61838 37408 61844 37460
rect 61896 37448 61902 37460
rect 64417 37451 64475 37457
rect 64417 37448 64429 37451
rect 61896 37420 64429 37448
rect 61896 37408 61902 37420
rect 64417 37417 64429 37420
rect 64463 37417 64475 37451
rect 64417 37411 64475 37417
rect 64506 37408 64512 37460
rect 64564 37448 64570 37460
rect 67085 37451 67143 37457
rect 67085 37448 67097 37451
rect 64564 37420 67097 37448
rect 64564 37408 64570 37420
rect 67085 37417 67097 37420
rect 67131 37417 67143 37451
rect 67085 37411 67143 37417
rect 67174 37408 67180 37460
rect 67232 37448 67238 37460
rect 69661 37451 69719 37457
rect 69661 37448 69673 37451
rect 67232 37420 69673 37448
rect 67232 37408 67238 37420
rect 69661 37417 69673 37420
rect 69707 37417 69719 37451
rect 69661 37411 69719 37417
rect 69750 37408 69756 37460
rect 69808 37448 69814 37460
rect 69808 37420 71728 37448
rect 69808 37408 69814 37420
rect 43346 37380 43352 37392
rect 41656 37352 43116 37380
rect 43307 37352 43352 37380
rect 41656 37340 41662 37352
rect 43346 37340 43352 37352
rect 43404 37340 43410 37392
rect 47670 37340 47676 37392
rect 47728 37380 47734 37392
rect 47765 37383 47823 37389
rect 47765 37380 47777 37383
rect 47728 37352 47777 37380
rect 47728 37340 47734 37352
rect 47765 37349 47777 37352
rect 47811 37349 47823 37383
rect 48498 37380 48504 37392
rect 48459 37352 48504 37380
rect 47765 37343 47823 37349
rect 48498 37340 48504 37352
rect 48556 37340 48562 37392
rect 49418 37340 49424 37392
rect 49476 37380 49482 37392
rect 49476 37352 50108 37380
rect 49476 37340 49482 37352
rect 23845 37315 23903 37321
rect 23845 37281 23857 37315
rect 23891 37281 23903 37315
rect 24118 37312 24124 37324
rect 24079 37284 24124 37312
rect 23845 37275 23903 37281
rect 24118 37272 24124 37284
rect 24176 37272 24182 37324
rect 25685 37315 25743 37321
rect 25685 37281 25697 37315
rect 25731 37312 25743 37315
rect 26142 37312 26148 37324
rect 25731 37284 26148 37312
rect 25731 37281 25743 37284
rect 25685 37275 25743 37281
rect 26142 37272 26148 37284
rect 26200 37272 26206 37324
rect 26237 37315 26295 37321
rect 26237 37281 26249 37315
rect 26283 37312 26295 37315
rect 26528 37312 26556 37340
rect 27154 37312 27160 37324
rect 26283 37284 26556 37312
rect 27115 37284 27160 37312
rect 26283 37281 26295 37284
rect 26237 37275 26295 37281
rect 27154 37272 27160 37284
rect 27212 37272 27218 37324
rect 28350 37312 28356 37324
rect 28311 37284 28356 37312
rect 28350 37272 28356 37284
rect 28408 37272 28414 37324
rect 29089 37315 29147 37321
rect 29089 37281 29101 37315
rect 29135 37312 29147 37315
rect 29638 37312 29644 37324
rect 29135 37284 29644 37312
rect 29135 37281 29147 37284
rect 29089 37275 29147 37281
rect 29638 37272 29644 37284
rect 29696 37272 29702 37324
rect 29825 37315 29883 37321
rect 29825 37281 29837 37315
rect 29871 37312 29883 37315
rect 31478 37312 31484 37324
rect 29871 37284 31484 37312
rect 29871 37281 29883 37284
rect 29825 37275 29883 37281
rect 31478 37272 31484 37284
rect 31536 37272 31542 37324
rect 33689 37315 33747 37321
rect 33689 37281 33701 37315
rect 33735 37312 33747 37315
rect 34054 37312 34060 37324
rect 33735 37284 34060 37312
rect 33735 37281 33747 37284
rect 33689 37275 33747 37281
rect 34054 37272 34060 37284
rect 34112 37272 34118 37324
rect 36078 37272 36084 37324
rect 36136 37312 36142 37324
rect 36630 37312 36636 37324
rect 36136 37284 36636 37312
rect 36136 37272 36142 37284
rect 36630 37272 36636 37284
rect 36688 37272 36694 37324
rect 37182 37312 37188 37324
rect 37143 37284 37188 37312
rect 37182 37272 37188 37284
rect 37240 37272 37246 37324
rect 38654 37272 38660 37324
rect 38712 37312 38718 37324
rect 39025 37315 39083 37321
rect 39025 37312 39037 37315
rect 38712 37284 39037 37312
rect 38712 37272 38718 37284
rect 39025 37281 39037 37284
rect 39071 37281 39083 37315
rect 39850 37312 39856 37324
rect 39811 37284 39856 37312
rect 39025 37275 39083 37281
rect 39850 37272 39856 37284
rect 39908 37272 39914 37324
rect 41690 37312 41696 37324
rect 41651 37284 41696 37312
rect 41690 37272 41696 37284
rect 41748 37272 41754 37324
rect 42334 37272 42340 37324
rect 42392 37312 42398 37324
rect 42429 37315 42487 37321
rect 42429 37312 42441 37315
rect 42392 37284 42441 37312
rect 42392 37272 42398 37284
rect 42429 37281 42441 37284
rect 42475 37281 42487 37315
rect 42429 37275 42487 37281
rect 42886 37272 42892 37324
rect 42944 37312 42950 37324
rect 43165 37315 43223 37321
rect 43165 37312 43177 37315
rect 42944 37284 43177 37312
rect 42944 37272 42950 37284
rect 43165 37281 43177 37284
rect 43211 37281 43223 37315
rect 44358 37312 44364 37324
rect 44319 37284 44364 37312
rect 43165 37275 43223 37281
rect 44358 37272 44364 37284
rect 44416 37272 44422 37324
rect 45094 37312 45100 37324
rect 45055 37284 45100 37312
rect 45094 37272 45100 37284
rect 45152 37272 45158 37324
rect 47029 37315 47087 37321
rect 47029 37281 47041 37315
rect 47075 37312 47087 37315
rect 47946 37312 47952 37324
rect 47075 37284 47952 37312
rect 47075 37281 47087 37284
rect 47029 37275 47087 37281
rect 47946 37272 47952 37284
rect 48004 37272 48010 37324
rect 49694 37312 49700 37324
rect 49655 37284 49700 37312
rect 49694 37272 49700 37284
rect 49752 37272 49758 37324
rect 49878 37312 49884 37324
rect 49839 37284 49884 37312
rect 49878 37272 49884 37284
rect 49936 37272 49942 37324
rect 50080 37312 50108 37352
rect 50154 37340 50160 37392
rect 50212 37380 50218 37392
rect 50433 37383 50491 37389
rect 50433 37380 50445 37383
rect 50212 37352 50445 37380
rect 50212 37340 50218 37352
rect 50433 37349 50445 37352
rect 50479 37349 50491 37383
rect 52549 37383 52607 37389
rect 52549 37380 52561 37383
rect 50433 37343 50491 37349
rect 51046 37352 52561 37380
rect 51046 37312 51074 37352
rect 52549 37349 52561 37352
rect 52595 37349 52607 37383
rect 52549 37343 52607 37349
rect 53006 37340 53012 37392
rect 53064 37380 53070 37392
rect 53101 37383 53159 37389
rect 53101 37380 53113 37383
rect 53064 37352 53113 37380
rect 53064 37340 53070 37352
rect 53101 37349 53113 37352
rect 53147 37349 53159 37383
rect 53101 37343 53159 37349
rect 53834 37340 53840 37392
rect 53892 37380 53898 37392
rect 55217 37383 55275 37389
rect 55217 37380 55229 37383
rect 53892 37352 55229 37380
rect 53892 37340 53898 37352
rect 55217 37349 55229 37352
rect 55263 37349 55275 37383
rect 55217 37343 55275 37349
rect 55398 37340 55404 37392
rect 55456 37380 55462 37392
rect 57701 37383 57759 37389
rect 55456 37352 56548 37380
rect 55456 37340 55462 37352
rect 51166 37312 51172 37324
rect 50080 37284 51074 37312
rect 51127 37284 51172 37312
rect 51166 37272 51172 37284
rect 51224 37272 51230 37324
rect 52362 37312 52368 37324
rect 52323 37284 52368 37312
rect 52362 37272 52368 37284
rect 52420 37272 52426 37324
rect 53466 37312 53472 37324
rect 53427 37284 53472 37312
rect 53466 37272 53472 37284
rect 53524 37272 53530 37324
rect 54662 37272 54668 37324
rect 54720 37312 54726 37324
rect 55033 37315 55091 37321
rect 55033 37312 55045 37315
rect 54720 37284 55045 37312
rect 54720 37272 54726 37284
rect 55033 37281 55045 37284
rect 55079 37281 55091 37315
rect 55033 37275 55091 37281
rect 55674 37272 55680 37324
rect 55732 37312 55738 37324
rect 56520 37321 56548 37352
rect 57701 37349 57713 37383
rect 57747 37380 57759 37383
rect 58250 37380 58256 37392
rect 57747 37352 58256 37380
rect 57747 37349 57759 37352
rect 57701 37343 57759 37349
rect 58250 37340 58256 37352
rect 58308 37340 58314 37392
rect 60826 37340 60832 37392
rect 60884 37380 60890 37392
rect 60921 37383 60979 37389
rect 60921 37380 60933 37383
rect 60884 37352 60933 37380
rect 60884 37340 60890 37352
rect 60921 37349 60933 37352
rect 60967 37349 60979 37383
rect 61102 37380 61108 37392
rect 61063 37352 61108 37380
rect 60921 37343 60979 37349
rect 61102 37340 61108 37352
rect 61160 37340 61166 37392
rect 63494 37340 63500 37392
rect 63552 37380 63558 37392
rect 63589 37383 63647 37389
rect 63589 37380 63601 37383
rect 63552 37352 63601 37380
rect 63552 37340 63558 37352
rect 63589 37349 63601 37352
rect 63635 37349 63647 37383
rect 63770 37380 63776 37392
rect 63731 37352 63776 37380
rect 63589 37343 63647 37349
rect 63770 37340 63776 37352
rect 63828 37340 63834 37392
rect 66162 37340 66168 37392
rect 66220 37380 66226 37392
rect 66257 37383 66315 37389
rect 66257 37380 66269 37383
rect 66220 37352 66269 37380
rect 66220 37340 66226 37352
rect 66257 37349 66269 37352
rect 66303 37349 66315 37383
rect 66438 37380 66444 37392
rect 66399 37352 66444 37380
rect 66257 37343 66315 37349
rect 66438 37340 66444 37352
rect 66496 37340 66502 37392
rect 71406 37340 71412 37392
rect 71464 37380 71470 37392
rect 71501 37383 71559 37389
rect 71501 37380 71513 37383
rect 71464 37352 71513 37380
rect 71464 37340 71470 37352
rect 71501 37349 71513 37352
rect 71547 37349 71559 37383
rect 71700 37380 71728 37420
rect 77570 37408 77576 37460
rect 77628 37448 77634 37460
rect 79137 37451 79195 37457
rect 79137 37448 79149 37451
rect 77628 37420 79149 37448
rect 77628 37408 77634 37420
rect 79137 37417 79149 37420
rect 79183 37417 79195 37451
rect 79137 37411 79195 37417
rect 80146 37408 80152 37460
rect 80204 37448 80210 37460
rect 80333 37451 80391 37457
rect 80333 37448 80345 37451
rect 80204 37420 80345 37448
rect 80204 37408 80210 37420
rect 80333 37417 80345 37420
rect 80379 37417 80391 37451
rect 80333 37411 80391 37417
rect 81342 37408 81348 37460
rect 81400 37448 81406 37460
rect 81400 37420 82584 37448
rect 81400 37408 81406 37420
rect 72421 37383 72479 37389
rect 72421 37380 72433 37383
rect 71700 37352 72433 37380
rect 71501 37343 71559 37349
rect 72421 37349 72433 37352
rect 72467 37349 72479 37383
rect 72421 37343 72479 37349
rect 73982 37340 73988 37392
rect 74040 37380 74046 37392
rect 74077 37383 74135 37389
rect 74077 37380 74089 37383
rect 74040 37352 74089 37380
rect 74040 37340 74046 37352
rect 74077 37349 74089 37352
rect 74123 37349 74135 37383
rect 74997 37383 75055 37389
rect 74997 37380 75009 37383
rect 74077 37343 74135 37349
rect 74184 37352 75009 37380
rect 55769 37315 55827 37321
rect 55769 37312 55781 37315
rect 55732 37284 55781 37312
rect 55732 37272 55738 37284
rect 55769 37281 55781 37284
rect 55815 37281 55827 37315
rect 55769 37275 55827 37281
rect 56505 37315 56563 37321
rect 56505 37281 56517 37315
rect 56551 37281 56563 37315
rect 58434 37312 58440 37324
rect 58395 37284 58440 37312
rect 56505 37275 56563 37281
rect 58434 37272 58440 37284
rect 58492 37272 58498 37324
rect 58894 37312 58900 37324
rect 58855 37284 58900 37312
rect 58894 37272 58900 37284
rect 58952 37272 58958 37324
rect 61654 37312 61660 37324
rect 61615 37284 61660 37312
rect 61654 37272 61660 37284
rect 61712 37272 61718 37324
rect 64322 37312 64328 37324
rect 64283 37284 64328 37312
rect 64322 37272 64328 37284
rect 64380 37272 64386 37324
rect 66990 37312 66996 37324
rect 66951 37284 66996 37312
rect 66990 37272 66996 37284
rect 67048 37272 67054 37324
rect 68738 37312 68744 37324
rect 68699 37284 68744 37312
rect 68738 37272 68744 37284
rect 68796 37272 68802 37324
rect 68848 37284 69060 37312
rect 22094 37244 22100 37256
rect 13832 37216 22100 37244
rect 2372 37204 2378 37216
rect 22094 37204 22100 37216
rect 22152 37204 22158 37256
rect 40957 37247 41015 37253
rect 40957 37244 40969 37247
rect 22204 37216 40969 37244
rect 1673 37179 1731 37185
rect 1673 37145 1685 37179
rect 1719 37176 1731 37179
rect 2133 37179 2191 37185
rect 2133 37176 2145 37179
rect 1719 37148 2145 37176
rect 1719 37145 1731 37148
rect 1673 37139 1731 37145
rect 2133 37145 2145 37148
rect 2179 37176 2191 37179
rect 2409 37179 2467 37185
rect 2409 37176 2421 37179
rect 2179 37148 2421 37176
rect 2179 37145 2191 37148
rect 2133 37139 2191 37145
rect 2409 37145 2421 37148
rect 2455 37176 2467 37179
rect 22204 37176 22232 37216
rect 40957 37213 40969 37216
rect 41003 37213 41015 37247
rect 40957 37207 41015 37213
rect 41046 37204 41052 37256
rect 41104 37244 41110 37256
rect 64966 37244 64972 37256
rect 41104 37216 64972 37244
rect 41104 37204 41110 37216
rect 64966 37204 64972 37216
rect 65024 37204 65030 37256
rect 65058 37204 65064 37256
rect 65116 37244 65122 37256
rect 68554 37244 68560 37256
rect 65116 37216 68560 37244
rect 65116 37204 65122 37216
rect 68554 37204 68560 37216
rect 68612 37204 68618 37256
rect 68848 37244 68876 37284
rect 68756 37216 68876 37244
rect 2455 37148 22232 37176
rect 2455 37145 2467 37148
rect 2409 37139 2467 37145
rect 28534 37136 28540 37188
rect 28592 37176 28598 37188
rect 68756 37176 68784 37216
rect 68922 37176 68928 37188
rect 28592 37148 68784 37176
rect 68883 37148 68928 37176
rect 28592 37136 28598 37148
rect 68922 37136 68928 37148
rect 68980 37136 68986 37188
rect 69032 37176 69060 37284
rect 69474 37272 69480 37324
rect 69532 37312 69538 37324
rect 69569 37315 69627 37321
rect 69569 37312 69581 37315
rect 69532 37284 69581 37312
rect 69532 37272 69538 37284
rect 69569 37281 69581 37284
rect 69615 37281 69627 37315
rect 69569 37275 69627 37281
rect 71682 37272 71688 37324
rect 71740 37312 71746 37324
rect 72237 37315 72295 37321
rect 72237 37312 72249 37315
rect 71740 37284 72249 37312
rect 71740 37272 71746 37284
rect 72237 37281 72249 37284
rect 72283 37281 72295 37315
rect 72237 37275 72295 37281
rect 72326 37272 72332 37324
rect 72384 37312 72390 37324
rect 74184 37312 74212 37352
rect 74997 37349 75009 37352
rect 75043 37349 75055 37383
rect 74997 37343 75055 37349
rect 76650 37340 76656 37392
rect 76708 37380 76714 37392
rect 76745 37383 76803 37389
rect 76745 37380 76757 37383
rect 76708 37352 76757 37380
rect 76708 37340 76714 37352
rect 76745 37349 76757 37352
rect 76791 37349 76803 37383
rect 76745 37343 76803 37349
rect 76834 37340 76840 37392
rect 76892 37380 76898 37392
rect 81802 37380 81808 37392
rect 76892 37352 81808 37380
rect 76892 37340 76898 37352
rect 81802 37340 81808 37352
rect 81860 37340 81866 37392
rect 81894 37340 81900 37392
rect 81952 37380 81958 37392
rect 81989 37383 82047 37389
rect 81989 37380 82001 37383
rect 81952 37352 82001 37380
rect 81952 37340 81958 37352
rect 81989 37349 82001 37352
rect 82035 37349 82047 37383
rect 82556 37380 82584 37420
rect 82814 37408 82820 37460
rect 82872 37448 82878 37460
rect 83001 37451 83059 37457
rect 83001 37448 83013 37451
rect 82872 37420 83013 37448
rect 82872 37408 82878 37420
rect 83001 37417 83013 37420
rect 83047 37417 83059 37451
rect 83001 37411 83059 37417
rect 83642 37408 83648 37460
rect 83700 37448 83706 37460
rect 83700 37420 86264 37448
rect 83700 37408 83706 37420
rect 84565 37383 84623 37389
rect 84565 37380 84577 37383
rect 82556 37352 84577 37380
rect 81989 37343 82047 37349
rect 84565 37349 84577 37352
rect 84611 37349 84623 37383
rect 85206 37380 85212 37392
rect 85167 37352 85212 37380
rect 84565 37343 84623 37349
rect 85206 37340 85212 37352
rect 85264 37340 85270 37392
rect 85390 37380 85396 37392
rect 85351 37352 85396 37380
rect 85390 37340 85396 37352
rect 85448 37340 85454 37392
rect 85482 37340 85488 37392
rect 85540 37380 85546 37392
rect 86236 37380 86264 37420
rect 86310 37408 86316 37460
rect 86368 37448 86374 37460
rect 86368 37420 89668 37448
rect 86368 37408 86374 37420
rect 87233 37383 87291 37389
rect 87233 37380 87245 37383
rect 85540 37352 85712 37380
rect 86236 37352 87245 37380
rect 85540 37340 85546 37352
rect 72384 37284 74212 37312
rect 72384 37272 72390 37284
rect 74258 37272 74264 37324
rect 74316 37312 74322 37324
rect 74316 37284 74361 37312
rect 74316 37272 74322 37284
rect 74718 37272 74724 37324
rect 74776 37312 74782 37324
rect 74813 37315 74871 37321
rect 74813 37312 74825 37315
rect 74776 37284 74825 37312
rect 74776 37272 74782 37284
rect 74813 37281 74825 37284
rect 74859 37281 74871 37315
rect 74813 37275 74871 37281
rect 74902 37272 74908 37324
rect 74960 37312 74966 37324
rect 77478 37312 77484 37324
rect 74960 37284 77340 37312
rect 77439 37284 77484 37312
rect 74960 37272 74966 37284
rect 70670 37204 70676 37256
rect 70728 37244 70734 37256
rect 73246 37244 73252 37256
rect 70728 37216 73252 37244
rect 70728 37204 70734 37216
rect 73246 37204 73252 37216
rect 73304 37204 73310 37256
rect 73522 37204 73528 37256
rect 73580 37244 73586 37256
rect 76190 37244 76196 37256
rect 73580 37216 76196 37244
rect 73580 37204 73586 37216
rect 76190 37204 76196 37216
rect 76248 37204 76254 37256
rect 76926 37244 76932 37256
rect 76887 37216 76932 37244
rect 76926 37204 76932 37216
rect 76984 37204 76990 37256
rect 77312 37244 77340 37284
rect 77478 37272 77484 37284
rect 77536 37272 77542 37324
rect 77665 37315 77723 37321
rect 77665 37312 77677 37315
rect 77588 37284 77677 37312
rect 77588 37244 77616 37284
rect 77665 37281 77677 37284
rect 77711 37281 77723 37315
rect 79042 37312 79048 37324
rect 79003 37284 79048 37312
rect 77665 37275 77723 37281
rect 79042 37272 79048 37284
rect 79100 37272 79106 37324
rect 80238 37312 80244 37324
rect 80199 37284 80244 37312
rect 80238 37272 80244 37284
rect 80296 37272 80302 37324
rect 81434 37272 81440 37324
rect 81492 37312 81498 37324
rect 82173 37315 82231 37321
rect 82173 37312 82185 37315
rect 81492 37284 82185 37312
rect 81492 37272 81498 37284
rect 82173 37281 82185 37284
rect 82219 37281 82231 37315
rect 82906 37312 82912 37324
rect 82867 37284 82912 37312
rect 82173 37275 82231 37281
rect 82906 37272 82912 37284
rect 82964 37272 82970 37324
rect 84194 37272 84200 37324
rect 84252 37312 84258 37324
rect 84381 37315 84439 37321
rect 84381 37312 84393 37315
rect 84252 37284 84393 37312
rect 84252 37272 84258 37284
rect 84381 37281 84393 37284
rect 84427 37281 84439 37315
rect 85224 37312 85252 37340
rect 85577 37315 85635 37321
rect 85577 37312 85589 37315
rect 85224 37284 85589 37312
rect 84381 37275 84439 37281
rect 85577 37281 85589 37284
rect 85623 37281 85635 37315
rect 85684 37312 85712 37352
rect 87233 37349 87245 37352
rect 87279 37349 87291 37383
rect 87874 37380 87880 37392
rect 87835 37352 87880 37380
rect 87233 37343 87291 37349
rect 87874 37340 87880 37352
rect 87932 37340 87938 37392
rect 88058 37380 88064 37392
rect 88019 37352 88064 37380
rect 88058 37340 88064 37352
rect 88116 37340 88122 37392
rect 89438 37380 89444 37392
rect 89399 37352 89444 37380
rect 89438 37340 89444 37352
rect 89496 37340 89502 37392
rect 89640 37389 89668 37420
rect 89714 37408 89720 37460
rect 89772 37448 89778 37460
rect 92385 37451 92443 37457
rect 92385 37448 92397 37451
rect 89772 37420 92397 37448
rect 89772 37408 89778 37420
rect 92385 37417 92397 37420
rect 92431 37417 92443 37451
rect 92385 37411 92443 37417
rect 95970 37408 95976 37460
rect 96028 37448 96034 37460
rect 96157 37451 96215 37457
rect 96157 37448 96169 37451
rect 96028 37420 96169 37448
rect 96028 37408 96034 37420
rect 96157 37417 96169 37420
rect 96203 37417 96215 37451
rect 97626 37448 97632 37460
rect 97587 37420 97632 37448
rect 96157 37411 96215 37417
rect 97626 37408 97632 37420
rect 97684 37408 97690 37460
rect 89625 37383 89683 37389
rect 89625 37349 89637 37383
rect 89671 37349 89683 37383
rect 90542 37380 90548 37392
rect 90503 37352 90548 37380
rect 89625 37343 89683 37349
rect 90542 37340 90548 37352
rect 90600 37340 90606 37392
rect 90726 37380 90732 37392
rect 90687 37352 90732 37380
rect 90726 37340 90732 37352
rect 90784 37340 90790 37392
rect 93302 37380 93308 37392
rect 93263 37352 93308 37380
rect 93302 37340 93308 37352
rect 93360 37340 93366 37392
rect 96062 37380 96068 37392
rect 96023 37352 96068 37380
rect 96062 37340 96068 37352
rect 96120 37340 96126 37392
rect 97644 37380 97672 37408
rect 97905 37383 97963 37389
rect 97905 37380 97917 37383
rect 97644 37352 97917 37380
rect 97905 37349 97917 37352
rect 97951 37349 97963 37383
rect 97905 37343 97963 37349
rect 98089 37383 98147 37389
rect 98089 37349 98101 37383
rect 98135 37380 98147 37383
rect 98546 37380 98552 37392
rect 98135 37352 98552 37380
rect 98135 37349 98147 37352
rect 98089 37343 98147 37349
rect 87049 37315 87107 37321
rect 87049 37312 87061 37315
rect 85684 37284 87061 37312
rect 85577 37275 85635 37281
rect 87049 37281 87061 37284
rect 87095 37281 87107 37315
rect 87892 37312 87920 37340
rect 88245 37315 88303 37321
rect 88245 37312 88257 37315
rect 87892 37284 88257 37312
rect 87049 37275 87107 37281
rect 88245 37281 88257 37284
rect 88291 37281 88303 37315
rect 89456 37312 89484 37340
rect 89809 37315 89867 37321
rect 89809 37312 89821 37315
rect 89456 37284 89821 37312
rect 88245 37275 88303 37281
rect 89809 37281 89821 37284
rect 89855 37281 89867 37315
rect 90560 37312 90588 37340
rect 90913 37315 90971 37321
rect 90913 37312 90925 37315
rect 90560 37284 90925 37312
rect 89809 37275 89867 37281
rect 90913 37281 90925 37284
rect 90959 37312 90971 37315
rect 91097 37315 91155 37321
rect 91097 37312 91109 37315
rect 90959 37284 91109 37312
rect 90959 37281 90971 37284
rect 90913 37275 90971 37281
rect 91097 37281 91109 37284
rect 91143 37281 91155 37315
rect 92477 37315 92535 37321
rect 92477 37312 92489 37315
rect 91097 37275 91155 37281
rect 92124 37284 92489 37312
rect 77312 37216 77616 37244
rect 92124 37185 92152 37284
rect 92477 37281 92489 37284
rect 92523 37312 92535 37315
rect 92661 37315 92719 37321
rect 92661 37312 92673 37315
rect 92523 37284 92673 37312
rect 92523 37281 92535 37284
rect 92477 37275 92535 37281
rect 92661 37281 92673 37284
rect 92707 37281 92719 37315
rect 92661 37275 92719 37281
rect 93213 37315 93271 37321
rect 93213 37281 93225 37315
rect 93259 37312 93271 37315
rect 93486 37312 93492 37324
rect 93259 37284 93492 37312
rect 93259 37281 93271 37284
rect 93213 37275 93271 37281
rect 93486 37272 93492 37284
rect 93544 37272 93550 37324
rect 94130 37272 94136 37324
rect 94188 37312 94194 37324
rect 95053 37315 95111 37321
rect 95053 37312 95065 37315
rect 94188 37284 95065 37312
rect 94188 37272 94194 37284
rect 95053 37281 95065 37284
rect 95099 37281 95111 37315
rect 95234 37312 95240 37324
rect 95195 37284 95240 37312
rect 95053 37275 95111 37281
rect 95234 37272 95240 37284
rect 95292 37272 95298 37324
rect 97920 37312 97948 37343
rect 98546 37340 98552 37352
rect 98604 37340 98610 37392
rect 98181 37315 98239 37321
rect 98181 37312 98193 37315
rect 97920 37284 98193 37312
rect 98181 37281 98193 37284
rect 98227 37281 98239 37315
rect 98181 37275 98239 37281
rect 92109 37179 92167 37185
rect 92109 37176 92121 37179
rect 69032 37148 89576 37176
rect 3142 37108 3148 37120
rect 3103 37080 3148 37108
rect 3142 37068 3148 37080
rect 3200 37068 3206 37120
rect 23474 37068 23480 37120
rect 23532 37108 23538 37120
rect 29638 37108 29644 37120
rect 23532 37080 29644 37108
rect 23532 37068 23538 37080
rect 29638 37068 29644 37080
rect 29696 37068 29702 37120
rect 32858 37068 32864 37120
rect 32916 37108 32922 37120
rect 40862 37108 40868 37120
rect 32916 37080 40868 37108
rect 32916 37068 32922 37080
rect 40862 37068 40868 37080
rect 40920 37068 40926 37120
rect 40957 37111 41015 37117
rect 40957 37077 40969 37111
rect 41003 37108 41015 37111
rect 48314 37108 48320 37120
rect 41003 37080 48320 37108
rect 41003 37077 41015 37080
rect 40957 37071 41015 37077
rect 48314 37068 48320 37080
rect 48372 37068 48378 37120
rect 48498 37068 48504 37120
rect 48556 37108 48562 37120
rect 50706 37108 50712 37120
rect 48556 37080 50712 37108
rect 48556 37068 48562 37080
rect 50706 37068 50712 37080
rect 50764 37108 50770 37120
rect 65058 37108 65064 37120
rect 50764 37080 65064 37108
rect 50764 37068 50770 37080
rect 65058 37068 65064 37080
rect 65116 37068 65122 37120
rect 65150 37068 65156 37120
rect 65208 37108 65214 37120
rect 70026 37108 70032 37120
rect 65208 37080 70032 37108
rect 65208 37068 65214 37080
rect 70026 37068 70032 37080
rect 70084 37068 70090 37120
rect 71498 37068 71504 37120
rect 71556 37108 71562 37120
rect 71593 37111 71651 37117
rect 71593 37108 71605 37111
rect 71556 37080 71605 37108
rect 71556 37068 71562 37080
rect 71593 37077 71605 37080
rect 71639 37077 71651 37111
rect 89548 37108 89576 37148
rect 89686 37148 92121 37176
rect 89686 37108 89714 37148
rect 92109 37145 92121 37148
rect 92155 37145 92167 37179
rect 92109 37139 92167 37145
rect 89548 37080 89714 37108
rect 71593 37071 71651 37077
rect 1104 37018 98808 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 65686 37018
rect 65738 36966 65750 37018
rect 65802 36966 65814 37018
rect 65866 36966 65878 37018
rect 65930 36966 96406 37018
rect 96458 36966 96470 37018
rect 96522 36966 96534 37018
rect 96586 36966 96598 37018
rect 96650 36966 98808 37018
rect 1104 36944 98808 36966
rect 2590 36864 2596 36916
rect 2648 36904 2654 36916
rect 42058 36904 42064 36916
rect 2648 36876 42064 36904
rect 2648 36864 2654 36876
rect 42058 36864 42064 36876
rect 42116 36864 42122 36916
rect 42242 36864 42248 36916
rect 42300 36904 42306 36916
rect 46753 36907 46811 36913
rect 46753 36904 46765 36907
rect 42300 36876 46765 36904
rect 42300 36864 42306 36876
rect 46753 36873 46765 36876
rect 46799 36873 46811 36907
rect 46753 36867 46811 36873
rect 46934 36864 46940 36916
rect 46992 36904 46998 36916
rect 47029 36907 47087 36913
rect 47029 36904 47041 36907
rect 46992 36876 47041 36904
rect 46992 36864 46998 36876
rect 47029 36873 47041 36876
rect 47075 36873 47087 36907
rect 53558 36904 53564 36916
rect 47029 36867 47087 36873
rect 47136 36876 53564 36904
rect 2130 36836 2136 36848
rect 2091 36808 2136 36836
rect 2130 36796 2136 36808
rect 2188 36796 2194 36848
rect 7374 36796 7380 36848
rect 7432 36836 7438 36848
rect 7653 36839 7711 36845
rect 7653 36836 7665 36839
rect 7432 36808 7665 36836
rect 7432 36796 7438 36808
rect 7653 36805 7665 36808
rect 7699 36805 7711 36839
rect 7653 36799 7711 36805
rect 9950 36796 9956 36848
rect 10008 36836 10014 36848
rect 10229 36839 10287 36845
rect 10229 36836 10241 36839
rect 10008 36808 10241 36836
rect 10008 36796 10014 36808
rect 10229 36805 10241 36808
rect 10275 36805 10287 36839
rect 10229 36799 10287 36805
rect 12618 36796 12624 36848
rect 12676 36836 12682 36848
rect 12897 36839 12955 36845
rect 12897 36836 12909 36839
rect 12676 36808 12909 36836
rect 12676 36796 12682 36808
rect 12897 36805 12909 36808
rect 12943 36805 12955 36839
rect 12897 36799 12955 36805
rect 15286 36796 15292 36848
rect 15344 36836 15350 36848
rect 15565 36839 15623 36845
rect 15565 36836 15577 36839
rect 15344 36808 15577 36836
rect 15344 36796 15350 36808
rect 15565 36805 15577 36808
rect 15611 36805 15623 36839
rect 17862 36836 17868 36848
rect 17823 36808 17868 36836
rect 15565 36799 15623 36805
rect 17862 36796 17868 36808
rect 17920 36796 17926 36848
rect 19334 36796 19340 36848
rect 19392 36836 19398 36848
rect 19429 36839 19487 36845
rect 19429 36836 19441 36839
rect 19392 36808 19441 36836
rect 19392 36796 19398 36808
rect 19429 36805 19441 36808
rect 19475 36805 19487 36839
rect 19429 36799 19487 36805
rect 19518 36796 19524 36848
rect 19576 36836 19582 36848
rect 20346 36836 20352 36848
rect 19576 36808 20352 36836
rect 19576 36796 19582 36808
rect 20346 36796 20352 36808
rect 20404 36796 20410 36848
rect 20714 36796 20720 36848
rect 20772 36836 20778 36848
rect 20809 36839 20867 36845
rect 20809 36836 20821 36839
rect 20772 36808 20821 36836
rect 20772 36796 20778 36808
rect 20809 36805 20821 36808
rect 20855 36805 20867 36839
rect 20809 36799 20867 36805
rect 24486 36796 24492 36848
rect 24544 36836 24550 36848
rect 24544 36808 33640 36836
rect 24544 36796 24550 36808
rect 3234 36768 3240 36780
rect 3195 36740 3240 36768
rect 3234 36728 3240 36740
rect 3292 36728 3298 36780
rect 4617 36771 4675 36777
rect 4617 36737 4629 36771
rect 4663 36768 4675 36771
rect 23474 36768 23480 36780
rect 4663 36740 23480 36768
rect 4663 36737 4675 36740
rect 4617 36731 4675 36737
rect 23474 36728 23480 36740
rect 23532 36728 23538 36780
rect 33612 36768 33640 36808
rect 33686 36796 33692 36848
rect 33744 36836 33750 36848
rect 33965 36839 34023 36845
rect 33965 36836 33977 36839
rect 33744 36808 33977 36836
rect 33744 36796 33750 36808
rect 33965 36805 33977 36808
rect 34011 36805 34023 36839
rect 33965 36799 34023 36805
rect 36262 36796 36268 36848
rect 36320 36836 36326 36848
rect 36541 36839 36599 36845
rect 36541 36836 36553 36839
rect 36320 36808 36553 36836
rect 36320 36796 36326 36808
rect 36541 36805 36553 36808
rect 36587 36805 36599 36839
rect 36541 36799 36599 36805
rect 36630 36796 36636 36848
rect 36688 36836 36694 36848
rect 36688 36808 43484 36836
rect 36688 36796 36694 36808
rect 43456 36768 43484 36808
rect 47136 36768 47164 36876
rect 53558 36864 53564 36876
rect 53616 36864 53622 36916
rect 54496 36876 54708 36904
rect 54496 36836 54524 36876
rect 23584 36740 33548 36768
rect 33612 36740 43392 36768
rect 43456 36740 47164 36768
rect 47228 36808 54524 36836
rect 54680 36836 54708 36876
rect 54754 36864 54760 36916
rect 54812 36904 54818 36916
rect 54941 36907 54999 36913
rect 54941 36904 54953 36907
rect 54812 36876 54953 36904
rect 54812 36864 54818 36876
rect 54941 36873 54953 36876
rect 54987 36873 54999 36907
rect 54941 36867 54999 36873
rect 55214 36864 55220 36916
rect 55272 36904 55278 36916
rect 55309 36907 55367 36913
rect 55309 36904 55321 36907
rect 55272 36876 55321 36904
rect 55272 36864 55278 36876
rect 55309 36873 55321 36876
rect 55355 36904 55367 36907
rect 55493 36907 55551 36913
rect 55493 36904 55505 36907
rect 55355 36876 55505 36904
rect 55355 36873 55367 36876
rect 55309 36867 55367 36873
rect 55493 36873 55505 36876
rect 55539 36873 55551 36907
rect 55493 36867 55551 36873
rect 57330 36864 57336 36916
rect 57388 36904 57394 36916
rect 57517 36907 57575 36913
rect 57517 36904 57529 36907
rect 57388 36876 57529 36904
rect 57388 36864 57394 36876
rect 57517 36873 57529 36876
rect 57563 36873 57575 36907
rect 57517 36867 57575 36873
rect 59998 36864 60004 36916
rect 60056 36904 60062 36916
rect 60185 36907 60243 36913
rect 60185 36904 60197 36907
rect 60056 36876 60197 36904
rect 60056 36864 60062 36876
rect 60185 36873 60197 36876
rect 60231 36873 60243 36907
rect 60185 36867 60243 36873
rect 62574 36864 62580 36916
rect 62632 36904 62638 36916
rect 62761 36907 62819 36913
rect 62761 36904 62773 36907
rect 62632 36876 62773 36904
rect 62632 36864 62638 36876
rect 62761 36873 62773 36876
rect 62807 36873 62819 36907
rect 62761 36867 62819 36873
rect 65058 36864 65064 36916
rect 65116 36904 65122 36916
rect 70486 36904 70492 36916
rect 65116 36876 70492 36904
rect 65116 36864 65122 36876
rect 70486 36864 70492 36876
rect 70544 36864 70550 36916
rect 70578 36864 70584 36916
rect 70636 36904 70642 36916
rect 70673 36907 70731 36913
rect 70673 36904 70685 36907
rect 70636 36876 70685 36904
rect 70636 36864 70642 36876
rect 70673 36873 70685 36876
rect 70719 36873 70731 36907
rect 70673 36867 70731 36873
rect 72973 36907 73031 36913
rect 72973 36873 72985 36907
rect 73019 36904 73031 36907
rect 73154 36904 73160 36916
rect 73019 36876 73160 36904
rect 73019 36873 73031 36876
rect 72973 36867 73031 36873
rect 73154 36864 73160 36876
rect 73212 36864 73218 36916
rect 73246 36864 73252 36916
rect 73304 36904 73310 36916
rect 86954 36904 86960 36916
rect 73304 36876 86960 36904
rect 73304 36864 73310 36876
rect 86954 36864 86960 36876
rect 87012 36864 87018 36916
rect 88978 36836 88984 36848
rect 54680 36808 88984 36836
rect 2041 36703 2099 36709
rect 2041 36669 2053 36703
rect 2087 36700 2099 36703
rect 2314 36700 2320 36712
rect 2087 36672 2320 36700
rect 2087 36669 2099 36672
rect 2041 36663 2099 36669
rect 2314 36660 2320 36672
rect 2372 36660 2378 36712
rect 2961 36703 3019 36709
rect 2961 36669 2973 36703
rect 3007 36700 3019 36703
rect 3510 36700 3516 36712
rect 3007 36672 3516 36700
rect 3007 36669 3019 36672
rect 2961 36663 3019 36669
rect 3510 36660 3516 36672
rect 3568 36660 3574 36712
rect 8202 36700 8208 36712
rect 8163 36672 8208 36700
rect 8202 36660 8208 36672
rect 8260 36660 8266 36712
rect 15381 36703 15439 36709
rect 15381 36669 15393 36703
rect 15427 36700 15439 36703
rect 15470 36700 15476 36712
rect 15427 36672 15476 36700
rect 15427 36669 15439 36672
rect 15381 36663 15439 36669
rect 15470 36660 15476 36672
rect 15528 36660 15534 36712
rect 18693 36703 18751 36709
rect 18693 36669 18705 36703
rect 18739 36700 18751 36703
rect 19245 36703 19303 36709
rect 19245 36700 19257 36703
rect 18739 36672 19257 36700
rect 18739 36669 18751 36672
rect 18693 36663 18751 36669
rect 19245 36669 19257 36672
rect 19291 36700 19303 36703
rect 19291 36672 19472 36700
rect 19291 36669 19303 36672
rect 19245 36663 19303 36669
rect 7466 36632 7472 36644
rect 7427 36604 7472 36632
rect 7466 36592 7472 36604
rect 7524 36592 7530 36644
rect 10045 36635 10103 36641
rect 10045 36601 10057 36635
rect 10091 36632 10103 36635
rect 10318 36632 10324 36644
rect 10091 36604 10324 36632
rect 10091 36601 10103 36604
rect 10045 36595 10103 36601
rect 10318 36592 10324 36604
rect 10376 36592 10382 36644
rect 12713 36635 12771 36641
rect 12713 36601 12725 36635
rect 12759 36632 12771 36635
rect 17402 36632 17408 36644
rect 12759 36604 17408 36632
rect 12759 36601 12771 36604
rect 12713 36595 12771 36601
rect 17402 36592 17408 36604
rect 17460 36592 17466 36644
rect 17773 36635 17831 36641
rect 17773 36601 17785 36635
rect 17819 36632 17831 36635
rect 18049 36635 18107 36641
rect 18049 36632 18061 36635
rect 17819 36604 18061 36632
rect 17819 36601 17831 36604
rect 17773 36595 17831 36601
rect 18049 36601 18061 36604
rect 18095 36632 18107 36635
rect 19444 36632 19472 36672
rect 19518 36660 19524 36712
rect 19576 36700 19582 36712
rect 23584 36700 23612 36740
rect 26694 36700 26700 36712
rect 19576 36672 19621 36700
rect 19720 36672 23612 36700
rect 26655 36672 26700 36700
rect 19576 36660 19582 36672
rect 19720 36632 19748 36672
rect 26694 36660 26700 36672
rect 26752 36660 26758 36712
rect 28626 36700 28632 36712
rect 28587 36672 28632 36700
rect 28626 36660 28632 36672
rect 28684 36660 28690 36712
rect 29270 36660 29276 36712
rect 29328 36700 29334 36712
rect 29917 36703 29975 36709
rect 29917 36700 29929 36703
rect 29328 36672 29929 36700
rect 29328 36660 29334 36672
rect 29917 36669 29929 36672
rect 29963 36669 29975 36703
rect 29917 36663 29975 36669
rect 31389 36703 31447 36709
rect 31389 36669 31401 36703
rect 31435 36700 31447 36703
rect 31662 36700 31668 36712
rect 31435 36672 31668 36700
rect 31435 36669 31447 36672
rect 31389 36663 31447 36669
rect 31662 36660 31668 36672
rect 31720 36660 31726 36712
rect 33520 36700 33548 36740
rect 36630 36700 36636 36712
rect 33520 36672 36636 36700
rect 36630 36660 36636 36672
rect 36688 36660 36694 36712
rect 36722 36660 36728 36712
rect 36780 36700 36786 36712
rect 39942 36700 39948 36712
rect 36780 36672 39948 36700
rect 36780 36660 36786 36672
rect 39942 36660 39948 36672
rect 40000 36660 40006 36712
rect 42426 36700 42432 36712
rect 42387 36672 42432 36700
rect 42426 36660 42432 36672
rect 42484 36660 42490 36712
rect 18095 36604 19288 36632
rect 19444 36604 19748 36632
rect 18095 36601 18107 36604
rect 18049 36595 18107 36601
rect 8386 36564 8392 36576
rect 8347 36536 8392 36564
rect 8386 36524 8392 36536
rect 8444 36524 8450 36576
rect 19058 36564 19064 36576
rect 19019 36536 19064 36564
rect 19058 36524 19064 36536
rect 19116 36524 19122 36576
rect 19260 36564 19288 36604
rect 20254 36592 20260 36644
rect 20312 36632 20318 36644
rect 20625 36635 20683 36641
rect 20625 36632 20637 36635
rect 20312 36604 20637 36632
rect 20312 36592 20318 36604
rect 20625 36601 20637 36604
rect 20671 36601 20683 36635
rect 28258 36632 28264 36644
rect 20625 36595 20683 36601
rect 22066 36604 28264 36632
rect 22066 36564 22094 36604
rect 28258 36592 28264 36604
rect 28316 36592 28322 36644
rect 28994 36632 29000 36644
rect 28955 36604 29000 36632
rect 28994 36592 29000 36604
rect 29052 36592 29058 36644
rect 33781 36635 33839 36641
rect 29656 36604 31754 36632
rect 19260 36536 22094 36564
rect 26694 36524 26700 36576
rect 26752 36564 26758 36576
rect 26881 36567 26939 36573
rect 26881 36564 26893 36567
rect 26752 36536 26893 36564
rect 26752 36524 26758 36536
rect 26881 36533 26893 36536
rect 26927 36533 26939 36567
rect 26881 36527 26939 36533
rect 27430 36524 27436 36576
rect 27488 36564 27494 36576
rect 29656 36564 29684 36604
rect 27488 36536 29684 36564
rect 29733 36567 29791 36573
rect 27488 36524 27494 36536
rect 29733 36533 29745 36567
rect 29779 36564 29791 36567
rect 30282 36564 30288 36576
rect 29779 36536 30288 36564
rect 29779 36533 29791 36536
rect 29733 36527 29791 36533
rect 30282 36524 30288 36536
rect 30340 36524 30346 36576
rect 31726 36564 31754 36604
rect 33781 36601 33793 36635
rect 33827 36632 33839 36635
rect 33962 36632 33968 36644
rect 33827 36604 33968 36632
rect 33827 36601 33839 36604
rect 33781 36595 33839 36601
rect 33962 36592 33968 36604
rect 34020 36592 34026 36644
rect 36262 36592 36268 36644
rect 36320 36632 36326 36644
rect 36357 36635 36415 36641
rect 36357 36632 36369 36635
rect 36320 36604 36369 36632
rect 36320 36592 36326 36604
rect 36357 36601 36369 36604
rect 36403 36601 36415 36635
rect 42242 36632 42248 36644
rect 36357 36595 36415 36601
rect 36556 36604 42248 36632
rect 36556 36564 36584 36604
rect 42242 36592 42248 36604
rect 42300 36592 42306 36644
rect 31726 36536 36584 36564
rect 38102 36524 38108 36576
rect 38160 36564 38166 36576
rect 42613 36567 42671 36573
rect 42613 36564 42625 36567
rect 38160 36536 42625 36564
rect 38160 36524 38166 36536
rect 42613 36533 42625 36536
rect 42659 36533 42671 36567
rect 43364 36564 43392 36740
rect 43530 36700 43536 36712
rect 43491 36672 43536 36700
rect 43530 36660 43536 36672
rect 43588 36660 43594 36712
rect 43806 36700 43812 36712
rect 43767 36672 43812 36700
rect 43806 36660 43812 36672
rect 43864 36660 43870 36712
rect 47228 36700 47256 36808
rect 88978 36796 88984 36808
rect 89036 36796 89042 36848
rect 94222 36836 94228 36848
rect 94183 36808 94228 36836
rect 94222 36796 94228 36808
rect 94280 36796 94286 36848
rect 96798 36836 96804 36848
rect 96759 36808 96804 36836
rect 96798 36796 96804 36808
rect 96856 36796 96862 36848
rect 98089 36839 98147 36845
rect 98089 36805 98101 36839
rect 98135 36836 98147 36839
rect 99466 36836 99472 36848
rect 98135 36808 99472 36836
rect 98135 36805 98147 36808
rect 98089 36799 98147 36805
rect 99466 36796 99472 36808
rect 99524 36796 99530 36848
rect 47302 36728 47308 36780
rect 47360 36768 47366 36780
rect 53466 36768 53472 36780
rect 47360 36740 53472 36768
rect 47360 36728 47366 36740
rect 53466 36728 53472 36740
rect 53524 36728 53530 36780
rect 53558 36728 53564 36780
rect 53616 36768 53622 36780
rect 65150 36768 65156 36780
rect 53616 36740 65156 36768
rect 53616 36728 53622 36740
rect 65150 36728 65156 36740
rect 65208 36728 65214 36780
rect 67726 36768 67732 36780
rect 65260 36740 67732 36768
rect 44468 36672 47256 36700
rect 44468 36564 44496 36672
rect 47394 36660 47400 36712
rect 47452 36700 47458 36712
rect 47452 36672 55444 36700
rect 47452 36660 47458 36672
rect 46937 36635 46995 36641
rect 46937 36601 46949 36635
rect 46983 36632 46995 36635
rect 48222 36632 48228 36644
rect 46983 36604 48228 36632
rect 46983 36601 46995 36604
rect 46937 36595 46995 36601
rect 48222 36592 48228 36604
rect 48280 36592 48286 36644
rect 48314 36592 48320 36644
rect 48372 36632 48378 36644
rect 52914 36632 52920 36644
rect 48372 36604 52920 36632
rect 48372 36592 48378 36604
rect 52914 36592 52920 36604
rect 52972 36592 52978 36644
rect 54570 36592 54576 36644
rect 54628 36632 54634 36644
rect 54849 36635 54907 36641
rect 54849 36632 54861 36635
rect 54628 36604 54861 36632
rect 54628 36592 54634 36604
rect 54849 36601 54861 36604
rect 54895 36601 54907 36635
rect 55416 36632 55444 36672
rect 55582 36660 55588 36712
rect 55640 36700 55646 36712
rect 56137 36703 56195 36709
rect 56137 36700 56149 36703
rect 55640 36672 56149 36700
rect 55640 36660 55646 36672
rect 56137 36669 56149 36672
rect 56183 36669 56195 36703
rect 65260 36700 65288 36740
rect 67726 36728 67732 36740
rect 67784 36728 67790 36780
rect 68186 36728 68192 36780
rect 68244 36768 68250 36780
rect 93854 36768 93860 36780
rect 68244 36740 93860 36768
rect 68244 36728 68250 36740
rect 93854 36728 93860 36740
rect 93912 36728 93918 36780
rect 65426 36700 65432 36712
rect 56137 36663 56195 36669
rect 56244 36672 65288 36700
rect 65387 36672 65432 36700
rect 56244 36632 56272 36672
rect 65426 36660 65432 36672
rect 65484 36700 65490 36712
rect 67818 36700 67824 36712
rect 65484 36672 67824 36700
rect 65484 36660 65490 36672
rect 67818 36660 67824 36672
rect 67876 36660 67882 36712
rect 68462 36660 68468 36712
rect 68520 36700 68526 36712
rect 68649 36703 68707 36709
rect 68649 36700 68661 36703
rect 68520 36672 68661 36700
rect 68520 36660 68526 36672
rect 68649 36669 68661 36672
rect 68695 36669 68707 36703
rect 70578 36700 70584 36712
rect 70539 36672 70584 36700
rect 68649 36663 68707 36669
rect 70578 36660 70584 36672
rect 70636 36660 70642 36712
rect 73709 36703 73767 36709
rect 73709 36700 73721 36703
rect 71976 36672 73721 36700
rect 57422 36632 57428 36644
rect 54849 36595 54907 36601
rect 54956 36604 55352 36632
rect 55416 36604 56272 36632
rect 57383 36604 57428 36632
rect 45094 36564 45100 36576
rect 43364 36536 44496 36564
rect 45007 36536 45100 36564
rect 42613 36527 42671 36533
rect 45094 36524 45100 36536
rect 45152 36564 45158 36576
rect 46658 36564 46664 36576
rect 45152 36536 46664 36564
rect 45152 36524 45158 36536
rect 46658 36524 46664 36536
rect 46716 36524 46722 36576
rect 46753 36567 46811 36573
rect 46753 36533 46765 36567
rect 46799 36564 46811 36567
rect 52086 36564 52092 36576
rect 46799 36536 52092 36564
rect 46799 36533 46811 36536
rect 46753 36527 46811 36533
rect 52086 36524 52092 36536
rect 52144 36524 52150 36576
rect 52178 36524 52184 36576
rect 52236 36564 52242 36576
rect 54956 36564 54984 36604
rect 52236 36536 54984 36564
rect 55324 36564 55352 36604
rect 57422 36592 57428 36604
rect 57480 36592 57486 36644
rect 60090 36632 60096 36644
rect 60051 36604 60096 36632
rect 60090 36592 60096 36604
rect 60148 36592 60154 36644
rect 62666 36632 62672 36644
rect 62627 36604 62672 36632
rect 62666 36592 62672 36604
rect 62724 36592 62730 36644
rect 65610 36632 65616 36644
rect 62960 36604 65616 36632
rect 55766 36564 55772 36576
rect 55324 36536 55772 36564
rect 52236 36524 52242 36536
rect 55766 36524 55772 36536
rect 55824 36524 55830 36576
rect 56318 36564 56324 36576
rect 56279 36536 56324 36564
rect 56318 36524 56324 36536
rect 56376 36524 56382 36576
rect 56502 36524 56508 36576
rect 56560 36564 56566 36576
rect 62960 36564 62988 36604
rect 65610 36592 65616 36604
rect 65668 36592 65674 36644
rect 65794 36632 65800 36644
rect 65755 36604 65800 36632
rect 65794 36592 65800 36604
rect 65852 36592 65858 36644
rect 68002 36632 68008 36644
rect 67963 36604 68008 36632
rect 68002 36592 68008 36604
rect 68060 36592 68066 36644
rect 68189 36635 68247 36641
rect 68189 36601 68201 36635
rect 68235 36632 68247 36635
rect 68278 36632 68284 36644
rect 68235 36604 68284 36632
rect 68235 36601 68247 36604
rect 68189 36595 68247 36601
rect 68278 36592 68284 36604
rect 68336 36592 68342 36644
rect 56560 36536 62988 36564
rect 56560 36524 56566 36536
rect 63034 36524 63040 36576
rect 63092 36564 63098 36576
rect 65518 36564 65524 36576
rect 63092 36536 65524 36564
rect 63092 36524 63098 36536
rect 65518 36524 65524 36536
rect 65576 36524 65582 36576
rect 68462 36564 68468 36576
rect 68423 36536 68468 36564
rect 68462 36524 68468 36536
rect 68520 36524 68526 36576
rect 68554 36524 68560 36576
rect 68612 36564 68618 36576
rect 71976 36564 72004 36672
rect 73709 36669 73721 36672
rect 73755 36669 73767 36703
rect 73982 36700 73988 36712
rect 73943 36672 73988 36700
rect 73709 36663 73767 36669
rect 73982 36660 73988 36672
rect 74040 36660 74046 36712
rect 75822 36660 75828 36712
rect 75880 36700 75886 36712
rect 76101 36703 76159 36709
rect 76101 36700 76113 36703
rect 75880 36672 76113 36700
rect 75880 36660 75886 36672
rect 76101 36669 76113 36672
rect 76147 36669 76159 36703
rect 76101 36663 76159 36669
rect 76190 36660 76196 36712
rect 76248 36700 76254 36712
rect 78493 36703 78551 36709
rect 78493 36700 78505 36703
rect 76248 36672 78505 36700
rect 76248 36660 76254 36672
rect 78493 36669 78505 36672
rect 78539 36669 78551 36703
rect 78674 36700 78680 36712
rect 78635 36672 78680 36700
rect 78493 36663 78551 36669
rect 78674 36660 78680 36672
rect 78732 36660 78738 36712
rect 79137 36703 79195 36709
rect 79137 36669 79149 36703
rect 79183 36700 79195 36703
rect 79318 36700 79324 36712
rect 79183 36672 79324 36700
rect 79183 36669 79195 36672
rect 79137 36663 79195 36669
rect 79318 36660 79324 36672
rect 79376 36660 79382 36712
rect 84381 36703 84439 36709
rect 84381 36669 84393 36703
rect 84427 36700 84439 36703
rect 84562 36700 84568 36712
rect 84427 36672 84568 36700
rect 84427 36669 84439 36672
rect 84381 36663 84439 36669
rect 84562 36660 84568 36672
rect 84620 36660 84626 36712
rect 87138 36700 87144 36712
rect 87099 36672 87144 36700
rect 87138 36660 87144 36672
rect 87196 36660 87202 36712
rect 89625 36703 89683 36709
rect 89625 36669 89637 36703
rect 89671 36700 89683 36703
rect 89806 36700 89812 36712
rect 89671 36672 89812 36700
rect 89671 36669 89683 36672
rect 89625 36663 89683 36669
rect 89806 36660 89812 36672
rect 89864 36660 89870 36712
rect 92474 36700 92480 36712
rect 92435 36672 92480 36700
rect 92474 36660 92480 36672
rect 92532 36660 92538 36712
rect 72878 36632 72884 36644
rect 72839 36604 72884 36632
rect 72878 36592 72884 36604
rect 72936 36592 72942 36644
rect 75914 36632 75920 36644
rect 72988 36604 74028 36632
rect 75875 36604 75920 36632
rect 68612 36536 72004 36564
rect 68612 36524 68618 36536
rect 72050 36524 72056 36576
rect 72108 36564 72114 36576
rect 72988 36564 73016 36604
rect 72108 36536 73016 36564
rect 72108 36524 72114 36536
rect 73430 36524 73436 36576
rect 73488 36564 73494 36576
rect 73525 36567 73583 36573
rect 73525 36564 73537 36567
rect 73488 36536 73537 36564
rect 73488 36524 73494 36536
rect 73525 36533 73537 36536
rect 73571 36533 73583 36567
rect 73525 36527 73583 36533
rect 73798 36524 73804 36576
rect 73856 36564 73862 36576
rect 73893 36567 73951 36573
rect 73893 36564 73905 36567
rect 73856 36536 73905 36564
rect 73856 36524 73862 36536
rect 73893 36533 73905 36536
rect 73939 36533 73951 36567
rect 74000 36564 74028 36604
rect 75914 36592 75920 36604
rect 75972 36592 75978 36644
rect 94133 36635 94191 36641
rect 94133 36632 94145 36635
rect 76024 36604 94145 36632
rect 76024 36564 76052 36604
rect 94133 36601 94145 36604
rect 94179 36632 94191 36635
rect 94409 36635 94467 36641
rect 94409 36632 94421 36635
rect 94179 36604 94421 36632
rect 94179 36601 94191 36604
rect 94133 36595 94191 36601
rect 94409 36601 94421 36604
rect 94455 36601 94467 36635
rect 94409 36595 94467 36601
rect 96985 36635 97043 36641
rect 96985 36601 96997 36635
rect 97031 36601 97043 36635
rect 97626 36632 97632 36644
rect 97587 36604 97632 36632
rect 96985 36595 97043 36601
rect 74000 36536 76052 36564
rect 79321 36567 79379 36573
rect 73893 36527 73951 36533
rect 79321 36533 79333 36567
rect 79367 36564 79379 36567
rect 79410 36564 79416 36576
rect 79367 36536 79416 36564
rect 79367 36533 79379 36536
rect 79321 36527 79379 36533
rect 79410 36524 79416 36536
rect 79468 36524 79474 36576
rect 96614 36564 96620 36576
rect 96575 36536 96620 36564
rect 96614 36524 96620 36536
rect 96672 36564 96678 36576
rect 97000 36564 97028 36595
rect 97626 36592 97632 36604
rect 97684 36632 97690 36644
rect 97905 36635 97963 36641
rect 97905 36632 97917 36635
rect 97684 36604 97917 36632
rect 97684 36592 97690 36604
rect 97905 36601 97917 36604
rect 97951 36632 97963 36635
rect 98181 36635 98239 36641
rect 98181 36632 98193 36635
rect 97951 36604 98193 36632
rect 97951 36601 97963 36604
rect 97905 36595 97963 36601
rect 98181 36601 98193 36604
rect 98227 36601 98239 36635
rect 98181 36595 98239 36601
rect 96672 36536 97028 36564
rect 96672 36524 96678 36536
rect 1104 36474 98808 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 50326 36474
rect 50378 36422 50390 36474
rect 50442 36422 50454 36474
rect 50506 36422 50518 36474
rect 50570 36422 81046 36474
rect 81098 36422 81110 36474
rect 81162 36422 81174 36474
rect 81226 36422 81238 36474
rect 81290 36422 98808 36474
rect 1104 36400 98808 36422
rect 8294 36360 8300 36372
rect 5644 36332 8300 36360
rect 4890 36184 4896 36236
rect 4948 36224 4954 36236
rect 5644 36233 5672 36332
rect 8294 36320 8300 36332
rect 8352 36320 8358 36372
rect 8386 36320 8392 36372
rect 8444 36360 8450 36372
rect 24762 36360 24768 36372
rect 8444 36332 24768 36360
rect 8444 36320 8450 36332
rect 24762 36320 24768 36332
rect 24820 36320 24826 36372
rect 24946 36320 24952 36372
rect 25004 36360 25010 36372
rect 26786 36360 26792 36372
rect 25004 36332 26792 36360
rect 25004 36320 25010 36332
rect 26786 36320 26792 36332
rect 26844 36320 26850 36372
rect 50893 36363 50951 36369
rect 50893 36360 50905 36363
rect 28184 36332 50905 36360
rect 12805 36295 12863 36301
rect 12805 36292 12817 36295
rect 5736 36264 12817 36292
rect 5736 36233 5764 36264
rect 12805 36261 12817 36264
rect 12851 36261 12863 36295
rect 28184 36292 28212 36332
rect 50893 36329 50905 36332
rect 50939 36329 50951 36363
rect 50893 36323 50951 36329
rect 51000 36332 55720 36360
rect 12805 36255 12863 36261
rect 12912 36264 28212 36292
rect 5261 36227 5319 36233
rect 5261 36224 5273 36227
rect 4948 36196 5273 36224
rect 4948 36184 4954 36196
rect 5261 36193 5273 36196
rect 5307 36193 5319 36227
rect 5261 36187 5319 36193
rect 5629 36227 5687 36233
rect 5629 36193 5641 36227
rect 5675 36193 5687 36227
rect 5629 36187 5687 36193
rect 5721 36227 5779 36233
rect 5721 36193 5733 36227
rect 5767 36193 5779 36227
rect 5721 36187 5779 36193
rect 5997 36227 6055 36233
rect 5997 36193 6009 36227
rect 6043 36224 6055 36227
rect 6178 36224 6184 36236
rect 6043 36196 6184 36224
rect 6043 36193 6055 36196
rect 5997 36187 6055 36193
rect 6178 36184 6184 36196
rect 6236 36184 6242 36236
rect 6089 36159 6147 36165
rect 6089 36125 6101 36159
rect 6135 36125 6147 36159
rect 6089 36119 6147 36125
rect 6104 36088 6132 36119
rect 10962 36116 10968 36168
rect 11020 36156 11026 36168
rect 12912 36156 12940 36264
rect 12986 36184 12992 36236
rect 13044 36224 13050 36236
rect 18417 36227 18475 36233
rect 13044 36196 13089 36224
rect 13044 36184 13050 36196
rect 18417 36193 18429 36227
rect 18463 36224 18475 36227
rect 18690 36224 18696 36236
rect 18463 36196 18696 36224
rect 18463 36193 18475 36196
rect 18417 36187 18475 36193
rect 18690 36184 18696 36196
rect 18748 36184 18754 36236
rect 27430 36224 27436 36236
rect 27391 36196 27436 36224
rect 27430 36184 27436 36196
rect 27488 36184 27494 36236
rect 27798 36224 27804 36236
rect 27759 36196 27804 36224
rect 27798 36184 27804 36196
rect 27856 36184 27862 36236
rect 28184 36233 28212 36264
rect 28258 36252 28264 36304
rect 28316 36292 28322 36304
rect 33410 36292 33416 36304
rect 28316 36264 33416 36292
rect 28316 36252 28322 36264
rect 33410 36252 33416 36264
rect 33468 36252 33474 36304
rect 34146 36252 34152 36304
rect 34204 36292 34210 36304
rect 42150 36292 42156 36304
rect 34204 36264 42156 36292
rect 34204 36252 34210 36264
rect 42150 36252 42156 36264
rect 42208 36252 42214 36304
rect 42242 36252 42248 36304
rect 42300 36292 42306 36304
rect 46934 36292 46940 36304
rect 42300 36264 46940 36292
rect 42300 36252 42306 36264
rect 46934 36252 46940 36264
rect 46992 36252 46998 36304
rect 51000 36292 51028 36332
rect 48286 36264 51028 36292
rect 52104 36264 55444 36292
rect 28169 36227 28227 36233
rect 28169 36193 28181 36227
rect 28215 36193 28227 36227
rect 28169 36187 28227 36193
rect 33686 36184 33692 36236
rect 33744 36224 33750 36236
rect 36722 36224 36728 36236
rect 33744 36196 36728 36224
rect 33744 36184 33750 36196
rect 36722 36184 36728 36196
rect 36780 36184 36786 36236
rect 37458 36184 37464 36236
rect 37516 36224 37522 36236
rect 43346 36224 43352 36236
rect 37516 36196 43352 36224
rect 37516 36184 37522 36196
rect 43346 36184 43352 36196
rect 43404 36184 43410 36236
rect 43530 36184 43536 36236
rect 43588 36224 43594 36236
rect 47213 36227 47271 36233
rect 47213 36224 47225 36227
rect 43588 36196 47225 36224
rect 43588 36184 43594 36196
rect 47213 36193 47225 36196
rect 47259 36193 47271 36227
rect 47213 36187 47271 36193
rect 47762 36184 47768 36236
rect 47820 36224 47826 36236
rect 48286 36224 48314 36264
rect 47820 36196 48314 36224
rect 47820 36184 47826 36196
rect 48682 36184 48688 36236
rect 48740 36224 48746 36236
rect 49602 36224 49608 36236
rect 48740 36196 49608 36224
rect 48740 36184 48746 36196
rect 49602 36184 49608 36196
rect 49660 36224 49666 36236
rect 52104 36224 52132 36264
rect 49660 36196 52132 36224
rect 49660 36184 49666 36196
rect 52178 36184 52184 36236
rect 52236 36224 52242 36236
rect 52236 36196 52281 36224
rect 52236 36184 52242 36196
rect 52362 36184 52368 36236
rect 52420 36224 52426 36236
rect 54846 36224 54852 36236
rect 52420 36196 54852 36224
rect 52420 36184 52426 36196
rect 54846 36184 54852 36196
rect 54904 36184 54910 36236
rect 55032 36227 55090 36233
rect 55032 36193 55044 36227
rect 55078 36193 55090 36227
rect 55032 36187 55090 36193
rect 55217 36227 55275 36233
rect 55217 36193 55229 36227
rect 55263 36224 55275 36227
rect 55306 36224 55312 36236
rect 55263 36196 55312 36224
rect 55263 36193 55275 36196
rect 55217 36187 55275 36193
rect 11020 36128 12940 36156
rect 13541 36159 13599 36165
rect 11020 36116 11026 36128
rect 13541 36125 13553 36159
rect 13587 36156 13599 36159
rect 14090 36156 14096 36168
rect 13587 36128 14096 36156
rect 13587 36125 13599 36128
rect 13541 36119 13599 36125
rect 14090 36116 14096 36128
rect 14148 36116 14154 36168
rect 22094 36116 22100 36168
rect 22152 36156 22158 36168
rect 22152 36128 22876 36156
rect 22152 36116 22158 36128
rect 22848 36088 22876 36128
rect 24302 36116 24308 36168
rect 24360 36156 24366 36168
rect 27617 36159 27675 36165
rect 27617 36156 27629 36159
rect 24360 36128 27629 36156
rect 24360 36116 24366 36128
rect 27617 36125 27629 36128
rect 27663 36125 27675 36159
rect 28074 36156 28080 36168
rect 28035 36128 28080 36156
rect 27617 36119 27675 36125
rect 28074 36116 28080 36128
rect 28132 36116 28138 36168
rect 28718 36156 28724 36168
rect 28679 36128 28724 36156
rect 28718 36116 28724 36128
rect 28776 36116 28782 36168
rect 31662 36116 31668 36168
rect 31720 36156 31726 36168
rect 41414 36156 41420 36168
rect 31720 36128 41420 36156
rect 31720 36116 31726 36128
rect 41414 36116 41420 36128
rect 41472 36116 41478 36168
rect 41506 36116 41512 36168
rect 41564 36156 41570 36168
rect 46934 36156 46940 36168
rect 41564 36128 46940 36156
rect 41564 36116 41570 36128
rect 46934 36116 46940 36128
rect 46992 36116 46998 36168
rect 47394 36116 47400 36168
rect 47452 36156 47458 36168
rect 47489 36159 47547 36165
rect 47489 36156 47501 36159
rect 47452 36128 47501 36156
rect 47452 36116 47458 36128
rect 47489 36125 47501 36128
rect 47535 36125 47547 36159
rect 47489 36119 47547 36125
rect 47578 36116 47584 36168
rect 47636 36156 47642 36168
rect 51166 36156 51172 36168
rect 47636 36128 51172 36156
rect 47636 36116 47642 36128
rect 51166 36116 51172 36128
rect 51224 36156 51230 36168
rect 52270 36156 52276 36168
rect 51224 36128 52276 36156
rect 51224 36116 51230 36128
rect 52270 36116 52276 36128
rect 52328 36116 52334 36168
rect 52730 36156 52736 36168
rect 52691 36128 52736 36156
rect 52730 36116 52736 36128
rect 52788 36116 52794 36168
rect 53006 36116 53012 36168
rect 53064 36156 53070 36168
rect 55048 36156 55076 36187
rect 55306 36184 55312 36196
rect 55364 36184 55370 36236
rect 55416 36233 55444 36264
rect 55490 36252 55496 36304
rect 55548 36292 55554 36304
rect 55585 36295 55643 36301
rect 55585 36292 55597 36295
rect 55548 36264 55597 36292
rect 55548 36252 55554 36264
rect 55585 36261 55597 36264
rect 55631 36261 55643 36295
rect 55585 36255 55643 36261
rect 55401 36227 55459 36233
rect 55401 36193 55413 36227
rect 55447 36193 55459 36227
rect 55692 36224 55720 36332
rect 55766 36320 55772 36372
rect 55824 36360 55830 36372
rect 65426 36360 65432 36372
rect 55824 36332 65432 36360
rect 55824 36320 55830 36332
rect 65426 36320 65432 36332
rect 65484 36320 65490 36372
rect 65518 36320 65524 36372
rect 65576 36360 65582 36372
rect 70486 36360 70492 36372
rect 65576 36332 70492 36360
rect 65576 36320 65582 36332
rect 70486 36320 70492 36332
rect 70544 36320 70550 36372
rect 70578 36320 70584 36372
rect 70636 36360 70642 36372
rect 70636 36332 75316 36360
rect 70636 36320 70642 36332
rect 55858 36252 55864 36304
rect 55916 36292 55922 36304
rect 59814 36292 59820 36304
rect 55916 36264 59820 36292
rect 55916 36252 55922 36264
rect 59814 36252 59820 36264
rect 59872 36252 59878 36304
rect 72878 36292 72884 36304
rect 64064 36264 72884 36292
rect 55401 36187 55459 36193
rect 55600 36196 55720 36224
rect 55600 36168 55628 36196
rect 56594 36184 56600 36236
rect 56652 36224 56658 36236
rect 64064 36224 64092 36264
rect 72878 36252 72884 36264
rect 72936 36252 72942 36304
rect 73816 36264 74028 36292
rect 65334 36224 65340 36236
rect 56652 36196 64092 36224
rect 65295 36196 65340 36224
rect 56652 36184 56658 36196
rect 65334 36184 65340 36196
rect 65392 36184 65398 36236
rect 70210 36224 70216 36236
rect 65444 36196 70216 36224
rect 53064 36128 55076 36156
rect 53064 36116 53070 36128
rect 55122 36116 55128 36168
rect 55180 36156 55186 36168
rect 55180 36128 55225 36156
rect 55180 36116 55186 36128
rect 55582 36116 55588 36168
rect 55640 36116 55646 36168
rect 55950 36116 55956 36168
rect 56008 36156 56014 36168
rect 59354 36156 59360 36168
rect 56008 36128 59360 36156
rect 56008 36116 56014 36128
rect 59354 36116 59360 36128
rect 59412 36116 59418 36168
rect 63126 36156 63132 36168
rect 63087 36128 63132 36156
rect 63126 36116 63132 36128
rect 63184 36116 63190 36168
rect 63402 36156 63408 36168
rect 63363 36128 63408 36156
rect 63402 36116 63408 36128
rect 63460 36116 63466 36168
rect 64966 36116 64972 36168
rect 65024 36156 65030 36168
rect 65444 36156 65472 36196
rect 70210 36184 70216 36196
rect 70268 36184 70274 36236
rect 70302 36184 70308 36236
rect 70360 36224 70366 36236
rect 73816 36224 73844 36264
rect 70360 36196 73844 36224
rect 73893 36227 73951 36233
rect 70360 36184 70366 36196
rect 73893 36193 73905 36227
rect 73939 36193 73951 36227
rect 73893 36187 73951 36193
rect 65024 36128 65472 36156
rect 65024 36116 65030 36128
rect 65610 36116 65616 36168
rect 65668 36156 65674 36168
rect 73908 36156 73936 36187
rect 65668 36128 73936 36156
rect 74000 36156 74028 36264
rect 75288 36224 75316 36332
rect 76006 36320 76012 36372
rect 76064 36360 76070 36372
rect 96614 36360 96620 36372
rect 76064 36332 96620 36360
rect 76064 36320 76070 36332
rect 96614 36320 96620 36332
rect 96672 36320 96678 36372
rect 81618 36224 81624 36236
rect 75288 36196 81624 36224
rect 81618 36184 81624 36196
rect 81676 36184 81682 36236
rect 93489 36227 93547 36233
rect 93489 36193 93501 36227
rect 93535 36224 93547 36227
rect 93854 36224 93860 36236
rect 93535 36196 93860 36224
rect 93535 36193 93547 36196
rect 93489 36187 93547 36193
rect 93854 36184 93860 36196
rect 93912 36224 93918 36236
rect 94590 36224 94596 36236
rect 93912 36196 94596 36224
rect 93912 36184 93918 36196
rect 94590 36184 94596 36196
rect 94648 36184 94654 36236
rect 95050 36224 95056 36236
rect 95011 36196 95056 36224
rect 95050 36184 95056 36196
rect 95108 36184 95114 36236
rect 97537 36227 97595 36233
rect 97537 36193 97549 36227
rect 97583 36224 97595 36227
rect 97718 36224 97724 36236
rect 97583 36196 97724 36224
rect 97583 36193 97595 36196
rect 97537 36187 97595 36193
rect 97718 36184 97724 36196
rect 97776 36184 97782 36236
rect 74261 36159 74319 36165
rect 74261 36156 74273 36159
rect 74000 36128 74273 36156
rect 65668 36116 65674 36128
rect 74261 36125 74273 36128
rect 74307 36125 74319 36159
rect 94038 36156 94044 36168
rect 93999 36128 94044 36156
rect 74261 36119 74319 36125
rect 94038 36116 94044 36128
rect 94096 36116 94102 36168
rect 35250 36088 35256 36100
rect 6104 36060 22094 36088
rect 22848 36060 35256 36088
rect 6454 36020 6460 36032
rect 6415 35992 6460 36020
rect 6454 35980 6460 35992
rect 6512 35980 6518 36032
rect 12805 36023 12863 36029
rect 12805 35989 12817 36023
rect 12851 36020 12863 36023
rect 13906 36020 13912 36032
rect 12851 35992 13912 36020
rect 12851 35989 12863 35992
rect 12805 35983 12863 35989
rect 13906 35980 13912 35992
rect 13964 35980 13970 36032
rect 22066 36020 22094 36060
rect 35250 36048 35256 36060
rect 35308 36048 35314 36100
rect 37185 36091 37243 36097
rect 37185 36057 37197 36091
rect 37231 36088 37243 36091
rect 37461 36091 37519 36097
rect 37461 36088 37473 36091
rect 37231 36060 37473 36088
rect 37231 36057 37243 36060
rect 37185 36051 37243 36057
rect 37461 36057 37473 36060
rect 37507 36088 37519 36091
rect 47118 36088 47124 36100
rect 37507 36060 43576 36088
rect 47079 36060 47124 36088
rect 37507 36057 37519 36060
rect 37461 36051 37519 36057
rect 33318 36020 33324 36032
rect 22066 35992 33324 36020
rect 33318 35980 33324 35992
rect 33376 35980 33382 36032
rect 33410 35980 33416 36032
rect 33468 36020 33474 36032
rect 43438 36020 43444 36032
rect 33468 35992 43444 36020
rect 33468 35980 33474 35992
rect 43438 35980 43444 35992
rect 43496 35980 43502 36032
rect 43548 36020 43576 36060
rect 47118 36048 47124 36060
rect 47176 36048 47182 36100
rect 48406 36048 48412 36100
rect 48464 36088 48470 36100
rect 48777 36091 48835 36097
rect 48777 36088 48789 36091
rect 48464 36060 48789 36088
rect 48464 36048 48470 36060
rect 48777 36057 48789 36060
rect 48823 36057 48835 36091
rect 48777 36051 48835 36057
rect 55858 36048 55864 36100
rect 55916 36088 55922 36100
rect 63034 36088 63040 36100
rect 55916 36060 63040 36088
rect 55916 36048 55922 36060
rect 63034 36048 63040 36060
rect 63092 36048 63098 36100
rect 65150 36048 65156 36100
rect 65208 36088 65214 36100
rect 65521 36091 65579 36097
rect 65521 36088 65533 36091
rect 65208 36060 65533 36088
rect 65208 36048 65214 36060
rect 65521 36057 65533 36060
rect 65567 36057 65579 36091
rect 75914 36088 75920 36100
rect 65521 36051 65579 36057
rect 66088 36060 75920 36088
rect 48590 36020 48596 36032
rect 43548 35992 48596 36020
rect 48590 35980 48596 35992
rect 48648 35980 48654 36032
rect 50893 36023 50951 36029
rect 50893 35989 50905 36023
rect 50939 36020 50951 36023
rect 55306 36020 55312 36032
rect 50939 35992 55312 36020
rect 50939 35989 50951 35992
rect 50893 35983 50951 35989
rect 55306 35980 55312 35992
rect 55364 35980 55370 36032
rect 55582 35980 55588 36032
rect 55640 36020 55646 36032
rect 64509 36023 64567 36029
rect 64509 36020 64521 36023
rect 55640 35992 64521 36020
rect 55640 35980 55646 35992
rect 64509 35989 64521 35992
rect 64555 35989 64567 36023
rect 64509 35983 64567 35989
rect 64598 35980 64604 36032
rect 64656 36020 64662 36032
rect 66088 36020 66116 36060
rect 75914 36048 75920 36060
rect 75972 36048 75978 36100
rect 64656 35992 66116 36020
rect 64656 35980 64662 35992
rect 66162 35980 66168 36032
rect 66220 36020 66226 36032
rect 73522 36020 73528 36032
rect 66220 35992 73528 36020
rect 66220 35980 66226 35992
rect 73522 35980 73528 35992
rect 73580 35980 73586 36032
rect 73614 35980 73620 36032
rect 73672 36020 73678 36032
rect 74031 36023 74089 36029
rect 74031 36020 74043 36023
rect 73672 35992 74043 36020
rect 73672 35980 73678 35992
rect 74031 35989 74043 35992
rect 74077 35989 74089 36023
rect 74166 36020 74172 36032
rect 74127 35992 74172 36020
rect 74031 35983 74089 35989
rect 74166 35980 74172 35992
rect 74224 35980 74230 36032
rect 74534 36020 74540 36032
rect 74495 35992 74540 36020
rect 74534 35980 74540 35992
rect 74592 35980 74598 36032
rect 1104 35930 98808 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 65686 35930
rect 65738 35878 65750 35930
rect 65802 35878 65814 35930
rect 65866 35878 65878 35930
rect 65930 35878 96406 35930
rect 96458 35878 96470 35930
rect 96522 35878 96534 35930
rect 96586 35878 96598 35930
rect 96650 35878 98808 35930
rect 1104 35856 98808 35878
rect 24486 35816 24492 35828
rect 24447 35788 24492 35816
rect 24486 35776 24492 35788
rect 24544 35776 24550 35828
rect 28626 35776 28632 35828
rect 28684 35816 28690 35828
rect 33502 35816 33508 35828
rect 28684 35788 33508 35816
rect 28684 35776 28690 35788
rect 33502 35776 33508 35788
rect 33560 35776 33566 35828
rect 43530 35816 43536 35828
rect 33796 35788 43536 35816
rect 20162 35708 20168 35760
rect 20220 35748 20226 35760
rect 33796 35748 33824 35788
rect 43530 35776 43536 35788
rect 43588 35776 43594 35828
rect 44174 35776 44180 35828
rect 44232 35816 44238 35828
rect 48130 35816 48136 35828
rect 44232 35788 48136 35816
rect 44232 35776 44238 35788
rect 48130 35776 48136 35788
rect 48188 35776 48194 35828
rect 48222 35776 48228 35828
rect 48280 35816 48286 35828
rect 51074 35816 51080 35828
rect 48280 35788 51080 35816
rect 48280 35776 48286 35788
rect 51074 35776 51080 35788
rect 51132 35776 51138 35828
rect 51166 35776 51172 35828
rect 51224 35816 51230 35828
rect 57057 35819 57115 35825
rect 57057 35816 57069 35819
rect 51224 35788 57069 35816
rect 51224 35776 51230 35788
rect 57057 35785 57069 35788
rect 57103 35785 57115 35819
rect 57057 35779 57115 35785
rect 57146 35776 57152 35828
rect 57204 35816 57210 35828
rect 79134 35816 79140 35828
rect 57204 35788 79140 35816
rect 57204 35776 57210 35788
rect 79134 35776 79140 35788
rect 79192 35776 79198 35828
rect 91554 35776 91560 35828
rect 91612 35816 91618 35828
rect 95234 35816 95240 35828
rect 91612 35788 95240 35816
rect 91612 35776 91618 35788
rect 95234 35776 95240 35788
rect 95292 35776 95298 35828
rect 20220 35720 33824 35748
rect 20220 35708 20226 35720
rect 33870 35708 33876 35760
rect 33928 35748 33934 35760
rect 39022 35748 39028 35760
rect 33928 35720 39028 35748
rect 33928 35708 33934 35720
rect 39022 35708 39028 35720
rect 39080 35708 39086 35760
rect 46750 35708 46756 35760
rect 46808 35748 46814 35760
rect 55582 35748 55588 35760
rect 46808 35720 55588 35748
rect 46808 35708 46814 35720
rect 55582 35708 55588 35720
rect 55640 35708 55646 35760
rect 66990 35748 66996 35760
rect 56612 35720 66996 35748
rect 11882 35640 11888 35692
rect 11940 35680 11946 35692
rect 39482 35680 39488 35692
rect 11940 35652 39488 35680
rect 11940 35640 11946 35652
rect 39482 35640 39488 35652
rect 39540 35640 39546 35692
rect 39574 35640 39580 35692
rect 39632 35680 39638 35692
rect 40034 35680 40040 35692
rect 39632 35652 40040 35680
rect 39632 35640 39638 35652
rect 40034 35640 40040 35652
rect 40092 35680 40098 35692
rect 43622 35680 43628 35692
rect 40092 35652 43628 35680
rect 40092 35640 40098 35652
rect 43622 35640 43628 35652
rect 43680 35640 43686 35692
rect 45094 35680 45100 35692
rect 43732 35652 45100 35680
rect 18877 35615 18935 35621
rect 18877 35581 18889 35615
rect 18923 35612 18935 35615
rect 19150 35612 19156 35624
rect 18923 35584 19156 35612
rect 18923 35581 18935 35584
rect 18877 35575 18935 35581
rect 19150 35572 19156 35584
rect 19208 35572 19214 35624
rect 24670 35612 24676 35624
rect 24631 35584 24676 35612
rect 24670 35572 24676 35584
rect 24728 35572 24734 35624
rect 24762 35572 24768 35624
rect 24820 35612 24826 35624
rect 24857 35615 24915 35621
rect 24857 35612 24869 35615
rect 24820 35584 24869 35612
rect 24820 35572 24826 35584
rect 24857 35581 24869 35584
rect 24903 35581 24915 35615
rect 25222 35612 25228 35624
rect 25183 35584 25228 35612
rect 24857 35575 24915 35581
rect 25222 35572 25228 35584
rect 25280 35572 25286 35624
rect 25409 35615 25467 35621
rect 25409 35581 25421 35615
rect 25455 35612 25467 35615
rect 39298 35612 39304 35624
rect 25455 35584 39304 35612
rect 25455 35581 25467 35584
rect 25409 35575 25467 35581
rect 39298 35572 39304 35584
rect 39356 35572 39362 35624
rect 39390 35572 39396 35624
rect 39448 35612 39454 35624
rect 39847 35615 39905 35621
rect 39847 35612 39859 35615
rect 39448 35584 39859 35612
rect 39448 35572 39454 35584
rect 39847 35581 39859 35584
rect 39893 35581 39905 35615
rect 39847 35575 39905 35581
rect 41138 35572 41144 35624
rect 41196 35612 41202 35624
rect 43732 35612 43760 35652
rect 45094 35640 45100 35652
rect 45152 35640 45158 35692
rect 46566 35640 46572 35692
rect 46624 35680 46630 35692
rect 47486 35680 47492 35692
rect 46624 35652 47492 35680
rect 46624 35640 46630 35652
rect 47486 35640 47492 35652
rect 47544 35640 47550 35692
rect 48314 35640 48320 35692
rect 48372 35680 48378 35692
rect 49878 35680 49884 35692
rect 48372 35652 49884 35680
rect 48372 35640 48378 35652
rect 49878 35640 49884 35652
rect 49936 35640 49942 35692
rect 56612 35680 56640 35720
rect 66990 35708 66996 35720
rect 67048 35708 67054 35760
rect 67726 35708 67732 35760
rect 67784 35748 67790 35760
rect 72694 35748 72700 35760
rect 67784 35720 72700 35748
rect 67784 35708 67790 35720
rect 72694 35708 72700 35720
rect 72752 35708 72758 35760
rect 88334 35748 88340 35760
rect 80026 35720 88340 35748
rect 49988 35652 56640 35680
rect 41196 35584 43760 35612
rect 41196 35572 41202 35584
rect 43806 35572 43812 35624
rect 43864 35612 43870 35624
rect 46106 35612 46112 35624
rect 43864 35584 46112 35612
rect 43864 35572 43870 35584
rect 46106 35572 46112 35584
rect 46164 35572 46170 35624
rect 46658 35572 46664 35624
rect 46716 35612 46722 35624
rect 49988 35612 50016 35652
rect 56686 35640 56692 35692
rect 56744 35680 56750 35692
rect 80026 35680 80054 35720
rect 88334 35708 88340 35720
rect 88392 35708 88398 35760
rect 56744 35652 80054 35680
rect 82265 35683 82323 35689
rect 56744 35640 56750 35652
rect 82265 35649 82277 35683
rect 82311 35680 82323 35683
rect 82354 35680 82360 35692
rect 82311 35652 82360 35680
rect 82311 35649 82323 35652
rect 82265 35643 82323 35649
rect 82354 35640 82360 35652
rect 82412 35640 82418 35692
rect 46716 35584 50016 35612
rect 46716 35572 46722 35584
rect 51074 35572 51080 35624
rect 51132 35612 51138 35624
rect 55490 35612 55496 35624
rect 51132 35584 55496 35612
rect 51132 35572 51138 35584
rect 55490 35572 55496 35584
rect 55548 35572 55554 35624
rect 55677 35615 55735 35621
rect 55677 35581 55689 35615
rect 55723 35612 55735 35615
rect 55766 35612 55772 35624
rect 55723 35584 55772 35612
rect 55723 35581 55735 35584
rect 55677 35575 55735 35581
rect 55766 35572 55772 35584
rect 55824 35572 55830 35624
rect 55950 35612 55956 35624
rect 55911 35584 55956 35612
rect 55950 35572 55956 35584
rect 56008 35572 56014 35624
rect 56042 35572 56048 35624
rect 56100 35612 56106 35624
rect 57146 35612 57152 35624
rect 56100 35584 57152 35612
rect 56100 35572 56106 35584
rect 57146 35572 57152 35584
rect 57204 35572 57210 35624
rect 61838 35572 61844 35624
rect 61896 35612 61902 35624
rect 66714 35612 66720 35624
rect 61896 35584 66720 35612
rect 61896 35572 61902 35584
rect 66714 35572 66720 35584
rect 66772 35572 66778 35624
rect 66990 35572 66996 35624
rect 67048 35612 67054 35624
rect 81894 35612 81900 35624
rect 67048 35584 80054 35612
rect 81855 35584 81900 35612
rect 67048 35572 67054 35584
rect 12986 35504 12992 35556
rect 13044 35544 13050 35556
rect 35986 35544 35992 35556
rect 13044 35516 35992 35544
rect 13044 35504 13050 35516
rect 35986 35504 35992 35516
rect 36044 35504 36050 35556
rect 36354 35504 36360 35556
rect 36412 35544 36418 35556
rect 39666 35544 39672 35556
rect 36412 35516 39672 35544
rect 36412 35504 36418 35516
rect 39666 35504 39672 35516
rect 39724 35504 39730 35556
rect 41046 35504 41052 35556
rect 41104 35544 41110 35556
rect 55306 35544 55312 35556
rect 41104 35516 55312 35544
rect 41104 35504 41110 35516
rect 55306 35504 55312 35516
rect 55364 35504 55370 35556
rect 56612 35516 60734 35544
rect 28994 35436 29000 35488
rect 29052 35476 29058 35488
rect 36446 35476 36452 35488
rect 29052 35448 36452 35476
rect 29052 35436 29058 35448
rect 36446 35436 36452 35448
rect 36504 35436 36510 35488
rect 36538 35436 36544 35488
rect 36596 35476 36602 35488
rect 39390 35476 39396 35488
rect 36596 35448 39396 35476
rect 36596 35436 36602 35448
rect 39390 35436 39396 35448
rect 39448 35436 39454 35488
rect 40954 35476 40960 35488
rect 40915 35448 40960 35476
rect 40954 35436 40960 35448
rect 41012 35436 41018 35488
rect 41322 35436 41328 35488
rect 41380 35476 41386 35488
rect 43898 35476 43904 35488
rect 41380 35448 43904 35476
rect 41380 35436 41386 35448
rect 43898 35436 43904 35448
rect 43956 35436 43962 35488
rect 46382 35436 46388 35488
rect 46440 35476 46446 35488
rect 56612 35476 56640 35516
rect 46440 35448 56640 35476
rect 60706 35476 60734 35516
rect 65150 35504 65156 35556
rect 65208 35544 65214 35556
rect 76006 35544 76012 35556
rect 65208 35516 76012 35544
rect 65208 35504 65214 35516
rect 76006 35504 76012 35516
rect 76064 35504 76070 35556
rect 80026 35544 80054 35584
rect 81894 35572 81900 35584
rect 81952 35572 81958 35624
rect 81986 35572 81992 35624
rect 82044 35621 82050 35624
rect 82044 35615 82103 35621
rect 82044 35581 82057 35615
rect 82091 35581 82103 35615
rect 82044 35575 82103 35581
rect 82044 35572 82050 35575
rect 82170 35572 82176 35624
rect 82228 35612 82234 35624
rect 82449 35615 82507 35621
rect 82228 35584 82273 35612
rect 82228 35572 82234 35584
rect 82449 35581 82461 35615
rect 82495 35581 82507 35615
rect 82449 35575 82507 35581
rect 82464 35544 82492 35575
rect 80026 35516 82492 35544
rect 82541 35479 82599 35485
rect 82541 35476 82553 35479
rect 60706 35448 82553 35476
rect 46440 35436 46446 35448
rect 82541 35445 82553 35448
rect 82587 35445 82599 35479
rect 82541 35439 82599 35445
rect 1104 35386 98808 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 50326 35386
rect 50378 35334 50390 35386
rect 50442 35334 50454 35386
rect 50506 35334 50518 35386
rect 50570 35334 81046 35386
rect 81098 35334 81110 35386
rect 81162 35334 81174 35386
rect 81226 35334 81238 35386
rect 81290 35334 98808 35386
rect 1104 35312 98808 35334
rect 19150 35232 19156 35284
rect 19208 35272 19214 35284
rect 46566 35272 46572 35284
rect 19208 35244 46572 35272
rect 19208 35232 19214 35244
rect 46566 35232 46572 35244
rect 46624 35232 46630 35284
rect 56318 35272 56324 35284
rect 46952 35244 56324 35272
rect 12158 35164 12164 35216
rect 12216 35204 12222 35216
rect 24302 35204 24308 35216
rect 12216 35176 24308 35204
rect 12216 35164 12222 35176
rect 24302 35164 24308 35176
rect 24360 35164 24366 35216
rect 36354 35204 36360 35216
rect 31726 35176 36360 35204
rect 17405 35139 17463 35145
rect 17405 35105 17417 35139
rect 17451 35136 17463 35139
rect 19978 35136 19984 35148
rect 17451 35108 19984 35136
rect 17451 35105 17463 35108
rect 17405 35099 17463 35105
rect 19978 35096 19984 35108
rect 20036 35096 20042 35148
rect 23658 35096 23664 35148
rect 23716 35136 23722 35148
rect 31726 35136 31754 35176
rect 36354 35164 36360 35176
rect 36412 35164 36418 35216
rect 36446 35164 36452 35216
rect 36504 35204 36510 35216
rect 43346 35204 43352 35216
rect 36504 35176 43352 35204
rect 36504 35164 36510 35176
rect 43346 35164 43352 35176
rect 43404 35164 43410 35216
rect 43530 35204 43536 35216
rect 43491 35176 43536 35204
rect 43530 35164 43536 35176
rect 43588 35164 43594 35216
rect 43993 35207 44051 35213
rect 43993 35173 44005 35207
rect 44039 35204 44051 35207
rect 44266 35204 44272 35216
rect 44039 35176 44272 35204
rect 44039 35173 44051 35176
rect 43993 35167 44051 35173
rect 44266 35164 44272 35176
rect 44324 35164 44330 35216
rect 46952 35213 46980 35244
rect 56318 35232 56324 35244
rect 56376 35232 56382 35284
rect 59354 35232 59360 35284
rect 59412 35272 59418 35284
rect 96706 35272 96712 35284
rect 59412 35244 96712 35272
rect 59412 35232 59418 35244
rect 96706 35232 96712 35244
rect 96764 35232 96770 35284
rect 46937 35207 46995 35213
rect 46937 35173 46949 35207
rect 46983 35173 46995 35207
rect 46937 35167 46995 35173
rect 47029 35207 47087 35213
rect 47029 35173 47041 35207
rect 47075 35204 47087 35207
rect 52178 35204 52184 35216
rect 47075 35176 52184 35204
rect 47075 35173 47087 35176
rect 47029 35167 47087 35173
rect 52178 35164 52184 35176
rect 52236 35164 52242 35216
rect 52270 35164 52276 35216
rect 52328 35204 52334 35216
rect 56686 35204 56692 35216
rect 52328 35176 56692 35204
rect 52328 35164 52334 35176
rect 56686 35164 56692 35176
rect 56744 35164 56750 35216
rect 56778 35164 56784 35216
rect 56836 35204 56842 35216
rect 56836 35176 62068 35204
rect 56836 35164 56842 35176
rect 62040 35148 62068 35176
rect 65978 35164 65984 35216
rect 66036 35204 66042 35216
rect 85945 35207 86003 35213
rect 85945 35204 85957 35207
rect 66036 35176 85957 35204
rect 66036 35164 66042 35176
rect 85945 35173 85957 35176
rect 85991 35204 86003 35207
rect 85991 35176 86172 35204
rect 85991 35173 86003 35176
rect 85945 35167 86003 35173
rect 23716 35108 31754 35136
rect 36541 35139 36599 35145
rect 23716 35096 23722 35108
rect 36541 35105 36553 35139
rect 36587 35136 36599 35139
rect 36814 35136 36820 35148
rect 36587 35108 36820 35136
rect 36587 35105 36599 35108
rect 36541 35099 36599 35105
rect 36814 35096 36820 35108
rect 36872 35096 36878 35148
rect 36906 35096 36912 35148
rect 36964 35136 36970 35148
rect 41322 35136 41328 35148
rect 36964 35108 41328 35136
rect 36964 35096 36970 35108
rect 41322 35096 41328 35108
rect 41380 35096 41386 35148
rect 41414 35096 41420 35148
rect 41472 35136 41478 35148
rect 42978 35136 42984 35148
rect 41472 35108 42984 35136
rect 41472 35096 41478 35108
rect 42978 35096 42984 35108
rect 43036 35096 43042 35148
rect 43714 35096 43720 35148
rect 43772 35136 43778 35148
rect 43898 35136 43904 35148
rect 43772 35108 43817 35136
rect 43859 35108 43904 35136
rect 43772 35096 43778 35108
rect 43898 35096 43904 35108
rect 43956 35096 43962 35148
rect 46750 35136 46756 35148
rect 46711 35108 46756 35136
rect 46750 35096 46756 35108
rect 46808 35096 46814 35148
rect 47118 35096 47124 35148
rect 47176 35145 47182 35148
rect 47176 35136 47184 35145
rect 47176 35108 47221 35136
rect 47176 35099 47184 35108
rect 47176 35096 47182 35099
rect 47302 35096 47308 35148
rect 47360 35145 47366 35148
rect 47360 35139 47380 35145
rect 47368 35105 47380 35139
rect 47360 35099 47380 35105
rect 47360 35096 47366 35099
rect 47486 35096 47492 35148
rect 47544 35136 47550 35148
rect 52362 35136 52368 35148
rect 47544 35108 52368 35136
rect 47544 35096 47550 35108
rect 52362 35096 52368 35108
rect 52420 35096 52426 35148
rect 53926 35096 53932 35148
rect 53984 35136 53990 35148
rect 54113 35139 54171 35145
rect 54113 35136 54125 35139
rect 53984 35108 54125 35136
rect 53984 35096 53990 35108
rect 54113 35105 54125 35108
rect 54159 35105 54171 35139
rect 54113 35099 54171 35105
rect 55582 35096 55588 35148
rect 55640 35136 55646 35148
rect 61838 35136 61844 35148
rect 55640 35108 61844 35136
rect 55640 35096 55646 35108
rect 61838 35096 61844 35108
rect 61896 35096 61902 35148
rect 62022 35136 62028 35148
rect 61983 35108 62028 35136
rect 62022 35096 62028 35108
rect 62080 35096 62086 35148
rect 62132 35108 62436 35136
rect 14458 35028 14464 35080
rect 14516 35068 14522 35080
rect 62132 35068 62160 35108
rect 14516 35040 62160 35068
rect 14516 35028 14522 35040
rect 62206 35028 62212 35080
rect 62264 35068 62270 35080
rect 62301 35071 62359 35077
rect 62301 35068 62313 35071
rect 62264 35040 62313 35068
rect 62264 35028 62270 35040
rect 62301 35037 62313 35040
rect 62347 35037 62359 35071
rect 62408 35068 62436 35108
rect 62574 35096 62580 35148
rect 62632 35136 62638 35148
rect 64598 35136 64604 35148
rect 62632 35108 64604 35136
rect 62632 35096 62638 35108
rect 64598 35096 64604 35108
rect 64656 35096 64662 35148
rect 68094 35136 68100 35148
rect 68055 35108 68100 35136
rect 68094 35096 68100 35108
rect 68152 35096 68158 35148
rect 68186 35096 68192 35148
rect 68244 35136 68250 35148
rect 68465 35139 68523 35145
rect 68465 35136 68477 35139
rect 68244 35108 68477 35136
rect 68244 35096 68250 35108
rect 68465 35105 68477 35108
rect 68511 35105 68523 35139
rect 68830 35136 68836 35148
rect 68791 35108 68836 35136
rect 68465 35099 68523 35105
rect 68830 35096 68836 35108
rect 68888 35096 68894 35148
rect 70026 35096 70032 35148
rect 70084 35136 70090 35148
rect 72326 35136 72332 35148
rect 70084 35108 72332 35136
rect 70084 35096 70090 35108
rect 72326 35096 72332 35108
rect 72384 35096 72390 35148
rect 78858 35136 78864 35148
rect 78819 35108 78864 35136
rect 78858 35096 78864 35108
rect 78916 35096 78922 35148
rect 86144 35145 86172 35176
rect 86236 35176 86724 35204
rect 86129 35139 86187 35145
rect 86129 35105 86141 35139
rect 86175 35105 86187 35139
rect 86129 35099 86187 35105
rect 68281 35071 68339 35077
rect 68281 35068 68293 35071
rect 62408 35040 68293 35068
rect 62301 35031 62359 35037
rect 68281 35037 68293 35040
rect 68327 35037 68339 35071
rect 68738 35068 68744 35080
rect 68699 35040 68744 35068
rect 68281 35031 68339 35037
rect 68738 35028 68744 35040
rect 68796 35028 68802 35080
rect 68922 35028 68928 35080
rect 68980 35068 68986 35080
rect 79137 35071 79195 35077
rect 79137 35068 79149 35071
rect 68980 35040 79149 35068
rect 68980 35028 68986 35040
rect 79137 35037 79149 35040
rect 79183 35037 79195 35071
rect 79137 35031 79195 35037
rect 85853 35071 85911 35077
rect 85853 35037 85865 35071
rect 85899 35068 85911 35071
rect 86236 35068 86264 35176
rect 86310 35096 86316 35148
rect 86368 35136 86374 35148
rect 86696 35145 86724 35176
rect 86681 35139 86739 35145
rect 86368 35108 86412 35136
rect 86368 35096 86374 35108
rect 86681 35105 86693 35139
rect 86727 35105 86739 35139
rect 86681 35099 86739 35105
rect 94958 35096 94964 35148
rect 95016 35136 95022 35148
rect 95053 35139 95111 35145
rect 95053 35136 95065 35139
rect 95016 35108 95065 35136
rect 95016 35096 95022 35108
rect 95053 35105 95065 35108
rect 95099 35105 95111 35139
rect 95053 35099 95111 35105
rect 86402 35068 86408 35080
rect 85899 35040 86264 35068
rect 86363 35040 86408 35068
rect 85899 35037 85911 35040
rect 85853 35031 85911 35037
rect 86402 35028 86408 35040
rect 86460 35028 86466 35080
rect 86497 35071 86555 35077
rect 86497 35037 86509 35071
rect 86543 35068 86555 35071
rect 95418 35068 95424 35080
rect 86543 35040 86724 35068
rect 95379 35040 95424 35068
rect 86543 35037 86555 35040
rect 86497 35031 86555 35037
rect 86696 35012 86724 35040
rect 95418 35028 95424 35040
rect 95476 35028 95482 35080
rect 6730 34960 6736 35012
rect 6788 35000 6794 35012
rect 6788 34972 17540 35000
rect 6788 34960 6794 34972
rect 17512 34932 17540 34972
rect 21542 34960 21548 35012
rect 21600 35000 21606 35012
rect 54110 35000 54116 35012
rect 21600 34972 54116 35000
rect 21600 34960 21606 34972
rect 54110 34960 54116 34972
rect 54168 34960 54174 35012
rect 67729 35003 67787 35009
rect 67729 35000 67741 35003
rect 54220 34972 62068 35000
rect 54220 34932 54248 34972
rect 54386 34932 54392 34944
rect 17512 34904 54248 34932
rect 54347 34904 54392 34932
rect 54386 34892 54392 34904
rect 54444 34892 54450 34944
rect 57146 34892 57152 34944
rect 57204 34932 57210 34944
rect 59354 34932 59360 34944
rect 57204 34904 59360 34932
rect 57204 34892 57210 34904
rect 59354 34892 59360 34904
rect 59412 34892 59418 34944
rect 61838 34932 61844 34944
rect 61799 34904 61844 34932
rect 61838 34892 61844 34904
rect 61896 34892 61902 34944
rect 62040 34932 62068 34972
rect 63420 34972 67741 35000
rect 63420 34932 63448 34972
rect 67729 34969 67741 34972
rect 67775 35000 67787 35003
rect 67913 35003 67971 35009
rect 67913 35000 67925 35003
rect 67775 34972 67925 35000
rect 67775 34969 67787 34972
rect 67729 34963 67787 34969
rect 67913 34969 67925 34972
rect 67959 35000 67971 35003
rect 69201 35003 69259 35009
rect 69201 35000 69213 35003
rect 67959 34972 69213 35000
rect 67959 34969 67971 34972
rect 67913 34963 67971 34969
rect 69201 34969 69213 34972
rect 69247 35000 69259 35003
rect 69569 35003 69627 35009
rect 69569 35000 69581 35003
rect 69247 34972 69581 35000
rect 69247 34969 69259 34972
rect 69201 34963 69259 34969
rect 69569 34969 69581 34972
rect 69615 35000 69627 35003
rect 69753 35003 69811 35009
rect 69753 35000 69765 35003
rect 69615 34972 69765 35000
rect 69615 34969 69627 34972
rect 69569 34963 69627 34969
rect 69753 34969 69765 34972
rect 69799 34969 69811 35003
rect 69753 34963 69811 34969
rect 70366 34972 86080 35000
rect 62040 34904 63448 34932
rect 63494 34892 63500 34944
rect 63552 34932 63558 34944
rect 63589 34935 63647 34941
rect 63589 34932 63601 34935
rect 63552 34904 63601 34932
rect 63552 34892 63558 34904
rect 63589 34901 63601 34904
rect 63635 34901 63647 34935
rect 63589 34895 63647 34901
rect 64230 34892 64236 34944
rect 64288 34932 64294 34944
rect 70366 34932 70394 34972
rect 64288 34904 70394 34932
rect 64288 34892 64294 34904
rect 76282 34892 76288 34944
rect 76340 34932 76346 34944
rect 77202 34932 77208 34944
rect 76340 34904 77208 34932
rect 76340 34892 76346 34904
rect 77202 34892 77208 34904
rect 77260 34932 77266 34944
rect 85853 34935 85911 34941
rect 85853 34932 85865 34935
rect 77260 34904 85865 34932
rect 77260 34892 77266 34904
rect 85853 34901 85865 34904
rect 85899 34901 85911 34935
rect 86052 34932 86080 34972
rect 86678 34960 86684 35012
rect 86736 34960 86742 35012
rect 86773 34935 86831 34941
rect 86773 34932 86785 34935
rect 86052 34904 86785 34932
rect 85853 34895 85911 34901
rect 86773 34901 86785 34904
rect 86819 34901 86831 34935
rect 86773 34895 86831 34901
rect 86862 34892 86868 34944
rect 86920 34932 86926 34944
rect 95191 34935 95249 34941
rect 95191 34932 95203 34935
rect 86920 34904 95203 34932
rect 86920 34892 86926 34904
rect 95191 34901 95203 34904
rect 95237 34901 95249 34935
rect 95326 34932 95332 34944
rect 95287 34904 95332 34932
rect 95191 34895 95249 34901
rect 95326 34892 95332 34904
rect 95384 34892 95390 34944
rect 95510 34932 95516 34944
rect 95471 34904 95516 34932
rect 95510 34892 95516 34904
rect 95568 34892 95574 34944
rect 1104 34842 98808 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 65686 34842
rect 65738 34790 65750 34842
rect 65802 34790 65814 34842
rect 65866 34790 65878 34842
rect 65930 34790 96406 34842
rect 96458 34790 96470 34842
rect 96522 34790 96534 34842
rect 96586 34790 96598 34842
rect 96650 34790 98808 34842
rect 1104 34768 98808 34790
rect 27709 34731 27767 34737
rect 27709 34697 27721 34731
rect 27755 34728 27767 34731
rect 27982 34728 27988 34740
rect 27755 34700 27988 34728
rect 27755 34697 27767 34700
rect 27709 34691 27767 34697
rect 27982 34688 27988 34700
rect 28040 34688 28046 34740
rect 31662 34688 31668 34740
rect 31720 34728 31726 34740
rect 31720 34700 36584 34728
rect 31720 34688 31726 34700
rect 7558 34620 7564 34672
rect 7616 34660 7622 34672
rect 36446 34660 36452 34672
rect 7616 34632 36452 34660
rect 7616 34620 7622 34632
rect 36446 34620 36452 34632
rect 36504 34620 36510 34672
rect 16114 34552 16120 34604
rect 16172 34592 16178 34604
rect 36556 34592 36584 34700
rect 36814 34688 36820 34740
rect 36872 34728 36878 34740
rect 92106 34728 92112 34740
rect 36872 34700 92112 34728
rect 36872 34688 36878 34700
rect 92106 34688 92112 34700
rect 92164 34688 92170 34740
rect 40773 34663 40831 34669
rect 40773 34629 40785 34663
rect 40819 34660 40831 34663
rect 40862 34660 40868 34672
rect 40819 34632 40868 34660
rect 40819 34629 40831 34632
rect 40773 34623 40831 34629
rect 40862 34620 40868 34632
rect 40920 34620 40926 34672
rect 41506 34620 41512 34672
rect 41564 34660 41570 34672
rect 43530 34660 43536 34672
rect 41564 34632 43536 34660
rect 41564 34620 41570 34632
rect 43530 34620 43536 34632
rect 43588 34620 43594 34672
rect 43622 34620 43628 34672
rect 43680 34660 43686 34672
rect 49694 34660 49700 34672
rect 43680 34632 49700 34660
rect 43680 34620 43686 34632
rect 49694 34620 49700 34632
rect 49752 34620 49758 34672
rect 49786 34620 49792 34672
rect 49844 34660 49850 34672
rect 50798 34660 50804 34672
rect 49844 34632 50804 34660
rect 49844 34620 49850 34632
rect 50798 34620 50804 34632
rect 50856 34660 50862 34672
rect 50982 34660 50988 34672
rect 50856 34632 50988 34660
rect 50856 34620 50862 34632
rect 50982 34620 50988 34632
rect 51040 34620 51046 34672
rect 53098 34620 53104 34672
rect 53156 34660 53162 34672
rect 86862 34660 86868 34672
rect 53156 34632 86868 34660
rect 53156 34620 53162 34632
rect 86862 34620 86868 34632
rect 86920 34620 86926 34672
rect 83458 34592 83464 34604
rect 16172 34564 36492 34592
rect 36556 34564 39528 34592
rect 16172 34552 16178 34564
rect 19334 34484 19340 34536
rect 19392 34524 19398 34536
rect 24394 34524 24400 34536
rect 19392 34496 24400 34524
rect 19392 34484 19398 34496
rect 24394 34484 24400 34496
rect 24452 34484 24458 34536
rect 25314 34484 25320 34536
rect 25372 34524 25378 34536
rect 27798 34524 27804 34536
rect 25372 34496 27804 34524
rect 25372 34484 25378 34496
rect 27798 34484 27804 34496
rect 27856 34524 27862 34536
rect 27856 34496 29132 34524
rect 27856 34484 27862 34496
rect 18690 34416 18696 34468
rect 18748 34456 18754 34468
rect 28994 34456 29000 34468
rect 18748 34428 29000 34456
rect 18748 34416 18754 34428
rect 28994 34416 29000 34428
rect 29052 34416 29058 34468
rect 29104 34456 29132 34496
rect 29822 34484 29828 34536
rect 29880 34524 29886 34536
rect 34146 34524 34152 34536
rect 29880 34496 34152 34524
rect 29880 34484 29886 34496
rect 34146 34484 34152 34496
rect 34204 34484 34210 34536
rect 34514 34524 34520 34536
rect 34475 34496 34520 34524
rect 34514 34484 34520 34496
rect 34572 34524 34578 34536
rect 34793 34527 34851 34533
rect 34793 34524 34805 34527
rect 34572 34496 34805 34524
rect 34572 34484 34578 34496
rect 34793 34493 34805 34496
rect 34839 34493 34851 34527
rect 36464 34524 36492 34564
rect 39500 34536 39528 34564
rect 40420 34564 83464 34592
rect 36906 34524 36912 34536
rect 36464 34496 36912 34524
rect 34793 34487 34851 34493
rect 36906 34484 36912 34496
rect 36964 34484 36970 34536
rect 37274 34484 37280 34536
rect 37332 34524 37338 34536
rect 38194 34524 38200 34536
rect 37332 34496 38200 34524
rect 37332 34484 37338 34496
rect 38194 34484 38200 34496
rect 38252 34484 38258 34536
rect 39390 34524 39396 34536
rect 39351 34496 39396 34524
rect 39390 34484 39396 34496
rect 39448 34484 39454 34536
rect 39482 34484 39488 34536
rect 39540 34484 39546 34536
rect 39666 34533 39672 34536
rect 39649 34527 39672 34533
rect 39649 34493 39661 34527
rect 39649 34487 39672 34493
rect 39666 34484 39672 34487
rect 39724 34484 39730 34536
rect 39942 34484 39948 34536
rect 40000 34524 40006 34536
rect 40420 34524 40448 34564
rect 83458 34552 83464 34564
rect 83516 34552 83522 34604
rect 87046 34552 87052 34604
rect 87104 34592 87110 34604
rect 88886 34592 88892 34604
rect 87104 34564 88892 34592
rect 87104 34552 87110 34564
rect 88886 34552 88892 34564
rect 88944 34552 88950 34604
rect 40000 34496 40448 34524
rect 40000 34484 40006 34496
rect 40494 34484 40500 34536
rect 40552 34524 40558 34536
rect 41506 34524 41512 34536
rect 40552 34496 41512 34524
rect 40552 34484 40558 34496
rect 41506 34484 41512 34496
rect 41564 34484 41570 34536
rect 43530 34484 43536 34536
rect 43588 34524 43594 34536
rect 46842 34524 46848 34536
rect 43588 34496 46848 34524
rect 43588 34484 43594 34496
rect 46842 34484 46848 34496
rect 46900 34484 46906 34536
rect 46934 34484 46940 34536
rect 46992 34524 46998 34536
rect 53098 34524 53104 34536
rect 46992 34496 53104 34524
rect 46992 34484 46998 34496
rect 53098 34484 53104 34496
rect 53156 34484 53162 34536
rect 54202 34484 54208 34536
rect 54260 34524 54266 34536
rect 54260 34496 59308 34524
rect 54260 34484 54266 34496
rect 54846 34456 54852 34468
rect 29104 34428 54852 34456
rect 54846 34416 54852 34428
rect 54904 34456 54910 34468
rect 55122 34456 55128 34468
rect 54904 34428 55128 34456
rect 54904 34416 54910 34428
rect 55122 34416 55128 34428
rect 55180 34416 55186 34468
rect 55306 34416 55312 34468
rect 55364 34456 55370 34468
rect 58618 34456 58624 34468
rect 55364 34428 58624 34456
rect 55364 34416 55370 34428
rect 58618 34416 58624 34428
rect 58676 34416 58682 34468
rect 59280 34456 59308 34496
rect 59354 34484 59360 34536
rect 59412 34524 59418 34536
rect 59412 34496 59457 34524
rect 59412 34484 59418 34496
rect 59630 34484 59636 34536
rect 59688 34524 59694 34536
rect 59725 34527 59783 34533
rect 59725 34524 59737 34527
rect 59688 34496 59737 34524
rect 59688 34484 59694 34496
rect 59725 34493 59737 34496
rect 59771 34493 59783 34527
rect 64966 34524 64972 34536
rect 59725 34487 59783 34493
rect 59832 34496 64972 34524
rect 59832 34456 59860 34496
rect 64966 34484 64972 34496
rect 65024 34484 65030 34536
rect 65978 34484 65984 34536
rect 66036 34524 66042 34536
rect 67082 34524 67088 34536
rect 66036 34496 67088 34524
rect 66036 34484 66042 34496
rect 67082 34484 67088 34496
rect 67140 34484 67146 34536
rect 67177 34527 67235 34533
rect 67177 34493 67189 34527
rect 67223 34524 67235 34527
rect 67450 34524 67456 34536
rect 67223 34496 67456 34524
rect 67223 34493 67235 34496
rect 67177 34487 67235 34493
rect 67450 34484 67456 34496
rect 67508 34484 67514 34536
rect 67542 34484 67548 34536
rect 67600 34524 67606 34536
rect 68922 34524 68928 34536
rect 67600 34496 68928 34524
rect 67600 34484 67606 34496
rect 68922 34484 68928 34496
rect 68980 34484 68986 34536
rect 73709 34527 73767 34533
rect 73709 34493 73721 34527
rect 73755 34524 73767 34527
rect 73985 34527 74043 34533
rect 73985 34524 73997 34527
rect 73755 34496 73997 34524
rect 73755 34493 73767 34496
rect 73709 34487 73767 34493
rect 73985 34493 73997 34496
rect 74031 34524 74043 34527
rect 75178 34524 75184 34536
rect 74031 34496 75184 34524
rect 74031 34493 74043 34496
rect 73985 34487 74043 34493
rect 75178 34484 75184 34496
rect 75236 34484 75242 34536
rect 75546 34484 75552 34536
rect 75604 34524 75610 34536
rect 81713 34527 81771 34533
rect 81713 34524 81725 34527
rect 75604 34496 81725 34524
rect 75604 34484 75610 34496
rect 81713 34493 81725 34496
rect 81759 34493 81771 34527
rect 81713 34487 81771 34493
rect 82265 34527 82323 34533
rect 82265 34493 82277 34527
rect 82311 34524 82323 34527
rect 83274 34524 83280 34536
rect 82311 34496 83280 34524
rect 82311 34493 82323 34496
rect 82265 34487 82323 34493
rect 83274 34484 83280 34496
rect 83332 34484 83338 34536
rect 94222 34524 94228 34536
rect 94183 34496 94228 34524
rect 94222 34484 94228 34496
rect 94280 34524 94286 34536
rect 94593 34527 94651 34533
rect 94593 34524 94605 34527
rect 94280 34496 94605 34524
rect 94280 34484 94286 34496
rect 94593 34493 94605 34496
rect 94639 34493 94651 34527
rect 94593 34487 94651 34493
rect 88794 34456 88800 34468
rect 59280 34428 59860 34456
rect 60706 34428 88800 34456
rect 9950 34348 9956 34400
rect 10008 34388 10014 34400
rect 27982 34388 27988 34400
rect 10008 34360 27988 34388
rect 10008 34348 10014 34360
rect 27982 34348 27988 34360
rect 28040 34348 28046 34400
rect 28074 34348 28080 34400
rect 28132 34388 28138 34400
rect 33870 34388 33876 34400
rect 28132 34360 33876 34388
rect 28132 34348 28138 34360
rect 33870 34348 33876 34360
rect 33928 34348 33934 34400
rect 33962 34348 33968 34400
rect 34020 34388 34026 34400
rect 41322 34388 41328 34400
rect 34020 34360 41328 34388
rect 34020 34348 34026 34360
rect 41322 34348 41328 34360
rect 41380 34348 41386 34400
rect 41690 34348 41696 34400
rect 41748 34388 41754 34400
rect 52270 34388 52276 34400
rect 41748 34360 52276 34388
rect 41748 34348 41754 34360
rect 52270 34348 52276 34360
rect 52328 34348 52334 34400
rect 52362 34348 52368 34400
rect 52420 34388 52426 34400
rect 60706 34388 60734 34428
rect 88794 34416 88800 34428
rect 88852 34416 88858 34468
rect 52420 34360 60734 34388
rect 52420 34348 52426 34360
rect 67450 34348 67456 34400
rect 67508 34388 67514 34400
rect 69198 34388 69204 34400
rect 67508 34360 69204 34388
rect 67508 34348 67514 34360
rect 69198 34348 69204 34360
rect 69256 34348 69262 34400
rect 69290 34348 69296 34400
rect 69348 34388 69354 34400
rect 90634 34388 90640 34400
rect 69348 34360 90640 34388
rect 69348 34348 69354 34360
rect 90634 34348 90640 34360
rect 90692 34348 90698 34400
rect 1104 34298 98808 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 50326 34298
rect 50378 34246 50390 34298
rect 50442 34246 50454 34298
rect 50506 34246 50518 34298
rect 50570 34246 81046 34298
rect 81098 34246 81110 34298
rect 81162 34246 81174 34298
rect 81226 34246 81238 34298
rect 81290 34246 98808 34298
rect 1104 34224 98808 34246
rect 28074 34184 28080 34196
rect 12406 34156 28080 34184
rect 9950 34048 9956 34060
rect 9911 34020 9956 34048
rect 9950 34008 9956 34020
rect 10008 34008 10014 34060
rect 10321 34051 10379 34057
rect 10321 34017 10333 34051
rect 10367 34048 10379 34051
rect 12406 34048 12434 34156
rect 28074 34144 28080 34156
rect 28132 34144 28138 34196
rect 30466 34144 30472 34196
rect 30524 34184 30530 34196
rect 31478 34184 31484 34196
rect 30524 34156 31484 34184
rect 30524 34144 30530 34156
rect 31478 34144 31484 34156
rect 31536 34184 31542 34196
rect 34790 34184 34796 34196
rect 31536 34156 34796 34184
rect 31536 34144 31542 34156
rect 34790 34144 34796 34156
rect 34848 34144 34854 34196
rect 35250 34144 35256 34196
rect 35308 34184 35314 34196
rect 36354 34184 36360 34196
rect 35308 34156 36360 34184
rect 35308 34144 35314 34156
rect 36354 34144 36360 34156
rect 36412 34144 36418 34196
rect 40494 34184 40500 34196
rect 36464 34156 40500 34184
rect 17865 34119 17923 34125
rect 17865 34085 17877 34119
rect 17911 34116 17923 34119
rect 17911 34088 18736 34116
rect 17911 34085 17923 34088
rect 17865 34079 17923 34085
rect 18708 34060 18736 34088
rect 22830 34076 22836 34128
rect 22888 34116 22894 34128
rect 36464 34116 36492 34156
rect 40494 34144 40500 34156
rect 40552 34144 40558 34196
rect 40954 34144 40960 34196
rect 41012 34184 41018 34196
rect 41414 34184 41420 34196
rect 41012 34156 41420 34184
rect 41012 34144 41018 34156
rect 41414 34144 41420 34156
rect 41472 34144 41478 34196
rect 41506 34144 41512 34196
rect 41564 34184 41570 34196
rect 64782 34184 64788 34196
rect 41564 34156 64788 34184
rect 41564 34144 41570 34156
rect 64782 34144 64788 34156
rect 64840 34144 64846 34196
rect 64966 34144 64972 34196
rect 65024 34184 65030 34196
rect 71041 34187 71099 34193
rect 71041 34184 71053 34187
rect 65024 34156 71053 34184
rect 65024 34144 65030 34156
rect 71041 34153 71053 34156
rect 71087 34153 71099 34187
rect 71041 34147 71099 34153
rect 84838 34144 84844 34196
rect 84896 34184 84902 34196
rect 85482 34184 85488 34196
rect 84896 34156 85488 34184
rect 84896 34144 84902 34156
rect 85482 34144 85488 34156
rect 85540 34144 85546 34196
rect 22888 34088 36492 34116
rect 22888 34076 22894 34088
rect 36538 34076 36544 34128
rect 36596 34116 36602 34128
rect 46934 34116 46940 34128
rect 36596 34088 46940 34116
rect 36596 34076 36602 34088
rect 46934 34076 46940 34088
rect 46992 34076 46998 34128
rect 47302 34076 47308 34128
rect 47360 34116 47366 34128
rect 47360 34088 51120 34116
rect 47360 34076 47366 34088
rect 10367 34020 12434 34048
rect 18417 34051 18475 34057
rect 10367 34017 10379 34020
rect 10321 34011 10379 34017
rect 18417 34017 18429 34051
rect 18463 34017 18475 34051
rect 18690 34048 18696 34060
rect 18651 34020 18696 34048
rect 18417 34011 18475 34017
rect 10413 33983 10471 33989
rect 10413 33949 10425 33983
rect 10459 33980 10471 33983
rect 18230 33980 18236 33992
rect 10459 33952 17908 33980
rect 18191 33952 18236 33980
rect 10459 33949 10471 33952
rect 10413 33943 10471 33949
rect 9769 33915 9827 33921
rect 9769 33881 9781 33915
rect 9815 33912 9827 33915
rect 9950 33912 9956 33924
rect 9815 33884 9956 33912
rect 9815 33881 9827 33884
rect 9769 33875 9827 33881
rect 9950 33872 9956 33884
rect 10008 33872 10014 33924
rect 17880 33844 17908 33952
rect 18230 33940 18236 33952
rect 18288 33940 18294 33992
rect 18432 33980 18460 34011
rect 18690 34008 18696 34020
rect 18748 34008 18754 34060
rect 21634 34048 21640 34060
rect 18800 34020 21640 34048
rect 18800 33980 18828 34020
rect 21634 34008 21640 34020
rect 21692 34008 21698 34060
rect 24854 34008 24860 34060
rect 24912 34048 24918 34060
rect 29362 34048 29368 34060
rect 24912 34020 29368 34048
rect 24912 34008 24918 34020
rect 29362 34008 29368 34020
rect 29420 34008 29426 34060
rect 30374 34008 30380 34060
rect 30432 34048 30438 34060
rect 36446 34048 36452 34060
rect 30432 34020 36452 34048
rect 30432 34008 30438 34020
rect 36446 34008 36452 34020
rect 36504 34008 36510 34060
rect 36630 34008 36636 34060
rect 36688 34048 36694 34060
rect 37826 34048 37832 34060
rect 36688 34020 37832 34048
rect 36688 34008 36694 34020
rect 37826 34008 37832 34020
rect 37884 34008 37890 34060
rect 38654 34008 38660 34060
rect 38712 34048 38718 34060
rect 39942 34048 39948 34060
rect 38712 34020 39948 34048
rect 38712 34008 38718 34020
rect 39942 34008 39948 34020
rect 40000 34008 40006 34060
rect 40402 34008 40408 34060
rect 40460 34048 40466 34060
rect 40460 34020 42196 34048
rect 40460 34008 40466 34020
rect 18432 33952 18828 33980
rect 18874 33940 18880 33992
rect 18932 33980 18938 33992
rect 21545 33983 21603 33989
rect 21545 33980 21557 33983
rect 18932 33952 21557 33980
rect 18932 33940 18938 33952
rect 21545 33949 21557 33952
rect 21591 33949 21603 33983
rect 21818 33980 21824 33992
rect 21779 33952 21824 33980
rect 21545 33943 21603 33949
rect 21818 33940 21824 33952
rect 21876 33940 21882 33992
rect 33962 33980 33968 33992
rect 22848 33952 33968 33980
rect 18506 33872 18512 33924
rect 18564 33912 18570 33924
rect 18601 33915 18659 33921
rect 18601 33912 18613 33915
rect 18564 33884 18613 33912
rect 18564 33872 18570 33884
rect 18601 33881 18613 33884
rect 18647 33881 18659 33915
rect 18601 33875 18659 33881
rect 22848 33844 22876 33952
rect 33962 33940 33968 33952
rect 34020 33940 34026 33992
rect 34146 33940 34152 33992
rect 34204 33980 34210 33992
rect 42061 33983 42119 33989
rect 42061 33980 42073 33983
rect 34204 33952 42073 33980
rect 34204 33940 34210 33952
rect 42061 33949 42073 33952
rect 42107 33949 42119 33983
rect 42168 33980 42196 34020
rect 42242 34008 42248 34060
rect 42300 34048 42306 34060
rect 42426 34048 42432 34060
rect 42300 34020 42345 34048
rect 42387 34020 42432 34048
rect 42300 34008 42306 34020
rect 42426 34008 42432 34020
rect 42484 34008 42490 34060
rect 42521 34051 42579 34057
rect 42521 34017 42533 34051
rect 42567 34048 42579 34051
rect 42610 34048 42616 34060
rect 42567 34020 42616 34048
rect 42567 34017 42579 34020
rect 42521 34011 42579 34017
rect 42610 34008 42616 34020
rect 42668 34008 42674 34060
rect 44266 34008 44272 34060
rect 44324 34048 44330 34060
rect 50890 34048 50896 34060
rect 44324 34020 50896 34048
rect 44324 34008 44330 34020
rect 50890 34008 50896 34020
rect 50948 34008 50954 34060
rect 51092 34048 51120 34088
rect 51166 34076 51172 34128
rect 51224 34116 51230 34128
rect 58158 34116 58164 34128
rect 51224 34088 58164 34116
rect 51224 34076 51230 34088
rect 58158 34076 58164 34088
rect 58216 34076 58222 34128
rect 58618 34076 58624 34128
rect 58676 34116 58682 34128
rect 93397 34119 93455 34125
rect 93397 34116 93409 34119
rect 58676 34088 93409 34116
rect 58676 34076 58682 34088
rect 93397 34085 93409 34088
rect 93443 34085 93455 34119
rect 93397 34079 93455 34085
rect 68462 34048 68468 34060
rect 51092 34020 68468 34048
rect 68462 34008 68468 34020
rect 68520 34008 68526 34060
rect 70397 34051 70455 34057
rect 70397 34017 70409 34051
rect 70443 34048 70455 34051
rect 70670 34048 70676 34060
rect 70443 34020 70676 34048
rect 70443 34017 70455 34020
rect 70397 34011 70455 34017
rect 70670 34008 70676 34020
rect 70728 34008 70734 34060
rect 77754 34048 77760 34060
rect 77715 34020 77760 34048
rect 77754 34008 77760 34020
rect 77812 34008 77818 34060
rect 77846 34008 77852 34060
rect 77904 34048 77910 34060
rect 95418 34048 95424 34060
rect 77904 34020 95424 34048
rect 77904 34008 77910 34020
rect 95418 34008 95424 34020
rect 95476 34008 95482 34060
rect 42168 33952 42288 33980
rect 42061 33943 42119 33949
rect 24762 33872 24768 33924
rect 24820 33912 24826 33924
rect 36538 33912 36544 33924
rect 24820 33884 36544 33912
rect 24820 33872 24826 33884
rect 36538 33872 36544 33884
rect 36596 33872 36602 33924
rect 37734 33872 37740 33924
rect 37792 33912 37798 33924
rect 41138 33912 41144 33924
rect 37792 33884 41144 33912
rect 37792 33872 37798 33884
rect 41138 33872 41144 33884
rect 41196 33872 41202 33924
rect 42260 33912 42288 33952
rect 44450 33940 44456 33992
rect 44508 33980 44514 33992
rect 45462 33980 45468 33992
rect 44508 33952 45468 33980
rect 44508 33940 44514 33952
rect 45462 33940 45468 33952
rect 45520 33940 45526 33992
rect 45554 33940 45560 33992
rect 45612 33980 45618 33992
rect 50982 33980 50988 33992
rect 45612 33952 50988 33980
rect 45612 33940 45618 33952
rect 50982 33940 50988 33952
rect 51040 33940 51046 33992
rect 52270 33940 52276 33992
rect 52328 33980 52334 33992
rect 61654 33980 61660 33992
rect 52328 33952 61660 33980
rect 52328 33940 52334 33952
rect 61654 33940 61660 33952
rect 61712 33980 61718 33992
rect 62022 33980 62028 33992
rect 61712 33952 62028 33980
rect 61712 33940 61718 33952
rect 62022 33940 62028 33952
rect 62080 33940 62086 33992
rect 64782 33940 64788 33992
rect 64840 33980 64846 33992
rect 64840 33952 67634 33980
rect 64840 33940 64846 33952
rect 53098 33912 53104 33924
rect 41386 33884 42196 33912
rect 42260 33884 53104 33912
rect 17880 33816 22876 33844
rect 23109 33847 23167 33853
rect 23109 33813 23121 33847
rect 23155 33844 23167 33847
rect 24578 33844 24584 33856
rect 23155 33816 24584 33844
rect 23155 33813 23167 33816
rect 23109 33807 23167 33813
rect 24578 33804 24584 33816
rect 24636 33804 24642 33856
rect 27617 33847 27675 33853
rect 27617 33813 27629 33847
rect 27663 33844 27675 33847
rect 27893 33847 27951 33853
rect 27893 33844 27905 33847
rect 27663 33816 27905 33844
rect 27663 33813 27675 33816
rect 27617 33807 27675 33813
rect 27893 33813 27905 33816
rect 27939 33844 27951 33847
rect 41386 33844 41414 33884
rect 27939 33816 41414 33844
rect 42168 33844 42196 33884
rect 53098 33872 53104 33884
rect 53156 33872 53162 33924
rect 66898 33912 66904 33924
rect 54772 33884 66904 33912
rect 54772 33844 54800 33884
rect 66898 33872 66904 33884
rect 66956 33872 66962 33924
rect 67606 33912 67634 33952
rect 70578 33940 70584 33992
rect 70636 33980 70642 33992
rect 70765 33983 70823 33989
rect 70765 33980 70777 33983
rect 70636 33952 70777 33980
rect 70636 33940 70642 33952
rect 70765 33949 70777 33952
rect 70811 33949 70823 33983
rect 70765 33943 70823 33949
rect 72418 33940 72424 33992
rect 72476 33980 72482 33992
rect 78033 33983 78091 33989
rect 78033 33980 78045 33983
rect 72476 33952 78045 33980
rect 72476 33940 72482 33952
rect 78033 33949 78045 33952
rect 78079 33949 78091 33983
rect 94777 33983 94835 33989
rect 94777 33980 94789 33983
rect 78033 33943 78091 33949
rect 93826 33952 94789 33980
rect 72970 33912 72976 33924
rect 67606 33884 72976 33912
rect 72970 33872 72976 33884
rect 73028 33912 73034 33924
rect 75546 33912 75552 33924
rect 73028 33884 75552 33912
rect 73028 33872 73034 33884
rect 75546 33872 75552 33884
rect 75604 33872 75610 33924
rect 42168 33816 54800 33844
rect 27939 33813 27951 33816
rect 27893 33807 27951 33813
rect 55030 33804 55036 33856
rect 55088 33844 55094 33856
rect 58066 33844 58072 33856
rect 55088 33816 58072 33844
rect 55088 33804 55094 33816
rect 58066 33804 58072 33816
rect 58124 33804 58130 33856
rect 59354 33804 59360 33856
rect 59412 33844 59418 33856
rect 63218 33844 63224 33856
rect 59412 33816 63224 33844
rect 59412 33804 59418 33816
rect 63218 33804 63224 33816
rect 63276 33804 63282 33856
rect 63310 33804 63316 33856
rect 63368 33844 63374 33856
rect 70535 33847 70593 33853
rect 70535 33844 70547 33847
rect 63368 33816 70547 33844
rect 63368 33804 63374 33816
rect 70535 33813 70547 33816
rect 70581 33813 70593 33847
rect 70535 33807 70593 33813
rect 70673 33847 70731 33853
rect 70673 33813 70685 33847
rect 70719 33844 70731 33847
rect 70762 33844 70768 33856
rect 70719 33816 70768 33844
rect 70719 33813 70731 33816
rect 70673 33807 70731 33813
rect 70762 33804 70768 33816
rect 70820 33804 70826 33856
rect 93210 33844 93216 33856
rect 93171 33816 93216 33844
rect 93210 33804 93216 33816
rect 93268 33844 93274 33856
rect 93826 33844 93854 33952
rect 94777 33949 94789 33952
rect 94823 33949 94835 33983
rect 94777 33943 94835 33949
rect 95053 33983 95111 33989
rect 95053 33949 95065 33983
rect 95099 33980 95111 33983
rect 95142 33980 95148 33992
rect 95099 33952 95148 33980
rect 95099 33949 95111 33952
rect 95053 33943 95111 33949
rect 95142 33940 95148 33952
rect 95200 33940 95206 33992
rect 93268 33816 93854 33844
rect 93268 33804 93274 33816
rect 1104 33754 98808 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 65686 33754
rect 65738 33702 65750 33754
rect 65802 33702 65814 33754
rect 65866 33702 65878 33754
rect 65930 33702 96406 33754
rect 96458 33702 96470 33754
rect 96522 33702 96534 33754
rect 96586 33702 96598 33754
rect 96650 33702 98808 33754
rect 1104 33680 98808 33702
rect 17678 33600 17684 33652
rect 17736 33640 17742 33652
rect 34146 33640 34152 33652
rect 17736 33612 34152 33640
rect 17736 33600 17742 33612
rect 34146 33600 34152 33612
rect 34204 33600 34210 33652
rect 34238 33600 34244 33652
rect 34296 33640 34302 33652
rect 34296 33612 41092 33640
rect 34296 33600 34302 33612
rect 19613 33575 19671 33581
rect 19613 33541 19625 33575
rect 19659 33572 19671 33575
rect 19659 33544 21220 33572
rect 19659 33541 19671 33544
rect 19613 33535 19671 33541
rect 17586 33504 17592 33516
rect 17547 33476 17592 33504
rect 17586 33464 17592 33476
rect 17644 33464 17650 33516
rect 19886 33464 19892 33516
rect 19944 33504 19950 33516
rect 19944 33476 20668 33504
rect 19944 33464 19950 33476
rect 17313 33439 17371 33445
rect 17313 33405 17325 33439
rect 17359 33436 17371 33439
rect 18874 33436 18880 33448
rect 17359 33408 18880 33436
rect 17359 33405 17371 33408
rect 17313 33399 17371 33405
rect 18874 33396 18880 33408
rect 18932 33436 18938 33448
rect 19150 33436 19156 33448
rect 18932 33408 19156 33436
rect 18932 33396 18938 33408
rect 19150 33396 19156 33408
rect 19208 33396 19214 33448
rect 20640 33445 20668 33476
rect 20257 33439 20315 33445
rect 20257 33405 20269 33439
rect 20303 33405 20315 33439
rect 20257 33399 20315 33405
rect 20625 33439 20683 33445
rect 20625 33405 20637 33439
rect 20671 33405 20683 33439
rect 20625 33399 20683 33405
rect 20717 33439 20775 33445
rect 20717 33405 20729 33439
rect 20763 33405 20775 33439
rect 20990 33436 20996 33448
rect 20951 33408 20996 33436
rect 20717 33399 20775 33405
rect 20272 33368 20300 33399
rect 20530 33368 20536 33380
rect 20272 33340 20536 33368
rect 20530 33328 20536 33340
rect 20588 33328 20594 33380
rect 20732 33368 20760 33399
rect 20990 33396 20996 33408
rect 21048 33396 21054 33448
rect 21192 33445 21220 33544
rect 27798 33532 27804 33584
rect 27856 33572 27862 33584
rect 30190 33572 30196 33584
rect 27856 33544 30196 33572
rect 27856 33532 27862 33544
rect 30190 33532 30196 33544
rect 30248 33532 30254 33584
rect 40126 33572 40132 33584
rect 35176 33544 40132 33572
rect 22066 33476 30880 33504
rect 21177 33439 21235 33445
rect 21177 33405 21189 33439
rect 21223 33436 21235 33439
rect 22066 33436 22094 33476
rect 24486 33436 24492 33448
rect 21223 33408 22094 33436
rect 24447 33408 24492 33436
rect 21223 33405 21235 33408
rect 21177 33399 21235 33405
rect 24486 33396 24492 33408
rect 24544 33396 24550 33448
rect 30190 33436 30196 33448
rect 30151 33408 30196 33436
rect 30190 33396 30196 33408
rect 30248 33396 30254 33448
rect 30282 33396 30288 33448
rect 30340 33436 30346 33448
rect 30466 33445 30472 33448
rect 30377 33439 30435 33445
rect 30377 33436 30389 33439
rect 30340 33408 30389 33436
rect 30340 33396 30346 33408
rect 30377 33405 30389 33408
rect 30423 33405 30435 33439
rect 30377 33399 30435 33405
rect 30465 33399 30472 33445
rect 30524 33436 30530 33448
rect 30607 33439 30665 33445
rect 30524 33408 30565 33436
rect 30466 33396 30472 33399
rect 30524 33396 30530 33408
rect 30607 33405 30619 33439
rect 30653 33436 30665 33439
rect 30852 33436 30880 33476
rect 30926 33464 30932 33516
rect 30984 33504 30990 33516
rect 35176 33504 35204 33544
rect 40126 33532 40132 33544
rect 40184 33532 40190 33584
rect 41064 33572 41092 33612
rect 41138 33600 41144 33652
rect 41196 33640 41202 33652
rect 67818 33640 67824 33652
rect 41196 33612 67824 33640
rect 41196 33600 41202 33612
rect 67818 33600 67824 33612
rect 67876 33600 67882 33652
rect 70118 33600 70124 33652
rect 70176 33640 70182 33652
rect 70302 33640 70308 33652
rect 70176 33612 70308 33640
rect 70176 33600 70182 33612
rect 70302 33600 70308 33612
rect 70360 33600 70366 33652
rect 72234 33572 72240 33584
rect 41064 33544 72240 33572
rect 72234 33532 72240 33544
rect 72292 33532 72298 33584
rect 30984 33476 35204 33504
rect 35268 33476 41276 33504
rect 30984 33464 30990 33476
rect 35268 33436 35296 33476
rect 30653 33408 30788 33436
rect 30852 33408 35296 33436
rect 30653 33405 30665 33408
rect 30607 33399 30665 33405
rect 21358 33368 21364 33380
rect 20732 33340 21364 33368
rect 21358 33328 21364 33340
rect 21416 33328 21422 33380
rect 22094 33328 22100 33380
rect 22152 33368 22158 33380
rect 24857 33371 24915 33377
rect 24857 33368 24869 33371
rect 22152 33340 24869 33368
rect 22152 33328 22158 33340
rect 24857 33337 24869 33340
rect 24903 33368 24915 33371
rect 25314 33368 25320 33380
rect 24903 33340 25320 33368
rect 24903 33337 24915 33340
rect 24857 33331 24915 33337
rect 25314 33328 25320 33340
rect 25372 33328 25378 33380
rect 27982 33328 27988 33380
rect 28040 33368 28046 33380
rect 28810 33368 28816 33380
rect 28040 33340 28816 33368
rect 28040 33328 28046 33340
rect 28810 33328 28816 33340
rect 28868 33368 28874 33380
rect 30006 33368 30012 33380
rect 28868 33340 30012 33368
rect 28868 33328 28874 33340
rect 30006 33328 30012 33340
rect 30064 33328 30070 33380
rect 30760 33368 30788 33408
rect 36446 33396 36452 33448
rect 36504 33436 36510 33448
rect 39945 33439 40003 33445
rect 39945 33436 39957 33439
rect 36504 33408 39957 33436
rect 36504 33396 36510 33408
rect 39945 33405 39957 33408
rect 39991 33405 40003 33439
rect 39945 33399 40003 33405
rect 32490 33368 32496 33380
rect 30760 33340 32496 33368
rect 32490 33328 32496 33340
rect 32548 33328 32554 33380
rect 39960 33368 39988 33399
rect 40034 33396 40040 33448
rect 40092 33436 40098 33448
rect 40129 33439 40187 33445
rect 40129 33436 40141 33439
rect 40092 33408 40141 33436
rect 40092 33396 40098 33408
rect 40129 33405 40141 33408
rect 40175 33405 40187 33439
rect 40405 33439 40463 33445
rect 40405 33436 40417 33439
rect 40129 33399 40187 33405
rect 40236 33408 40417 33436
rect 40236 33368 40264 33408
rect 40405 33405 40417 33408
rect 40451 33405 40463 33439
rect 41248 33436 41276 33476
rect 41322 33464 41328 33516
rect 41380 33504 41386 33516
rect 45554 33504 45560 33516
rect 41380 33476 45560 33504
rect 41380 33464 41386 33476
rect 45554 33464 45560 33476
rect 45612 33464 45618 33516
rect 45646 33464 45652 33516
rect 45704 33504 45710 33516
rect 49142 33504 49148 33516
rect 45704 33476 49148 33504
rect 45704 33464 45710 33476
rect 49142 33464 49148 33476
rect 49200 33464 49206 33516
rect 54478 33504 54484 33516
rect 49252 33476 54484 33504
rect 49050 33436 49056 33448
rect 41248 33408 49056 33436
rect 40405 33399 40463 33405
rect 49050 33396 49056 33408
rect 49108 33396 49114 33448
rect 49252 33445 49280 33476
rect 54478 33464 54484 33476
rect 54536 33464 54542 33516
rect 56134 33464 56140 33516
rect 56192 33504 56198 33516
rect 60366 33504 60372 33516
rect 56192 33476 60372 33504
rect 56192 33464 56198 33476
rect 60366 33464 60372 33476
rect 60424 33464 60430 33516
rect 60829 33507 60887 33513
rect 60829 33473 60841 33507
rect 60875 33504 60887 33507
rect 61378 33504 61384 33516
rect 60875 33476 61384 33504
rect 60875 33473 60887 33476
rect 60829 33467 60887 33473
rect 61378 33464 61384 33476
rect 61436 33464 61442 33516
rect 62022 33464 62028 33516
rect 62080 33504 62086 33516
rect 69290 33504 69296 33516
rect 62080 33476 69296 33504
rect 62080 33464 62086 33476
rect 69290 33464 69296 33476
rect 69348 33464 69354 33516
rect 49237 33439 49295 33445
rect 49237 33405 49249 33439
rect 49283 33405 49295 33439
rect 49237 33399 49295 33405
rect 53098 33396 53104 33448
rect 53156 33436 53162 33448
rect 59354 33436 59360 33448
rect 53156 33408 58848 33436
rect 59315 33408 59360 33436
rect 53156 33396 53162 33408
rect 39960 33340 40264 33368
rect 41386 33340 41644 33368
rect 18690 33300 18696 33312
rect 18651 33272 18696 33300
rect 18690 33260 18696 33272
rect 18748 33260 18754 33312
rect 19797 33303 19855 33309
rect 19797 33269 19809 33303
rect 19843 33300 19855 33303
rect 19889 33303 19947 33309
rect 19889 33300 19901 33303
rect 19843 33272 19901 33300
rect 19843 33269 19855 33272
rect 19797 33263 19855 33269
rect 19889 33269 19901 33272
rect 19935 33300 19947 33303
rect 20073 33303 20131 33309
rect 20073 33300 20085 33303
rect 19935 33272 20085 33300
rect 19935 33269 19947 33272
rect 19889 33263 19947 33269
rect 20073 33269 20085 33272
rect 20119 33300 20131 33303
rect 21453 33303 21511 33309
rect 21453 33300 21465 33303
rect 20119 33272 21465 33300
rect 20119 33269 20131 33272
rect 20073 33263 20131 33269
rect 21453 33269 21465 33272
rect 21499 33300 21511 33303
rect 21729 33303 21787 33309
rect 21729 33300 21741 33303
rect 21499 33272 21741 33300
rect 21499 33269 21511 33272
rect 21453 33263 21511 33269
rect 21729 33269 21741 33272
rect 21775 33300 21787 33303
rect 21913 33303 21971 33309
rect 21913 33300 21925 33303
rect 21775 33272 21925 33300
rect 21775 33269 21787 33272
rect 21729 33263 21787 33269
rect 21913 33269 21925 33272
rect 21959 33300 21971 33303
rect 22281 33303 22339 33309
rect 22281 33300 22293 33303
rect 21959 33272 22293 33300
rect 21959 33269 21971 33272
rect 21913 33263 21971 33269
rect 22281 33269 22293 33272
rect 22327 33300 22339 33303
rect 30466 33300 30472 33312
rect 22327 33272 30472 33300
rect 22327 33269 22339 33272
rect 22281 33263 22339 33269
rect 30466 33260 30472 33272
rect 30524 33260 30530 33312
rect 30742 33300 30748 33312
rect 30703 33272 30748 33300
rect 30742 33260 30748 33272
rect 30800 33260 30806 33312
rect 34790 33260 34796 33312
rect 34848 33300 34854 33312
rect 37918 33300 37924 33312
rect 34848 33272 37924 33300
rect 34848 33260 34854 33272
rect 37918 33260 37924 33272
rect 37976 33260 37982 33312
rect 38010 33260 38016 33312
rect 38068 33300 38074 33312
rect 41386 33300 41414 33340
rect 38068 33272 41414 33300
rect 41616 33300 41644 33340
rect 41690 33328 41696 33380
rect 41748 33368 41754 33380
rect 41785 33371 41843 33377
rect 41785 33368 41797 33371
rect 41748 33340 41797 33368
rect 41748 33328 41754 33340
rect 41785 33337 41797 33340
rect 41831 33368 41843 33371
rect 42702 33368 42708 33380
rect 41831 33340 42708 33368
rect 41831 33337 41843 33340
rect 41785 33331 41843 33337
rect 42702 33328 42708 33340
rect 42760 33328 42766 33380
rect 49510 33368 49516 33380
rect 49471 33340 49516 33368
rect 49510 33328 49516 33340
rect 49568 33328 49574 33380
rect 49602 33328 49608 33380
rect 49660 33368 49666 33380
rect 51074 33368 51080 33380
rect 49660 33340 51080 33368
rect 49660 33328 49666 33340
rect 51074 33328 51080 33340
rect 51132 33328 51138 33380
rect 55306 33328 55312 33380
rect 55364 33368 55370 33380
rect 58710 33368 58716 33380
rect 55364 33340 58716 33368
rect 55364 33328 55370 33340
rect 58710 33328 58716 33340
rect 58768 33328 58774 33380
rect 58820 33368 58848 33408
rect 59354 33396 59360 33408
rect 59412 33396 59418 33448
rect 60274 33396 60280 33448
rect 60332 33436 60338 33448
rect 60461 33439 60519 33445
rect 60461 33436 60473 33439
rect 60332 33408 60473 33436
rect 60332 33396 60338 33408
rect 60461 33405 60473 33408
rect 60507 33405 60519 33439
rect 60461 33399 60519 33405
rect 60609 33439 60667 33445
rect 60609 33405 60621 33439
rect 60655 33405 60667 33439
rect 60734 33436 60740 33448
rect 60695 33408 60740 33436
rect 60609 33399 60667 33405
rect 59446 33368 59452 33380
rect 58820 33340 59452 33368
rect 59446 33328 59452 33340
rect 59504 33328 59510 33380
rect 59722 33368 59728 33380
rect 59683 33340 59728 33368
rect 59722 33328 59728 33340
rect 59780 33328 59786 33380
rect 60366 33328 60372 33380
rect 60424 33368 60430 33380
rect 60624 33368 60652 33399
rect 60734 33396 60740 33408
rect 60792 33396 60798 33448
rect 60918 33396 60924 33448
rect 60976 33445 60982 33448
rect 60976 33439 61025 33445
rect 60976 33405 60979 33439
rect 61013 33405 61025 33439
rect 60976 33399 61025 33405
rect 60976 33396 60982 33399
rect 61286 33396 61292 33448
rect 61344 33436 61350 33448
rect 84838 33436 84844 33448
rect 61344 33408 84844 33436
rect 61344 33396 61350 33408
rect 84838 33396 84844 33408
rect 84896 33396 84902 33448
rect 60424 33340 60652 33368
rect 60424 33328 60430 33340
rect 61470 33328 61476 33380
rect 61528 33368 61534 33380
rect 61528 33340 70394 33368
rect 61528 33328 61534 33340
rect 60734 33300 60740 33312
rect 41616 33272 60740 33300
rect 38068 33260 38074 33272
rect 60734 33260 60740 33272
rect 60792 33260 60798 33312
rect 61102 33300 61108 33312
rect 61063 33272 61108 33300
rect 61102 33260 61108 33272
rect 61160 33260 61166 33312
rect 63218 33260 63224 33312
rect 63276 33300 63282 33312
rect 65978 33300 65984 33312
rect 63276 33272 65984 33300
rect 63276 33260 63282 33272
rect 65978 33260 65984 33272
rect 66036 33260 66042 33312
rect 70366 33300 70394 33340
rect 83826 33300 83832 33312
rect 70366 33272 83832 33300
rect 83826 33260 83832 33272
rect 83884 33260 83890 33312
rect 1104 33210 98808 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 50326 33210
rect 50378 33158 50390 33210
rect 50442 33158 50454 33210
rect 50506 33158 50518 33210
rect 50570 33158 81046 33210
rect 81098 33158 81110 33210
rect 81162 33158 81174 33210
rect 81226 33158 81238 33210
rect 81290 33158 98808 33210
rect 1104 33136 98808 33158
rect 16758 33056 16764 33108
rect 16816 33096 16822 33108
rect 90634 33096 90640 33108
rect 16816 33068 80054 33096
rect 90595 33068 90640 33096
rect 16816 33056 16822 33068
rect 22186 32988 22192 33040
rect 22244 33028 22250 33040
rect 38930 33028 38936 33040
rect 22244 33000 38936 33028
rect 22244 32988 22250 33000
rect 38930 32988 38936 33000
rect 38988 32988 38994 33040
rect 42150 33028 42156 33040
rect 39408 33000 42156 33028
rect 16666 32920 16672 32972
rect 16724 32960 16730 32972
rect 22002 32960 22008 32972
rect 16724 32932 22008 32960
rect 16724 32920 16730 32932
rect 22002 32920 22008 32932
rect 22060 32920 22066 32972
rect 22097 32963 22155 32969
rect 22097 32929 22109 32963
rect 22143 32960 22155 32963
rect 22370 32960 22376 32972
rect 22143 32932 22376 32960
rect 22143 32929 22155 32932
rect 22097 32923 22155 32929
rect 22370 32920 22376 32932
rect 22428 32920 22434 32972
rect 38286 32960 38292 32972
rect 22480 32932 38292 32960
rect 16850 32852 16856 32904
rect 16908 32892 16914 32904
rect 22480 32892 22508 32932
rect 38286 32920 38292 32932
rect 38344 32920 38350 32972
rect 38746 32920 38752 32972
rect 38804 32960 38810 32972
rect 39025 32963 39083 32969
rect 39025 32960 39037 32963
rect 38804 32932 39037 32960
rect 38804 32920 38810 32932
rect 39025 32929 39037 32932
rect 39071 32929 39083 32963
rect 39025 32923 39083 32929
rect 39209 32963 39267 32969
rect 39209 32929 39221 32963
rect 39255 32929 39267 32963
rect 39209 32923 39267 32929
rect 39301 32963 39359 32969
rect 39301 32929 39313 32963
rect 39347 32960 39359 32963
rect 39408 32960 39436 33000
rect 42150 32988 42156 33000
rect 42208 32988 42214 33040
rect 42426 32988 42432 33040
rect 42484 33028 42490 33040
rect 42484 33000 46980 33028
rect 42484 32988 42490 33000
rect 39347 32932 39436 32960
rect 39347 32929 39359 32932
rect 39301 32923 39359 32929
rect 22646 32892 22652 32904
rect 16908 32864 22508 32892
rect 22607 32864 22652 32892
rect 16908 32852 16914 32864
rect 22646 32852 22652 32864
rect 22704 32852 22710 32904
rect 26878 32852 26884 32904
rect 26936 32892 26942 32904
rect 35434 32892 35440 32904
rect 26936 32864 35440 32892
rect 26936 32852 26942 32864
rect 35434 32852 35440 32864
rect 35492 32852 35498 32904
rect 38838 32852 38844 32904
rect 38896 32892 38902 32904
rect 39224 32892 39252 32923
rect 39482 32920 39488 32972
rect 39540 32960 39546 32972
rect 39577 32963 39635 32969
rect 39577 32960 39589 32963
rect 39540 32932 39589 32960
rect 39540 32920 39546 32932
rect 39577 32929 39589 32932
rect 39623 32929 39635 32963
rect 42058 32960 42064 32972
rect 42019 32932 42064 32960
rect 39577 32923 39635 32929
rect 42058 32920 42064 32932
rect 42116 32920 42122 32972
rect 46952 32969 46980 33000
rect 49326 32988 49332 33040
rect 49384 33028 49390 33040
rect 71774 33028 71780 33040
rect 49384 33000 71780 33028
rect 49384 32988 49390 33000
rect 71774 32988 71780 33000
rect 71832 32988 71838 33040
rect 80026 33028 80054 33068
rect 90634 33056 90640 33068
rect 90692 33056 90698 33108
rect 95510 33028 95516 33040
rect 80026 33000 95516 33028
rect 95510 32988 95516 33000
rect 95568 32988 95574 33040
rect 42245 32963 42303 32969
rect 42245 32929 42257 32963
rect 42291 32929 42303 32963
rect 42245 32923 42303 32929
rect 42337 32963 42395 32969
rect 42337 32929 42349 32963
rect 42383 32960 42395 32963
rect 46937 32963 46995 32969
rect 42383 32932 42472 32960
rect 42383 32929 42395 32932
rect 42337 32923 42395 32929
rect 39390 32892 39396 32904
rect 38896 32864 39252 32892
rect 39351 32864 39396 32892
rect 38896 32852 38902 32864
rect 39390 32852 39396 32864
rect 39448 32852 39454 32904
rect 40494 32852 40500 32904
rect 40552 32892 40558 32904
rect 42260 32892 42288 32923
rect 40552 32864 42288 32892
rect 40552 32852 40558 32864
rect 6457 32827 6515 32833
rect 6457 32793 6469 32827
rect 6503 32824 6515 32827
rect 6733 32827 6791 32833
rect 6733 32824 6745 32827
rect 6503 32796 6745 32824
rect 6503 32793 6515 32796
rect 6457 32787 6515 32793
rect 6733 32793 6745 32796
rect 6779 32824 6791 32827
rect 6779 32796 13860 32824
rect 6779 32793 6791 32796
rect 6733 32787 6791 32793
rect 13357 32759 13415 32765
rect 13357 32725 13369 32759
rect 13403 32756 13415 32759
rect 13630 32756 13636 32768
rect 13403 32728 13636 32756
rect 13403 32725 13415 32728
rect 13357 32719 13415 32725
rect 13630 32716 13636 32728
rect 13688 32716 13694 32768
rect 13832 32756 13860 32796
rect 13998 32784 14004 32836
rect 14056 32824 14062 32836
rect 21266 32824 21272 32836
rect 14056 32796 21272 32824
rect 14056 32784 14062 32796
rect 21266 32784 21272 32796
rect 21324 32784 21330 32836
rect 22370 32784 22376 32836
rect 22428 32824 22434 32836
rect 26050 32824 26056 32836
rect 22428 32796 26056 32824
rect 22428 32784 22434 32796
rect 26050 32784 26056 32796
rect 26108 32784 26114 32836
rect 29362 32784 29368 32836
rect 29420 32824 29426 32836
rect 39574 32824 39580 32836
rect 29420 32796 39580 32824
rect 29420 32784 29426 32796
rect 39574 32784 39580 32796
rect 39632 32784 39638 32836
rect 39761 32827 39819 32833
rect 39761 32793 39773 32827
rect 39807 32824 39819 32827
rect 39807 32796 42288 32824
rect 39807 32793 39819 32796
rect 39761 32787 39819 32793
rect 32398 32756 32404 32768
rect 13832 32728 32404 32756
rect 32398 32716 32404 32728
rect 32456 32716 32462 32768
rect 32582 32716 32588 32768
rect 32640 32756 32646 32768
rect 38654 32756 38660 32768
rect 32640 32728 38660 32756
rect 32640 32716 32646 32728
rect 38654 32716 38660 32728
rect 38712 32716 38718 32768
rect 38838 32756 38844 32768
rect 38799 32728 38844 32756
rect 38838 32716 38844 32728
rect 38896 32716 38902 32768
rect 39942 32716 39948 32768
rect 40000 32756 40006 32768
rect 41877 32759 41935 32765
rect 41877 32756 41889 32759
rect 40000 32728 41889 32756
rect 40000 32716 40006 32728
rect 41877 32725 41889 32728
rect 41923 32725 41935 32759
rect 42260 32756 42288 32796
rect 42334 32784 42340 32836
rect 42392 32824 42398 32836
rect 42444 32824 42472 32932
rect 46937 32929 46949 32963
rect 46983 32929 46995 32963
rect 46937 32923 46995 32929
rect 47044 32932 50936 32960
rect 42794 32852 42800 32904
rect 42852 32892 42858 32904
rect 47044 32892 47072 32932
rect 47210 32892 47216 32904
rect 42852 32864 47072 32892
rect 47171 32864 47216 32892
rect 42852 32852 42858 32864
rect 47210 32852 47216 32864
rect 47268 32852 47274 32904
rect 47302 32852 47308 32904
rect 47360 32892 47366 32904
rect 49694 32892 49700 32904
rect 47360 32864 49700 32892
rect 47360 32852 47366 32864
rect 49694 32852 49700 32864
rect 49752 32852 49758 32904
rect 42392 32796 42472 32824
rect 42628 32796 43300 32824
rect 42392 32784 42398 32796
rect 42628 32756 42656 32796
rect 42260 32728 42656 32756
rect 41877 32719 41935 32725
rect 42702 32716 42708 32768
rect 42760 32756 42766 32768
rect 43162 32756 43168 32768
rect 42760 32728 43168 32756
rect 42760 32716 42766 32728
rect 43162 32716 43168 32728
rect 43220 32716 43226 32768
rect 43272 32756 43300 32796
rect 46566 32784 46572 32836
rect 46624 32824 46630 32836
rect 50614 32824 50620 32836
rect 46624 32796 50620 32824
rect 46624 32784 46630 32796
rect 50614 32784 50620 32796
rect 50672 32784 50678 32836
rect 50908 32824 50936 32932
rect 59722 32920 59728 32972
rect 59780 32960 59786 32972
rect 90453 32963 90511 32969
rect 90453 32960 90465 32963
rect 59780 32932 90465 32960
rect 59780 32920 59786 32932
rect 90453 32929 90465 32932
rect 90499 32929 90511 32963
rect 90453 32923 90511 32929
rect 90729 32963 90787 32969
rect 90729 32929 90741 32963
rect 90775 32960 90787 32963
rect 90818 32960 90824 32972
rect 90775 32932 90824 32960
rect 90775 32929 90787 32932
rect 90729 32923 90787 32929
rect 90818 32920 90824 32932
rect 90876 32920 90882 32972
rect 56042 32852 56048 32904
rect 56100 32892 56106 32904
rect 60918 32892 60924 32904
rect 56100 32864 60924 32892
rect 56100 32852 56106 32864
rect 60918 32852 60924 32864
rect 60976 32892 60982 32904
rect 64322 32892 64328 32904
rect 60976 32864 64328 32892
rect 60976 32852 60982 32864
rect 64322 32852 64328 32864
rect 64380 32892 64386 32904
rect 68922 32892 68928 32904
rect 64380 32864 68928 32892
rect 64380 32852 64386 32864
rect 68922 32852 68928 32864
rect 68980 32852 68986 32904
rect 58526 32824 58532 32836
rect 50908 32796 58532 32824
rect 58526 32784 58532 32796
rect 58584 32784 58590 32836
rect 59262 32784 59268 32836
rect 59320 32824 59326 32836
rect 70578 32824 70584 32836
rect 59320 32796 70584 32824
rect 59320 32784 59326 32796
rect 70578 32784 70584 32796
rect 70636 32784 70642 32836
rect 61838 32756 61844 32768
rect 43272 32728 61844 32756
rect 61838 32716 61844 32728
rect 61896 32716 61902 32768
rect 68830 32716 68836 32768
rect 68888 32756 68894 32768
rect 69658 32756 69664 32768
rect 68888 32728 69664 32756
rect 68888 32716 68894 32728
rect 69658 32716 69664 32728
rect 69716 32716 69722 32768
rect 90082 32716 90088 32768
rect 90140 32756 90146 32768
rect 90269 32759 90327 32765
rect 90269 32756 90281 32759
rect 90140 32728 90281 32756
rect 90140 32716 90146 32728
rect 90269 32725 90281 32728
rect 90315 32725 90327 32759
rect 90269 32719 90327 32725
rect 1104 32666 98808 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 65686 32666
rect 65738 32614 65750 32666
rect 65802 32614 65814 32666
rect 65866 32614 65878 32666
rect 65930 32614 96406 32666
rect 96458 32614 96470 32666
rect 96522 32614 96534 32666
rect 96586 32614 96598 32666
rect 96650 32614 98808 32666
rect 1104 32592 98808 32614
rect 13630 32512 13636 32564
rect 13688 32552 13694 32564
rect 26878 32552 26884 32564
rect 13688 32524 26884 32552
rect 13688 32512 13694 32524
rect 26878 32512 26884 32524
rect 26936 32512 26942 32564
rect 26970 32512 26976 32564
rect 27028 32552 27034 32564
rect 30374 32552 30380 32564
rect 27028 32524 30380 32552
rect 27028 32512 27034 32524
rect 30374 32512 30380 32524
rect 30432 32512 30438 32564
rect 31573 32555 31631 32561
rect 31573 32521 31585 32555
rect 31619 32552 31631 32555
rect 31662 32552 31668 32564
rect 31619 32524 31668 32552
rect 31619 32521 31631 32524
rect 31573 32515 31631 32521
rect 31662 32512 31668 32524
rect 31720 32552 31726 32564
rect 31849 32555 31907 32561
rect 31849 32552 31861 32555
rect 31720 32524 31861 32552
rect 31720 32512 31726 32524
rect 31849 32521 31861 32524
rect 31895 32521 31907 32555
rect 31849 32515 31907 32521
rect 32493 32555 32551 32561
rect 32493 32521 32505 32555
rect 32539 32552 32551 32555
rect 42981 32555 43039 32561
rect 42981 32552 42993 32555
rect 32539 32524 42993 32552
rect 32539 32521 32551 32524
rect 32493 32515 32551 32521
rect 42981 32521 42993 32524
rect 43027 32521 43039 32555
rect 42981 32515 43039 32521
rect 43162 32512 43168 32564
rect 43220 32552 43226 32564
rect 55030 32552 55036 32564
rect 43220 32524 55036 32552
rect 43220 32512 43226 32524
rect 55030 32512 55036 32524
rect 55088 32512 55094 32564
rect 58158 32512 58164 32564
rect 58216 32552 58222 32564
rect 85758 32552 85764 32564
rect 58216 32524 85764 32552
rect 58216 32512 58222 32524
rect 85758 32512 85764 32524
rect 85816 32512 85822 32564
rect 13449 32487 13507 32493
rect 13449 32453 13461 32487
rect 13495 32484 13507 32487
rect 13725 32487 13783 32493
rect 13725 32484 13737 32487
rect 13495 32456 13737 32484
rect 13495 32453 13507 32456
rect 13449 32447 13507 32453
rect 13725 32453 13737 32456
rect 13771 32484 13783 32487
rect 13998 32484 14004 32496
rect 13771 32456 14004 32484
rect 13771 32453 13783 32456
rect 13725 32447 13783 32453
rect 13998 32444 14004 32456
rect 14056 32444 14062 32496
rect 23014 32484 23020 32496
rect 22975 32456 23020 32484
rect 23014 32444 23020 32456
rect 23072 32444 23078 32496
rect 25406 32444 25412 32496
rect 25464 32484 25470 32496
rect 39942 32484 39948 32496
rect 25464 32456 39948 32484
rect 25464 32444 25470 32456
rect 39942 32444 39948 32456
rect 40000 32444 40006 32496
rect 41248 32456 56732 32484
rect 12250 32376 12256 32428
rect 12308 32416 12314 32428
rect 21910 32416 21916 32428
rect 12308 32388 21916 32416
rect 12308 32376 12314 32388
rect 21910 32376 21916 32388
rect 21968 32376 21974 32428
rect 22465 32419 22523 32425
rect 22465 32385 22477 32419
rect 22511 32416 22523 32419
rect 41248 32416 41276 32456
rect 22511 32388 24716 32416
rect 22511 32385 22523 32388
rect 22465 32379 22523 32385
rect 13814 32308 13820 32360
rect 13872 32348 13878 32360
rect 13998 32348 14004 32360
rect 13872 32320 14004 32348
rect 13872 32308 13878 32320
rect 13998 32308 14004 32320
rect 14056 32308 14062 32360
rect 22094 32348 22100 32360
rect 15948 32320 22100 32348
rect 11606 32240 11612 32292
rect 11664 32280 11670 32292
rect 15948 32280 15976 32320
rect 22094 32308 22100 32320
rect 22152 32308 22158 32360
rect 22557 32351 22615 32357
rect 22557 32348 22569 32351
rect 22480 32320 22569 32348
rect 22480 32292 22508 32320
rect 22557 32317 22569 32320
rect 22603 32317 22615 32351
rect 22557 32311 22615 32317
rect 11664 32252 15976 32280
rect 11664 32240 11670 32252
rect 16022 32240 16028 32292
rect 16080 32280 16086 32292
rect 22370 32280 22376 32292
rect 16080 32252 22376 32280
rect 16080 32240 16086 32252
rect 22370 32240 22376 32252
rect 22428 32240 22434 32292
rect 22462 32240 22468 32292
rect 22520 32240 22526 32292
rect 17310 32172 17316 32224
rect 17368 32212 17374 32224
rect 22278 32212 22284 32224
rect 17368 32184 22284 32212
rect 17368 32172 17374 32184
rect 22278 32172 22284 32184
rect 22336 32172 22342 32224
rect 22649 32215 22707 32221
rect 22649 32181 22661 32215
rect 22695 32212 22707 32215
rect 22756 32212 22784 32388
rect 22833 32351 22891 32357
rect 22833 32317 22845 32351
rect 22879 32317 22891 32351
rect 22833 32311 22891 32317
rect 22695 32184 22784 32212
rect 22848 32212 22876 32311
rect 24688 32280 24716 32388
rect 27908 32388 41276 32416
rect 27908 32360 27936 32388
rect 41966 32376 41972 32428
rect 42024 32416 42030 32428
rect 53742 32416 53748 32428
rect 42024 32388 53748 32416
rect 42024 32376 42030 32388
rect 53742 32376 53748 32388
rect 53800 32376 53806 32428
rect 56597 32419 56655 32425
rect 56597 32416 56609 32419
rect 53852 32388 56609 32416
rect 27890 32348 27896 32360
rect 27803 32320 27896 32348
rect 27890 32308 27896 32320
rect 27948 32308 27954 32360
rect 31389 32351 31447 32357
rect 31389 32348 31401 32351
rect 28000 32320 31401 32348
rect 28000 32280 28028 32320
rect 31389 32317 31401 32320
rect 31435 32317 31447 32351
rect 31389 32311 31447 32317
rect 36630 32308 36636 32360
rect 36688 32348 36694 32360
rect 39942 32348 39948 32360
rect 36688 32320 39948 32348
rect 36688 32308 36694 32320
rect 39942 32308 39948 32320
rect 40000 32308 40006 32360
rect 40034 32308 40040 32360
rect 40092 32348 40098 32360
rect 40129 32351 40187 32357
rect 40129 32348 40141 32351
rect 40092 32320 40141 32348
rect 40092 32308 40098 32320
rect 40129 32317 40141 32320
rect 40175 32317 40187 32351
rect 40402 32348 40408 32360
rect 40363 32320 40408 32348
rect 40129 32311 40187 32317
rect 40402 32308 40408 32320
rect 40460 32308 40466 32360
rect 40678 32308 40684 32360
rect 40736 32348 40742 32360
rect 53852 32348 53880 32388
rect 56597 32385 56609 32388
rect 56643 32385 56655 32419
rect 56597 32379 56655 32385
rect 55766 32348 55772 32360
rect 40736 32320 53880 32348
rect 55727 32320 55772 32348
rect 40736 32308 40742 32320
rect 55766 32308 55772 32320
rect 55824 32308 55830 32360
rect 55858 32308 55864 32360
rect 55916 32348 55922 32360
rect 55953 32351 56011 32357
rect 55953 32348 55965 32351
rect 55916 32320 55965 32348
rect 55916 32308 55922 32320
rect 55953 32317 55965 32320
rect 55999 32317 56011 32351
rect 56134 32348 56140 32360
rect 56095 32320 56140 32348
rect 55953 32311 56011 32317
rect 56134 32308 56140 32320
rect 56192 32308 56198 32360
rect 56410 32308 56416 32360
rect 56468 32348 56474 32360
rect 56505 32351 56563 32357
rect 56505 32348 56517 32351
rect 56468 32320 56517 32348
rect 56468 32308 56474 32320
rect 56505 32317 56517 32320
rect 56551 32317 56563 32351
rect 56704 32348 56732 32456
rect 56778 32444 56784 32496
rect 56836 32484 56842 32496
rect 77846 32484 77852 32496
rect 56836 32456 77852 32484
rect 56836 32444 56842 32456
rect 77846 32444 77852 32456
rect 77904 32444 77910 32496
rect 58066 32376 58072 32428
rect 58124 32416 58130 32428
rect 62850 32416 62856 32428
rect 58124 32388 62856 32416
rect 58124 32376 58130 32388
rect 62850 32376 62856 32388
rect 62908 32376 62914 32428
rect 78858 32348 78864 32360
rect 56704 32320 78864 32348
rect 56505 32311 56563 32317
rect 78858 32308 78864 32320
rect 78916 32348 78922 32360
rect 79686 32348 79692 32360
rect 78916 32320 79692 32348
rect 78916 32308 78922 32320
rect 79686 32308 79692 32320
rect 79744 32308 79750 32360
rect 84746 32308 84752 32360
rect 84804 32348 84810 32360
rect 95050 32348 95056 32360
rect 84804 32320 95056 32348
rect 84804 32308 84810 32320
rect 95050 32308 95056 32320
rect 95108 32308 95114 32360
rect 24688 32252 28028 32280
rect 28445 32283 28503 32289
rect 28445 32249 28457 32283
rect 28491 32280 28503 32283
rect 29822 32280 29828 32292
rect 28491 32252 29828 32280
rect 28491 32249 28503 32252
rect 28445 32243 28503 32249
rect 29822 32240 29828 32252
rect 29880 32240 29886 32292
rect 33686 32280 33692 32292
rect 30116 32252 33692 32280
rect 29914 32212 29920 32224
rect 22848 32184 29920 32212
rect 22695 32181 22707 32184
rect 22649 32175 22707 32181
rect 29914 32172 29920 32184
rect 29972 32212 29978 32224
rect 30116 32212 30144 32252
rect 33686 32240 33692 32252
rect 33744 32280 33750 32292
rect 41782 32280 41788 32292
rect 33744 32252 37136 32280
rect 41743 32252 41788 32280
rect 33744 32240 33750 32252
rect 29972 32184 30144 32212
rect 31389 32215 31447 32221
rect 29972 32172 29978 32184
rect 31389 32181 31401 32215
rect 31435 32212 31447 32215
rect 32493 32215 32551 32221
rect 32493 32212 32505 32215
rect 31435 32184 32505 32212
rect 31435 32181 31447 32184
rect 31389 32175 31447 32181
rect 32493 32181 32505 32184
rect 32539 32181 32551 32215
rect 32493 32175 32551 32181
rect 33870 32172 33876 32224
rect 33928 32212 33934 32224
rect 36998 32212 37004 32224
rect 33928 32184 37004 32212
rect 33928 32172 33934 32184
rect 36998 32172 37004 32184
rect 37056 32172 37062 32224
rect 37108 32212 37136 32252
rect 41782 32240 41788 32252
rect 41840 32240 41846 32292
rect 42981 32283 43039 32289
rect 42981 32249 42993 32283
rect 43027 32280 43039 32283
rect 56042 32280 56048 32292
rect 43027 32252 56048 32280
rect 43027 32249 43039 32252
rect 42981 32243 43039 32249
rect 56042 32240 56048 32252
rect 56100 32240 56106 32292
rect 59722 32280 59728 32292
rect 56888 32252 59728 32280
rect 41966 32212 41972 32224
rect 37108 32184 41972 32212
rect 41966 32172 41972 32184
rect 42024 32172 42030 32224
rect 42058 32172 42064 32224
rect 42116 32212 42122 32224
rect 46566 32212 46572 32224
rect 42116 32184 46572 32212
rect 42116 32172 42122 32184
rect 46566 32172 46572 32184
rect 46624 32172 46630 32224
rect 47026 32172 47032 32224
rect 47084 32212 47090 32224
rect 50982 32212 50988 32224
rect 47084 32184 50988 32212
rect 47084 32172 47090 32184
rect 50982 32172 50988 32184
rect 51040 32172 51046 32224
rect 51074 32172 51080 32224
rect 51132 32212 51138 32224
rect 52362 32212 52368 32224
rect 51132 32184 52368 32212
rect 51132 32172 51138 32184
rect 52362 32172 52368 32184
rect 52420 32172 52426 32224
rect 53742 32172 53748 32224
rect 53800 32212 53806 32224
rect 56888 32212 56916 32252
rect 59722 32240 59728 32252
rect 59780 32240 59786 32292
rect 68094 32240 68100 32292
rect 68152 32280 68158 32292
rect 89162 32280 89168 32292
rect 68152 32252 89168 32280
rect 68152 32240 68158 32252
rect 89162 32240 89168 32252
rect 89220 32240 89226 32292
rect 53800 32184 56916 32212
rect 56965 32215 57023 32221
rect 53800 32172 53806 32184
rect 56965 32181 56977 32215
rect 57011 32212 57023 32215
rect 87322 32212 87328 32224
rect 57011 32184 87328 32212
rect 57011 32181 57023 32184
rect 56965 32175 57023 32181
rect 87322 32172 87328 32184
rect 87380 32172 87386 32224
rect 87782 32172 87788 32224
rect 87840 32212 87846 32224
rect 95878 32212 95884 32224
rect 87840 32184 95884 32212
rect 87840 32172 87846 32184
rect 95878 32172 95884 32184
rect 95936 32172 95942 32224
rect 1104 32122 98808 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 50326 32122
rect 50378 32070 50390 32122
rect 50442 32070 50454 32122
rect 50506 32070 50518 32122
rect 50570 32070 81046 32122
rect 81098 32070 81110 32122
rect 81162 32070 81174 32122
rect 81226 32070 81238 32122
rect 81290 32070 98808 32122
rect 1104 32048 98808 32070
rect 13817 32011 13875 32017
rect 13817 31977 13829 32011
rect 13863 32008 13875 32011
rect 16022 32008 16028 32020
rect 13863 31980 16028 32008
rect 13863 31977 13875 31980
rect 13817 31971 13875 31977
rect 16022 31968 16028 31980
rect 16080 31968 16086 32020
rect 19429 32011 19487 32017
rect 16132 31980 18920 32008
rect 13722 31940 13728 31952
rect 13635 31912 13728 31940
rect 13078 31872 13084 31884
rect 13039 31844 13084 31872
rect 13078 31832 13084 31844
rect 13136 31832 13142 31884
rect 13262 31872 13268 31884
rect 13223 31844 13268 31872
rect 13262 31832 13268 31844
rect 13320 31832 13326 31884
rect 13648 31881 13676 31912
rect 13722 31900 13728 31912
rect 13780 31940 13786 31952
rect 16132 31940 16160 31980
rect 16758 31940 16764 31952
rect 13780 31912 16160 31940
rect 16719 31912 16764 31940
rect 13780 31900 13786 31912
rect 16758 31900 16764 31912
rect 16816 31900 16822 31952
rect 17034 31900 17040 31952
rect 17092 31940 17098 31952
rect 18892 31940 18920 31980
rect 19429 31977 19441 32011
rect 19475 32008 19487 32011
rect 58066 32008 58072 32020
rect 19475 31980 58072 32008
rect 19475 31977 19487 31980
rect 19429 31971 19487 31977
rect 58066 31968 58072 31980
rect 58124 31968 58130 32020
rect 58250 31968 58256 32020
rect 58308 32008 58314 32020
rect 58621 32011 58679 32017
rect 58621 32008 58633 32011
rect 58308 31980 58633 32008
rect 58308 31968 58314 31980
rect 58621 31977 58633 31980
rect 58667 31977 58679 32011
rect 58621 31971 58679 31977
rect 61010 31968 61016 32020
rect 61068 32008 61074 32020
rect 88889 32011 88947 32017
rect 88889 32008 88901 32011
rect 61068 31980 88901 32008
rect 61068 31968 61074 31980
rect 88889 31977 88901 31980
rect 88935 31977 88947 32011
rect 88889 31971 88947 31977
rect 88978 31968 88984 32020
rect 89036 32008 89042 32020
rect 89530 32008 89536 32020
rect 89036 31980 89536 32008
rect 89036 31968 89042 31980
rect 89530 31968 89536 31980
rect 89588 31968 89594 32020
rect 90358 32008 90364 32020
rect 90319 31980 90364 32008
rect 90358 31968 90364 31980
rect 90416 31968 90422 32020
rect 92566 31968 92572 32020
rect 92624 32008 92630 32020
rect 92624 31980 96660 32008
rect 92624 31968 92630 31980
rect 41414 31940 41420 31952
rect 17092 31912 18184 31940
rect 18892 31912 41420 31940
rect 17092 31900 17098 31912
rect 13633 31875 13691 31881
rect 13633 31841 13645 31875
rect 13679 31841 13691 31875
rect 15194 31872 15200 31884
rect 13633 31835 13691 31841
rect 13740 31844 15200 31872
rect 12434 31764 12440 31816
rect 12492 31804 12498 31816
rect 13357 31807 13415 31813
rect 13357 31804 13369 31807
rect 12492 31776 13369 31804
rect 12492 31764 12498 31776
rect 13357 31773 13369 31776
rect 13403 31773 13415 31807
rect 13357 31767 13415 31773
rect 13449 31807 13507 31813
rect 13449 31773 13461 31807
rect 13495 31804 13507 31807
rect 13740 31804 13768 31844
rect 15194 31832 15200 31844
rect 15252 31832 15258 31884
rect 18156 31872 18184 31912
rect 41414 31900 41420 31912
rect 41472 31900 41478 31952
rect 51074 31940 51080 31952
rect 43456 31912 51080 31940
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 18156 31844 19441 31872
rect 19429 31841 19441 31844
rect 19475 31841 19487 31875
rect 27246 31872 27252 31884
rect 19429 31835 19487 31841
rect 22066 31844 27252 31872
rect 13495 31776 13768 31804
rect 13495 31773 13507 31776
rect 13449 31767 13507 31773
rect 16850 31764 16856 31816
rect 16908 31813 16914 31816
rect 16908 31807 16966 31813
rect 16908 31773 16920 31807
rect 16954 31773 16966 31807
rect 17126 31804 17132 31816
rect 17087 31776 17132 31804
rect 16908 31767 16966 31773
rect 16908 31764 16914 31767
rect 17126 31764 17132 31776
rect 17184 31764 17190 31816
rect 19058 31764 19064 31816
rect 19116 31804 19122 31816
rect 22066 31804 22094 31844
rect 27246 31832 27252 31844
rect 27304 31832 27310 31884
rect 27706 31832 27712 31884
rect 27764 31872 27770 31884
rect 27764 31844 33640 31872
rect 27764 31832 27770 31844
rect 19116 31776 22094 31804
rect 19116 31764 19122 31776
rect 22278 31764 22284 31816
rect 22336 31804 22342 31816
rect 33505 31807 33563 31813
rect 33505 31804 33517 31807
rect 22336 31776 33517 31804
rect 22336 31764 22342 31776
rect 33505 31773 33517 31776
rect 33551 31773 33563 31807
rect 33612 31804 33640 31844
rect 33686 31832 33692 31884
rect 33744 31881 33750 31884
rect 33744 31875 33766 31881
rect 33754 31841 33766 31875
rect 33870 31872 33876 31884
rect 33831 31844 33876 31872
rect 33744 31835 33766 31841
rect 33744 31832 33750 31835
rect 33870 31832 33876 31844
rect 33928 31832 33934 31884
rect 33962 31832 33968 31884
rect 34020 31872 34026 31884
rect 41322 31872 41328 31884
rect 34020 31844 34065 31872
rect 34164 31844 41328 31872
rect 34020 31832 34026 31844
rect 34164 31804 34192 31844
rect 41322 31832 41328 31844
rect 41380 31832 41386 31884
rect 43456 31872 43484 31912
rect 51074 31900 51080 31912
rect 51132 31900 51138 31952
rect 58802 31900 58808 31952
rect 58860 31940 58866 31952
rect 84746 31940 84752 31952
rect 58860 31912 84752 31940
rect 58860 31900 58866 31912
rect 84746 31900 84752 31912
rect 84804 31900 84810 31952
rect 94685 31943 94743 31949
rect 94685 31940 94697 31943
rect 84856 31912 89944 31940
rect 41616 31844 43484 31872
rect 45005 31875 45063 31881
rect 33612 31776 34192 31804
rect 33505 31767 33563 31773
rect 37182 31764 37188 31816
rect 37240 31804 37246 31816
rect 37240 31776 38240 31804
rect 37240 31764 37246 31776
rect 17034 31736 17040 31748
rect 16995 31708 17040 31736
rect 17034 31696 17040 31708
rect 17092 31696 17098 31748
rect 17218 31736 17224 31748
rect 17179 31708 17224 31736
rect 17218 31696 17224 31708
rect 17276 31696 17282 31748
rect 17586 31696 17592 31748
rect 17644 31736 17650 31748
rect 19334 31736 19340 31748
rect 17644 31708 19340 31736
rect 17644 31696 17650 31708
rect 19334 31696 19340 31708
rect 19392 31696 19398 31748
rect 22554 31696 22560 31748
rect 22612 31736 22618 31748
rect 22612 31708 24440 31736
rect 22612 31696 22618 31708
rect 3602 31628 3608 31680
rect 3660 31668 3666 31680
rect 24026 31668 24032 31680
rect 3660 31640 24032 31668
rect 3660 31628 3666 31640
rect 24026 31628 24032 31640
rect 24084 31628 24090 31680
rect 24412 31668 24440 31708
rect 27522 31696 27528 31748
rect 27580 31736 27586 31748
rect 27580 31708 34100 31736
rect 27580 31696 27586 31708
rect 33962 31668 33968 31680
rect 24412 31640 33968 31668
rect 33962 31628 33968 31640
rect 34020 31628 34026 31680
rect 34072 31668 34100 31708
rect 36262 31696 36268 31748
rect 36320 31736 36326 31748
rect 37458 31736 37464 31748
rect 36320 31708 37464 31736
rect 36320 31696 36326 31708
rect 37458 31696 37464 31708
rect 37516 31696 37522 31748
rect 38212 31736 38240 31776
rect 38286 31764 38292 31816
rect 38344 31804 38350 31816
rect 40862 31804 40868 31816
rect 38344 31776 40868 31804
rect 38344 31764 38350 31776
rect 40862 31764 40868 31776
rect 40920 31764 40926 31816
rect 40494 31736 40500 31748
rect 38212 31708 40500 31736
rect 40494 31696 40500 31708
rect 40552 31696 40558 31748
rect 41322 31696 41328 31748
rect 41380 31736 41386 31748
rect 41616 31736 41644 31844
rect 45005 31841 45017 31875
rect 45051 31872 45063 31875
rect 45281 31875 45339 31881
rect 45281 31872 45293 31875
rect 45051 31844 45293 31872
rect 45051 31841 45063 31844
rect 45005 31835 45063 31841
rect 45281 31841 45293 31844
rect 45327 31872 45339 31875
rect 57882 31872 57888 31884
rect 45327 31844 57888 31872
rect 45327 31841 45339 31844
rect 45281 31835 45339 31841
rect 57882 31832 57888 31844
rect 57940 31832 57946 31884
rect 57974 31832 57980 31884
rect 58032 31872 58038 31884
rect 58032 31844 58076 31872
rect 58032 31832 58038 31844
rect 58158 31832 58164 31884
rect 58216 31872 58222 31884
rect 58316 31875 58374 31881
rect 58316 31872 58328 31875
rect 58216 31844 58328 31872
rect 58216 31832 58222 31844
rect 58316 31841 58328 31844
rect 58362 31841 58374 31875
rect 58316 31835 58374 31841
rect 58526 31832 58532 31884
rect 58584 31872 58590 31884
rect 66806 31872 66812 31884
rect 58584 31844 66812 31872
rect 58584 31832 58590 31844
rect 66806 31832 66812 31844
rect 66864 31832 66870 31884
rect 69658 31832 69664 31884
rect 69716 31872 69722 31884
rect 84856 31872 84884 31912
rect 89162 31872 89168 31884
rect 69716 31844 84884 31872
rect 89123 31844 89168 31872
rect 69716 31832 69722 31844
rect 89162 31832 89168 31844
rect 89220 31832 89226 31884
rect 89349 31875 89407 31881
rect 89349 31872 89361 31875
rect 89272 31844 89361 31872
rect 44174 31764 44180 31816
rect 44232 31804 44238 31816
rect 52822 31804 52828 31816
rect 44232 31776 52684 31804
rect 52783 31776 52828 31804
rect 44232 31764 44238 31776
rect 41380 31708 41644 31736
rect 41380 31696 41386 31708
rect 41782 31696 41788 31748
rect 41840 31736 41846 31748
rect 42886 31736 42892 31748
rect 41840 31708 42892 31736
rect 41840 31696 41846 31708
rect 42886 31696 42892 31708
rect 42944 31736 42950 31748
rect 44266 31736 44272 31748
rect 42944 31708 44272 31736
rect 42944 31696 42950 31708
rect 44266 31696 44272 31708
rect 44324 31696 44330 31748
rect 45830 31696 45836 31748
rect 45888 31736 45894 31748
rect 50154 31736 50160 31748
rect 45888 31708 50160 31736
rect 45888 31696 45894 31708
rect 50154 31696 50160 31708
rect 50212 31696 50218 31748
rect 38838 31668 38844 31680
rect 34072 31640 38844 31668
rect 38838 31628 38844 31640
rect 38896 31628 38902 31680
rect 39022 31628 39028 31680
rect 39080 31668 39086 31680
rect 41138 31668 41144 31680
rect 39080 31640 41144 31668
rect 39080 31628 39086 31640
rect 41138 31628 41144 31640
rect 41196 31628 41202 31680
rect 43530 31628 43536 31680
rect 43588 31668 43594 31680
rect 48406 31668 48412 31680
rect 43588 31640 48412 31668
rect 43588 31628 43594 31640
rect 48406 31628 48412 31640
rect 48464 31628 48470 31680
rect 52656 31668 52684 31776
rect 52822 31764 52828 31776
rect 52880 31764 52886 31816
rect 53101 31807 53159 31813
rect 53101 31773 53113 31807
rect 53147 31804 53159 31807
rect 53190 31804 53196 31816
rect 53147 31776 53196 31804
rect 53147 31773 53159 31776
rect 53101 31767 53159 31773
rect 53190 31764 53196 31776
rect 53248 31764 53254 31816
rect 56226 31804 56232 31816
rect 53760 31776 56232 31804
rect 53760 31668 53788 31776
rect 56226 31764 56232 31776
rect 56284 31764 56290 31816
rect 88889 31807 88947 31813
rect 58084 31776 88840 31804
rect 54202 31736 54208 31748
rect 54163 31708 54208 31736
rect 54202 31696 54208 31708
rect 54260 31696 54266 31748
rect 55030 31696 55036 31748
rect 55088 31736 55094 31748
rect 57514 31736 57520 31748
rect 55088 31708 57520 31736
rect 55088 31696 55094 31708
rect 57514 31696 57520 31708
rect 57572 31696 57578 31748
rect 58084 31736 58112 31776
rect 57992 31708 58112 31736
rect 52656 31640 53788 31668
rect 55674 31628 55680 31680
rect 55732 31668 55738 31680
rect 56134 31668 56140 31680
rect 55732 31640 56140 31668
rect 55732 31628 55738 31640
rect 56134 31628 56140 31640
rect 56192 31628 56198 31680
rect 56226 31628 56232 31680
rect 56284 31668 56290 31680
rect 57992 31668 58020 31708
rect 58342 31696 58348 31748
rect 58400 31736 58406 31748
rect 84194 31736 84200 31748
rect 58400 31708 84200 31736
rect 58400 31696 58406 31708
rect 84194 31696 84200 31708
rect 84252 31696 84258 31748
rect 56284 31640 58020 31668
rect 56284 31628 56290 31640
rect 58066 31628 58072 31680
rect 58124 31677 58130 31680
rect 58124 31671 58173 31677
rect 58124 31637 58127 31671
rect 58161 31637 58173 31671
rect 58124 31631 58173 31637
rect 58253 31671 58311 31677
rect 58253 31637 58265 31671
rect 58299 31668 58311 31671
rect 58802 31668 58808 31680
rect 58299 31640 58808 31668
rect 58299 31637 58311 31640
rect 58253 31631 58311 31637
rect 58124 31628 58130 31631
rect 58802 31628 58808 31640
rect 58860 31628 58866 31680
rect 59998 31628 60004 31680
rect 60056 31668 60062 31680
rect 60274 31668 60280 31680
rect 60056 31640 60280 31668
rect 60056 31628 60062 31640
rect 60274 31628 60280 31640
rect 60332 31628 60338 31680
rect 60550 31628 60556 31680
rect 60608 31668 60614 31680
rect 86586 31668 86592 31680
rect 60608 31640 86592 31668
rect 60608 31628 60614 31640
rect 86586 31628 86592 31640
rect 86644 31628 86650 31680
rect 88812 31668 88840 31776
rect 88889 31773 88901 31807
rect 88935 31804 88947 31807
rect 88935 31776 88969 31804
rect 88935 31773 88947 31776
rect 88889 31767 88947 31773
rect 88904 31736 88932 31767
rect 89272 31736 89300 31844
rect 89349 31841 89361 31844
rect 89395 31841 89407 31875
rect 89530 31872 89536 31884
rect 89491 31844 89536 31872
rect 89349 31835 89407 31841
rect 89530 31832 89536 31844
rect 89588 31832 89594 31884
rect 89916 31881 89944 31912
rect 90008 31912 94697 31940
rect 89901 31875 89959 31881
rect 89901 31841 89913 31875
rect 89947 31841 89959 31875
rect 89901 31835 89959 31841
rect 89806 31804 89812 31816
rect 89767 31776 89812 31804
rect 89806 31764 89812 31776
rect 89864 31764 89870 31816
rect 90008 31804 90036 31912
rect 94685 31909 94697 31912
rect 94731 31909 94743 31943
rect 94685 31903 94743 31909
rect 95712 31912 96292 31940
rect 92474 31832 92480 31884
rect 92532 31872 92538 31884
rect 95712 31872 95740 31912
rect 95878 31872 95884 31884
rect 92532 31844 95740 31872
rect 95839 31844 95884 31872
rect 92532 31832 92538 31844
rect 95878 31832 95884 31844
rect 95936 31832 95942 31884
rect 96264 31881 96292 31912
rect 96632 31881 96660 31980
rect 96249 31875 96307 31881
rect 96249 31841 96261 31875
rect 96295 31841 96307 31875
rect 96249 31835 96307 31841
rect 96617 31875 96675 31881
rect 96617 31841 96629 31875
rect 96663 31841 96675 31875
rect 96617 31835 96675 31841
rect 89916 31776 90036 31804
rect 88904 31708 89300 31736
rect 89916 31668 89944 31776
rect 90634 31764 90640 31816
rect 90692 31804 90698 31816
rect 90821 31807 90879 31813
rect 90821 31804 90833 31807
rect 90692 31776 90833 31804
rect 90692 31764 90698 31776
rect 90821 31773 90833 31776
rect 90867 31804 90879 31807
rect 91005 31807 91063 31813
rect 91005 31804 91017 31807
rect 90867 31776 91017 31804
rect 90867 31773 90879 31776
rect 90821 31767 90879 31773
rect 91005 31773 91017 31776
rect 91051 31773 91063 31807
rect 91005 31767 91063 31773
rect 94685 31807 94743 31813
rect 94685 31773 94697 31807
rect 94731 31804 94743 31807
rect 94869 31807 94927 31813
rect 94869 31804 94881 31807
rect 94731 31776 94881 31804
rect 94731 31773 94743 31776
rect 94685 31767 94743 31773
rect 94869 31773 94881 31776
rect 94915 31804 94927 31807
rect 96062 31804 96068 31816
rect 94915 31776 95924 31804
rect 96023 31776 96068 31804
rect 94915 31773 94927 31776
rect 94869 31767 94927 31773
rect 93854 31696 93860 31748
rect 93912 31736 93918 31748
rect 94961 31739 95019 31745
rect 94961 31736 94973 31739
rect 93912 31708 94973 31736
rect 93912 31696 93918 31708
rect 94961 31705 94973 31708
rect 95007 31736 95019 31739
rect 95145 31739 95203 31745
rect 95145 31736 95157 31739
rect 95007 31708 95157 31736
rect 95007 31705 95019 31708
rect 94961 31699 95019 31705
rect 95145 31705 95157 31708
rect 95191 31736 95203 31739
rect 95329 31739 95387 31745
rect 95329 31736 95341 31739
rect 95191 31708 95341 31736
rect 95191 31705 95203 31708
rect 95145 31699 95203 31705
rect 95329 31705 95341 31708
rect 95375 31736 95387 31739
rect 95513 31739 95571 31745
rect 95513 31736 95525 31739
rect 95375 31708 95525 31736
rect 95375 31705 95387 31708
rect 95329 31699 95387 31705
rect 95513 31705 95525 31708
rect 95559 31736 95571 31739
rect 95697 31739 95755 31745
rect 95697 31736 95709 31739
rect 95559 31708 95709 31736
rect 95559 31705 95571 31708
rect 95513 31699 95571 31705
rect 95697 31705 95709 31708
rect 95743 31705 95755 31739
rect 95896 31736 95924 31776
rect 96062 31764 96068 31776
rect 96120 31764 96126 31816
rect 96525 31807 96583 31813
rect 96525 31804 96537 31807
rect 96172 31776 96537 31804
rect 96172 31736 96200 31776
rect 96525 31773 96537 31776
rect 96571 31773 96583 31807
rect 96985 31807 97043 31813
rect 96985 31804 96997 31807
rect 96525 31767 96583 31773
rect 96632 31776 96997 31804
rect 96632 31736 96660 31776
rect 96985 31773 96997 31776
rect 97031 31804 97043 31807
rect 97353 31807 97411 31813
rect 97353 31804 97365 31807
rect 97031 31776 97365 31804
rect 97031 31773 97043 31776
rect 96985 31767 97043 31773
rect 97353 31773 97365 31776
rect 97399 31804 97411 31807
rect 97537 31807 97595 31813
rect 97537 31804 97549 31807
rect 97399 31776 97549 31804
rect 97399 31773 97411 31776
rect 97353 31767 97411 31773
rect 97537 31773 97549 31776
rect 97583 31804 97595 31807
rect 97721 31807 97779 31813
rect 97721 31804 97733 31807
rect 97583 31776 97733 31804
rect 97583 31773 97595 31776
rect 97537 31767 97595 31773
rect 97721 31773 97733 31776
rect 97767 31804 97779 31807
rect 97905 31807 97963 31813
rect 97905 31804 97917 31807
rect 97767 31776 97917 31804
rect 97767 31773 97779 31776
rect 97721 31767 97779 31773
rect 97905 31773 97917 31776
rect 97951 31773 97963 31807
rect 97905 31767 97963 31773
rect 95896 31708 96200 31736
rect 96540 31708 96660 31736
rect 95697 31699 95755 31705
rect 88812 31640 89944 31668
rect 95712 31668 95740 31699
rect 96540 31668 96568 31708
rect 95712 31640 96568 31668
rect 1104 31578 98808 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 65686 31578
rect 65738 31526 65750 31578
rect 65802 31526 65814 31578
rect 65866 31526 65878 31578
rect 65930 31526 96406 31578
rect 96458 31526 96470 31578
rect 96522 31526 96534 31578
rect 96586 31526 96598 31578
rect 96650 31526 98808 31578
rect 1104 31504 98808 31526
rect 3418 31424 3424 31476
rect 3476 31464 3482 31476
rect 40954 31464 40960 31476
rect 3476 31436 40960 31464
rect 3476 31424 3482 31436
rect 40954 31424 40960 31436
rect 41012 31424 41018 31476
rect 43901 31467 43959 31473
rect 43901 31433 43913 31467
rect 43947 31464 43959 31467
rect 44082 31464 44088 31476
rect 43947 31436 44088 31464
rect 43947 31433 43959 31436
rect 43901 31427 43959 31433
rect 44082 31424 44088 31436
rect 44140 31464 44146 31476
rect 44177 31467 44235 31473
rect 44177 31464 44189 31467
rect 44140 31436 44189 31464
rect 44140 31424 44146 31436
rect 44177 31433 44189 31436
rect 44223 31433 44235 31467
rect 44177 31427 44235 31433
rect 44266 31424 44272 31476
rect 44324 31464 44330 31476
rect 51810 31464 51816 31476
rect 44324 31436 51816 31464
rect 44324 31424 44330 31436
rect 51810 31424 51816 31436
rect 51868 31424 51874 31476
rect 51902 31424 51908 31476
rect 51960 31464 51966 31476
rect 51960 31436 60734 31464
rect 51960 31424 51966 31436
rect 17586 31396 17592 31408
rect 17547 31368 17592 31396
rect 17586 31356 17592 31368
rect 17644 31356 17650 31408
rect 19334 31356 19340 31408
rect 19392 31396 19398 31408
rect 19518 31396 19524 31408
rect 19392 31368 19524 31396
rect 19392 31356 19398 31368
rect 19518 31356 19524 31368
rect 19576 31356 19582 31408
rect 21266 31356 21272 31408
rect 21324 31396 21330 31408
rect 27614 31396 27620 31408
rect 21324 31368 27620 31396
rect 21324 31356 21330 31368
rect 27614 31356 27620 31368
rect 27672 31356 27678 31408
rect 27709 31399 27767 31405
rect 27709 31365 27721 31399
rect 27755 31396 27767 31399
rect 27985 31399 28043 31405
rect 27985 31396 27997 31399
rect 27755 31368 27997 31396
rect 27755 31365 27767 31368
rect 27709 31359 27767 31365
rect 27985 31365 27997 31368
rect 28031 31396 28043 31399
rect 28074 31396 28080 31408
rect 28031 31368 28080 31396
rect 28031 31365 28043 31368
rect 27985 31359 28043 31365
rect 28074 31356 28080 31368
rect 28132 31356 28138 31408
rect 28350 31356 28356 31408
rect 28408 31396 28414 31408
rect 43530 31396 43536 31408
rect 28408 31368 43536 31396
rect 28408 31356 28414 31368
rect 43530 31356 43536 31368
rect 43588 31356 43594 31408
rect 43622 31356 43628 31408
rect 43680 31396 43686 31408
rect 49326 31396 49332 31408
rect 43680 31368 49332 31396
rect 43680 31356 43686 31368
rect 49326 31356 49332 31368
rect 49384 31356 49390 31408
rect 49694 31356 49700 31408
rect 49752 31396 49758 31408
rect 52638 31396 52644 31408
rect 49752 31368 52644 31396
rect 49752 31356 49758 31368
rect 52638 31356 52644 31368
rect 52696 31356 52702 31408
rect 52822 31356 52828 31408
rect 52880 31396 52886 31408
rect 54110 31396 54116 31408
rect 52880 31368 54116 31396
rect 52880 31356 52886 31368
rect 54110 31356 54116 31368
rect 54168 31396 54174 31408
rect 54754 31396 54760 31408
rect 54168 31368 54760 31396
rect 54168 31356 54174 31368
rect 54754 31356 54760 31368
rect 54812 31356 54818 31408
rect 59633 31399 59691 31405
rect 59633 31365 59645 31399
rect 59679 31396 59691 31399
rect 60706 31396 60734 31436
rect 84194 31424 84200 31476
rect 84252 31464 84258 31476
rect 94498 31464 94504 31476
rect 84252 31436 94504 31464
rect 84252 31424 84258 31436
rect 94498 31424 94504 31436
rect 94556 31424 94562 31476
rect 94593 31399 94651 31405
rect 94593 31396 94605 31399
rect 59679 31368 60596 31396
rect 60706 31368 94605 31396
rect 59679 31365 59691 31368
rect 59633 31359 59691 31365
rect 8938 31288 8944 31340
rect 8996 31328 9002 31340
rect 18966 31328 18972 31340
rect 8996 31300 18972 31328
rect 8996 31288 9002 31300
rect 18966 31288 18972 31300
rect 19024 31288 19030 31340
rect 19061 31331 19119 31337
rect 19061 31297 19073 31331
rect 19107 31328 19119 31331
rect 19150 31328 19156 31340
rect 19107 31300 19156 31328
rect 19107 31297 19119 31300
rect 19061 31291 19119 31297
rect 19150 31288 19156 31300
rect 19208 31288 19214 31340
rect 19260 31300 19564 31328
rect 9306 31220 9312 31272
rect 9364 31260 9370 31272
rect 19260 31260 19288 31300
rect 9364 31232 19288 31260
rect 19337 31263 19395 31269
rect 9364 31220 9370 31232
rect 19337 31229 19349 31263
rect 19383 31260 19395 31263
rect 19426 31260 19432 31272
rect 19383 31232 19432 31260
rect 19383 31229 19395 31232
rect 19337 31223 19395 31229
rect 19426 31220 19432 31232
rect 19484 31220 19490 31272
rect 19536 31260 19564 31300
rect 19610 31288 19616 31340
rect 19668 31328 19674 31340
rect 59722 31328 59728 31340
rect 19668 31300 59728 31328
rect 19668 31288 19674 31300
rect 59722 31288 59728 31300
rect 59780 31288 59786 31340
rect 59909 31331 59967 31337
rect 59909 31297 59921 31331
rect 59955 31328 59967 31331
rect 60274 31328 60280 31340
rect 59955 31300 60280 31328
rect 59955 31297 59967 31300
rect 59909 31291 59967 31297
rect 54754 31260 54760 31272
rect 19536 31232 44128 31260
rect 54715 31232 54760 31260
rect 4890 31152 4896 31204
rect 4948 31192 4954 31204
rect 19518 31192 19524 31204
rect 4948 31164 17908 31192
rect 19431 31164 19524 31192
rect 4948 31152 4954 31164
rect 16850 31084 16856 31136
rect 16908 31124 16914 31136
rect 17773 31127 17831 31133
rect 17773 31124 17785 31127
rect 16908 31096 17785 31124
rect 16908 31084 16914 31096
rect 17773 31093 17785 31096
rect 17819 31093 17831 31127
rect 17880 31124 17908 31164
rect 19518 31152 19524 31164
rect 19576 31192 19582 31204
rect 20070 31192 20076 31204
rect 19576 31164 20076 31192
rect 19576 31152 19582 31164
rect 20070 31152 20076 31164
rect 20128 31152 20134 31204
rect 22066 31164 27752 31192
rect 22066 31124 22094 31164
rect 17880 31096 22094 31124
rect 17773 31087 17831 31093
rect 24302 31084 24308 31136
rect 24360 31124 24366 31136
rect 24578 31124 24584 31136
rect 24360 31096 24584 31124
rect 24360 31084 24366 31096
rect 24578 31084 24584 31096
rect 24636 31084 24642 31136
rect 26510 31084 26516 31136
rect 26568 31124 26574 31136
rect 27522 31124 27528 31136
rect 26568 31096 27528 31124
rect 26568 31084 26574 31096
rect 27522 31084 27528 31096
rect 27580 31084 27586 31136
rect 27724 31124 27752 31164
rect 28166 31152 28172 31204
rect 28224 31192 28230 31204
rect 43622 31192 43628 31204
rect 28224 31164 43628 31192
rect 28224 31152 28230 31164
rect 43622 31152 43628 31164
rect 43680 31152 43686 31204
rect 44100 31192 44128 31232
rect 54754 31220 54760 31232
rect 54812 31220 54818 31272
rect 55030 31260 55036 31272
rect 54991 31232 55036 31260
rect 55030 31220 55036 31232
rect 55088 31220 55094 31272
rect 55306 31220 55312 31272
rect 55364 31260 55370 31272
rect 59924 31260 59952 31291
rect 60274 31288 60280 31300
rect 60332 31328 60338 31340
rect 60461 31331 60519 31337
rect 60461 31328 60473 31331
rect 60332 31300 60473 31328
rect 60332 31288 60338 31300
rect 60461 31297 60473 31300
rect 60507 31297 60519 31331
rect 60461 31291 60519 31297
rect 55364 31232 59952 31260
rect 55364 31220 55370 31232
rect 59998 31220 60004 31272
rect 60056 31260 60062 31272
rect 60568 31269 60596 31368
rect 94593 31365 94605 31368
rect 94639 31365 94651 31399
rect 94593 31359 94651 31365
rect 60642 31288 60648 31340
rect 60700 31328 60706 31340
rect 93854 31328 93860 31340
rect 60700 31300 93860 31328
rect 60700 31288 60706 31300
rect 93854 31288 93860 31300
rect 93912 31288 93918 31340
rect 93946 31288 93952 31340
rect 94004 31328 94010 31340
rect 94004 31300 94176 31328
rect 94004 31288 94010 31300
rect 60185 31263 60243 31269
rect 60185 31260 60197 31263
rect 60056 31232 60197 31260
rect 60056 31220 60062 31232
rect 60185 31229 60197 31232
rect 60231 31229 60243 31263
rect 60185 31223 60243 31229
rect 60368 31263 60426 31269
rect 60368 31229 60380 31263
rect 60414 31229 60426 31263
rect 60368 31223 60426 31229
rect 60553 31263 60611 31269
rect 60553 31229 60565 31263
rect 60599 31229 60611 31263
rect 60553 31223 60611 31229
rect 43732 31164 43944 31192
rect 44100 31164 54616 31192
rect 43732 31124 43760 31164
rect 27724 31096 43760 31124
rect 43916 31124 43944 31164
rect 53742 31124 53748 31136
rect 43916 31096 53748 31124
rect 53742 31084 53748 31096
rect 53800 31084 53806 31136
rect 54588 31124 54616 31164
rect 57514 31152 57520 31204
rect 57572 31192 57578 31204
rect 59633 31195 59691 31201
rect 59633 31192 59645 31195
rect 57572 31164 59645 31192
rect 57572 31152 57578 31164
rect 59633 31161 59645 31164
rect 59679 31161 59691 31195
rect 60384 31192 60412 31223
rect 59633 31155 59691 31161
rect 60292 31164 60412 31192
rect 55306 31124 55312 31136
rect 54588 31096 55312 31124
rect 55306 31084 55312 31096
rect 55364 31084 55370 31136
rect 55674 31084 55680 31136
rect 55732 31124 55738 31136
rect 56042 31124 56048 31136
rect 55732 31096 56048 31124
rect 55732 31084 55738 31096
rect 56042 31084 56048 31096
rect 56100 31084 56106 31136
rect 56137 31127 56195 31133
rect 56137 31093 56149 31127
rect 56183 31124 56195 31127
rect 56226 31124 56232 31136
rect 56183 31096 56232 31124
rect 56183 31093 56195 31096
rect 56137 31087 56195 31093
rect 56226 31084 56232 31096
rect 56284 31084 56290 31136
rect 59998 31124 60004 31136
rect 59959 31096 60004 31124
rect 59998 31084 60004 31096
rect 60056 31084 60062 31136
rect 60182 31084 60188 31136
rect 60240 31124 60246 31136
rect 60292 31124 60320 31164
rect 60240 31096 60320 31124
rect 60568 31124 60596 31223
rect 60734 31220 60740 31272
rect 60792 31260 60798 31272
rect 60921 31263 60979 31269
rect 60792 31232 60837 31260
rect 60792 31220 60798 31232
rect 60921 31229 60933 31263
rect 60967 31260 60979 31263
rect 62022 31260 62028 31272
rect 60967 31232 62028 31260
rect 60967 31229 60979 31232
rect 60921 31223 60979 31229
rect 62022 31220 62028 31232
rect 62080 31220 62086 31272
rect 87230 31260 87236 31272
rect 87191 31232 87236 31260
rect 87230 31220 87236 31232
rect 87288 31220 87294 31272
rect 93394 31220 93400 31272
rect 93452 31260 93458 31272
rect 94041 31263 94099 31269
rect 94041 31260 94053 31263
rect 93452 31232 94053 31260
rect 93452 31220 93458 31232
rect 94041 31229 94053 31232
rect 94087 31229 94099 31263
rect 94148 31260 94176 31300
rect 94414 31263 94472 31269
rect 94414 31260 94426 31263
rect 94148 31232 94426 31260
rect 94041 31223 94099 31229
rect 94414 31229 94426 31232
rect 94460 31229 94472 31263
rect 94414 31223 94472 31229
rect 91738 31192 91744 31204
rect 86696 31164 91744 31192
rect 86696 31136 86724 31164
rect 91738 31152 91744 31164
rect 91796 31152 91802 31204
rect 91830 31152 91836 31204
rect 91888 31192 91894 31204
rect 93854 31192 93860 31204
rect 91888 31164 93860 31192
rect 91888 31152 91894 31164
rect 93854 31152 93860 31164
rect 93912 31152 93918 31204
rect 93949 31195 94007 31201
rect 93949 31161 93961 31195
rect 93995 31192 94007 31195
rect 94225 31195 94283 31201
rect 94225 31192 94237 31195
rect 93995 31164 94237 31192
rect 93995 31161 94007 31164
rect 93949 31155 94007 31161
rect 94225 31161 94237 31164
rect 94271 31161 94283 31195
rect 94225 31155 94283 31161
rect 61105 31127 61163 31133
rect 61105 31124 61117 31127
rect 60568 31096 61117 31124
rect 60240 31084 60246 31096
rect 61105 31093 61117 31096
rect 61151 31124 61163 31127
rect 86678 31124 86684 31136
rect 61151 31096 86684 31124
rect 61151 31093 61163 31096
rect 61105 31087 61163 31093
rect 86678 31084 86684 31096
rect 86736 31084 86742 31136
rect 87141 31127 87199 31133
rect 87141 31093 87153 31127
rect 87187 31124 87199 31127
rect 87230 31124 87236 31136
rect 87187 31096 87236 31124
rect 87187 31093 87199 31096
rect 87141 31087 87199 31093
rect 87230 31084 87236 31096
rect 87288 31084 87294 31136
rect 93578 31084 93584 31136
rect 93636 31124 93642 31136
rect 93964 31124 93992 31155
rect 94314 31152 94320 31204
rect 94372 31192 94378 31204
rect 94777 31195 94835 31201
rect 94777 31192 94789 31195
rect 94372 31164 94789 31192
rect 94372 31152 94378 31164
rect 94777 31161 94789 31164
rect 94823 31161 94835 31195
rect 94777 31155 94835 31161
rect 93636 31096 93992 31124
rect 93636 31084 93642 31096
rect 1104 31034 98808 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 50326 31034
rect 50378 30982 50390 31034
rect 50442 30982 50454 31034
rect 50506 30982 50518 31034
rect 50570 30982 81046 31034
rect 81098 30982 81110 31034
rect 81162 30982 81174 31034
rect 81226 30982 81238 31034
rect 81290 30982 98808 31034
rect 1104 30960 98808 30982
rect 10134 30880 10140 30932
rect 10192 30920 10198 30932
rect 57514 30920 57520 30932
rect 10192 30892 57520 30920
rect 10192 30880 10198 30892
rect 57514 30880 57520 30892
rect 57572 30880 57578 30932
rect 59354 30880 59360 30932
rect 59412 30920 59418 30932
rect 59906 30920 59912 30932
rect 59412 30892 59912 30920
rect 59412 30880 59418 30892
rect 59906 30880 59912 30892
rect 59964 30880 59970 30932
rect 60274 30880 60280 30932
rect 60332 30920 60338 30932
rect 86034 30920 86040 30932
rect 60332 30892 80054 30920
rect 85995 30892 86040 30920
rect 60332 30880 60338 30892
rect 19426 30812 19432 30864
rect 19484 30852 19490 30864
rect 20806 30852 20812 30864
rect 19484 30824 20812 30852
rect 19484 30812 19490 30824
rect 20806 30812 20812 30824
rect 20864 30812 20870 30864
rect 28350 30812 28356 30864
rect 28408 30852 28414 30864
rect 36630 30852 36636 30864
rect 28408 30824 36636 30852
rect 28408 30812 28414 30824
rect 36630 30812 36636 30824
rect 36688 30812 36694 30864
rect 36998 30812 37004 30864
rect 37056 30852 37062 30864
rect 37056 30824 60734 30852
rect 37056 30812 37062 30824
rect 11146 30744 11152 30796
rect 11204 30784 11210 30796
rect 11422 30784 11428 30796
rect 11204 30756 11428 30784
rect 11204 30744 11210 30756
rect 11422 30744 11428 30756
rect 11480 30784 11486 30796
rect 36538 30784 36544 30796
rect 11480 30756 36544 30784
rect 11480 30744 11486 30756
rect 36538 30744 36544 30756
rect 36596 30784 36602 30796
rect 37182 30784 37188 30796
rect 36596 30756 37188 30784
rect 36596 30744 36602 30756
rect 37182 30744 37188 30756
rect 37240 30744 37246 30796
rect 43625 30787 43683 30793
rect 43625 30753 43637 30787
rect 43671 30784 43683 30787
rect 43901 30787 43959 30793
rect 43901 30784 43913 30787
rect 43671 30756 43913 30784
rect 43671 30753 43683 30756
rect 43625 30747 43683 30753
rect 43901 30753 43913 30756
rect 43947 30784 43959 30787
rect 43990 30784 43996 30796
rect 43947 30756 43996 30784
rect 43947 30753 43959 30756
rect 43901 30747 43959 30753
rect 43990 30744 43996 30756
rect 44048 30744 44054 30796
rect 46014 30744 46020 30796
rect 46072 30784 46078 30796
rect 46569 30787 46627 30793
rect 46569 30784 46581 30787
rect 46072 30756 46581 30784
rect 46072 30744 46078 30756
rect 46569 30753 46581 30756
rect 46615 30753 46627 30787
rect 46569 30747 46627 30753
rect 46658 30744 46664 30796
rect 46716 30784 46722 30796
rect 46836 30787 46894 30793
rect 46836 30784 46848 30787
rect 46716 30756 46848 30784
rect 46716 30744 46722 30756
rect 46836 30753 46848 30756
rect 46882 30753 46894 30787
rect 46836 30747 46894 30753
rect 46937 30787 46995 30793
rect 46937 30753 46949 30787
rect 46983 30753 46995 30787
rect 46937 30747 46995 30753
rect 16942 30676 16948 30728
rect 17000 30716 17006 30728
rect 33870 30716 33876 30728
rect 17000 30688 33876 30716
rect 17000 30676 17006 30688
rect 33870 30676 33876 30688
rect 33928 30676 33934 30728
rect 33962 30676 33968 30728
rect 34020 30716 34026 30728
rect 35342 30716 35348 30728
rect 34020 30688 35348 30716
rect 34020 30676 34026 30688
rect 35342 30676 35348 30688
rect 35400 30676 35406 30728
rect 36722 30676 36728 30728
rect 36780 30716 36786 30728
rect 36780 30688 45968 30716
rect 36780 30676 36786 30688
rect 18506 30608 18512 30660
rect 18564 30648 18570 30660
rect 45830 30648 45836 30660
rect 18564 30620 45836 30648
rect 18564 30608 18570 30620
rect 45830 30608 45836 30620
rect 45888 30608 45894 30660
rect 45940 30648 45968 30688
rect 46290 30676 46296 30728
rect 46348 30716 46354 30728
rect 46385 30719 46443 30725
rect 46385 30716 46397 30719
rect 46348 30688 46397 30716
rect 46348 30676 46354 30688
rect 46385 30685 46397 30688
rect 46431 30685 46443 30719
rect 46750 30716 46756 30728
rect 46711 30688 46756 30716
rect 46385 30679 46443 30685
rect 46750 30676 46756 30688
rect 46808 30676 46814 30728
rect 46952 30716 46980 30747
rect 47026 30744 47032 30796
rect 47084 30784 47090 30796
rect 47121 30787 47179 30793
rect 47121 30784 47133 30787
rect 47084 30756 47133 30784
rect 47084 30744 47090 30756
rect 47121 30753 47133 30756
rect 47167 30753 47179 30787
rect 53650 30784 53656 30796
rect 47121 30747 47179 30753
rect 47504 30756 53656 30784
rect 47302 30716 47308 30728
rect 46952 30688 47308 30716
rect 47302 30676 47308 30688
rect 47360 30676 47366 30728
rect 47504 30648 47532 30756
rect 53650 30744 53656 30756
rect 53708 30744 53714 30796
rect 53742 30744 53748 30796
rect 53800 30784 53806 30796
rect 59998 30784 60004 30796
rect 53800 30756 60004 30784
rect 53800 30744 53806 30756
rect 59998 30744 60004 30756
rect 60056 30744 60062 30796
rect 60706 30784 60734 30824
rect 61102 30812 61108 30864
rect 61160 30852 61166 30864
rect 67542 30852 67548 30864
rect 61160 30824 67548 30852
rect 61160 30812 61166 30824
rect 67542 30812 67548 30824
rect 67600 30812 67606 30864
rect 72050 30812 72056 30864
rect 72108 30852 72114 30864
rect 72697 30855 72755 30861
rect 72108 30824 72556 30852
rect 72108 30812 72114 30824
rect 70670 30784 70676 30796
rect 60706 30756 70676 30784
rect 70670 30744 70676 30756
rect 70728 30784 70734 30796
rect 71682 30784 71688 30796
rect 70728 30756 71688 30784
rect 70728 30744 70734 30756
rect 71682 30744 71688 30756
rect 71740 30744 71746 30796
rect 72418 30784 72424 30796
rect 72379 30756 72424 30784
rect 72418 30744 72424 30756
rect 72476 30744 72482 30796
rect 72528 30793 72556 30824
rect 72697 30821 72709 30855
rect 72743 30852 72755 30855
rect 75454 30852 75460 30864
rect 72743 30824 75460 30852
rect 72743 30821 72755 30824
rect 72697 30815 72755 30821
rect 75454 30812 75460 30824
rect 75512 30812 75518 30864
rect 80026 30852 80054 30892
rect 86034 30880 86040 30892
rect 86092 30920 86098 30932
rect 86092 30892 86448 30920
rect 86092 30880 86098 30892
rect 86310 30852 86316 30864
rect 80026 30824 86316 30852
rect 86310 30812 86316 30824
rect 86368 30812 86374 30864
rect 86420 30861 86448 30892
rect 86405 30855 86463 30861
rect 86405 30821 86417 30855
rect 86451 30821 86463 30855
rect 86405 30815 86463 30821
rect 72514 30787 72572 30793
rect 72514 30753 72526 30787
rect 72560 30753 72572 30787
rect 72514 30747 72572 30753
rect 72786 30744 72792 30796
rect 72844 30784 72850 30796
rect 72927 30787 72985 30793
rect 72844 30756 72889 30784
rect 72844 30744 72850 30756
rect 72927 30753 72939 30787
rect 72973 30784 72985 30787
rect 73062 30784 73068 30796
rect 72973 30756 73068 30784
rect 72973 30753 72985 30756
rect 72927 30747 72985 30753
rect 73062 30744 73068 30756
rect 73120 30744 73126 30796
rect 85853 30787 85911 30793
rect 85853 30753 85865 30787
rect 85899 30784 85911 30787
rect 86221 30787 86279 30793
rect 86221 30784 86233 30787
rect 85899 30756 86233 30784
rect 85899 30753 85911 30756
rect 85853 30747 85911 30753
rect 86221 30753 86233 30756
rect 86267 30753 86279 30787
rect 86221 30747 86279 30753
rect 86497 30787 86555 30793
rect 86497 30753 86509 30787
rect 86543 30753 86555 30787
rect 86497 30747 86555 30753
rect 51074 30676 51080 30728
rect 51132 30716 51138 30728
rect 58802 30716 58808 30728
rect 51132 30688 58808 30716
rect 51132 30676 51138 30688
rect 58802 30676 58808 30688
rect 58860 30676 58866 30728
rect 59354 30716 59360 30728
rect 58912 30688 59360 30716
rect 45940 30620 47532 30648
rect 47578 30608 47584 30660
rect 47636 30648 47642 30660
rect 55214 30648 55220 30660
rect 47636 30620 55220 30648
rect 47636 30608 47642 30620
rect 55214 30608 55220 30620
rect 55272 30608 55278 30660
rect 58912 30648 58940 30688
rect 59354 30676 59360 30688
rect 59412 30676 59418 30728
rect 59630 30676 59636 30728
rect 59688 30716 59694 30728
rect 60550 30716 60556 30728
rect 59688 30688 60556 30716
rect 59688 30676 59694 30688
rect 60550 30676 60556 30688
rect 60608 30676 60614 30728
rect 63218 30676 63224 30728
rect 63276 30716 63282 30728
rect 86512 30716 86540 30747
rect 86586 30744 86592 30796
rect 86644 30793 86650 30796
rect 86644 30784 86652 30793
rect 86644 30756 86689 30784
rect 86644 30747 86652 30756
rect 86644 30744 86650 30747
rect 63276 30688 86540 30716
rect 63276 30676 63282 30688
rect 55324 30620 58940 30648
rect 13998 30540 14004 30592
rect 14056 30580 14062 30592
rect 14182 30580 14188 30592
rect 14056 30552 14188 30580
rect 14056 30540 14062 30552
rect 14182 30540 14188 30552
rect 14240 30540 14246 30592
rect 17126 30540 17132 30592
rect 17184 30580 17190 30592
rect 18782 30580 18788 30592
rect 17184 30552 18788 30580
rect 17184 30540 17190 30552
rect 18782 30540 18788 30552
rect 18840 30540 18846 30592
rect 23753 30583 23811 30589
rect 23753 30549 23765 30583
rect 23799 30580 23811 30583
rect 24029 30583 24087 30589
rect 24029 30580 24041 30583
rect 23799 30552 24041 30580
rect 23799 30549 23811 30552
rect 23753 30543 23811 30549
rect 24029 30549 24041 30552
rect 24075 30580 24087 30583
rect 45094 30580 45100 30592
rect 24075 30552 45100 30580
rect 24075 30549 24087 30552
rect 24029 30543 24087 30549
rect 45094 30540 45100 30552
rect 45152 30540 45158 30592
rect 46293 30583 46351 30589
rect 46293 30549 46305 30583
rect 46339 30580 46351 30583
rect 47026 30580 47032 30592
rect 46339 30552 47032 30580
rect 46339 30549 46351 30552
rect 46293 30543 46351 30549
rect 47026 30540 47032 30552
rect 47084 30540 47090 30592
rect 47210 30540 47216 30592
rect 47268 30580 47274 30592
rect 49142 30580 49148 30592
rect 47268 30552 49148 30580
rect 47268 30540 47274 30552
rect 49142 30540 49148 30552
rect 49200 30540 49206 30592
rect 51810 30540 51816 30592
rect 51868 30580 51874 30592
rect 55324 30580 55352 30620
rect 59078 30608 59084 30660
rect 59136 30648 59142 30660
rect 72050 30648 72056 30660
rect 59136 30620 72056 30648
rect 59136 30608 59142 30620
rect 72050 30608 72056 30620
rect 72108 30608 72114 30660
rect 85853 30651 85911 30657
rect 85853 30648 85865 30651
rect 72988 30620 85865 30648
rect 51868 30552 55352 30580
rect 51868 30540 51874 30552
rect 55490 30540 55496 30592
rect 55548 30580 55554 30592
rect 62482 30580 62488 30592
rect 55548 30552 62488 30580
rect 55548 30540 55554 30552
rect 62482 30540 62488 30552
rect 62540 30580 62546 30592
rect 63218 30580 63224 30592
rect 62540 30552 63224 30580
rect 62540 30540 62546 30552
rect 63218 30540 63224 30552
rect 63276 30540 63282 30592
rect 66898 30540 66904 30592
rect 66956 30580 66962 30592
rect 66993 30583 67051 30589
rect 66993 30580 67005 30583
rect 66956 30552 67005 30580
rect 66956 30540 66962 30552
rect 66993 30549 67005 30552
rect 67039 30580 67051 30583
rect 67177 30583 67235 30589
rect 67177 30580 67189 30583
rect 67039 30552 67189 30580
rect 67039 30549 67051 30552
rect 66993 30543 67051 30549
rect 67177 30549 67189 30552
rect 67223 30549 67235 30583
rect 67177 30543 67235 30549
rect 69474 30540 69480 30592
rect 69532 30580 69538 30592
rect 72988 30580 73016 30620
rect 85853 30617 85865 30620
rect 85899 30617 85911 30651
rect 85853 30611 85911 30617
rect 69532 30552 73016 30580
rect 73065 30583 73123 30589
rect 69532 30540 69538 30552
rect 73065 30549 73077 30583
rect 73111 30580 73123 30583
rect 74442 30580 74448 30592
rect 73111 30552 74448 30580
rect 73111 30549 73123 30552
rect 73065 30543 73123 30549
rect 74442 30540 74448 30552
rect 74500 30540 74506 30592
rect 86770 30580 86776 30592
rect 86731 30552 86776 30580
rect 86770 30540 86776 30552
rect 86828 30540 86834 30592
rect 88610 30580 88616 30592
rect 88571 30552 88616 30580
rect 88610 30540 88616 30552
rect 88668 30580 88674 30592
rect 88797 30583 88855 30589
rect 88797 30580 88809 30583
rect 88668 30552 88809 30580
rect 88668 30540 88674 30552
rect 88797 30549 88809 30552
rect 88843 30549 88855 30583
rect 88797 30543 88855 30549
rect 1104 30490 98808 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 65686 30490
rect 65738 30438 65750 30490
rect 65802 30438 65814 30490
rect 65866 30438 65878 30490
rect 65930 30438 96406 30490
rect 96458 30438 96470 30490
rect 96522 30438 96534 30490
rect 96586 30438 96598 30490
rect 96650 30438 98808 30490
rect 1104 30416 98808 30438
rect 8294 30336 8300 30388
rect 8352 30376 8358 30388
rect 9306 30376 9312 30388
rect 8352 30348 9312 30376
rect 8352 30336 8358 30348
rect 9306 30336 9312 30348
rect 9364 30336 9370 30388
rect 10318 30336 10324 30388
rect 10376 30376 10382 30388
rect 25222 30376 25228 30388
rect 10376 30348 25228 30376
rect 10376 30336 10382 30348
rect 25222 30336 25228 30348
rect 25280 30376 25286 30388
rect 30282 30376 30288 30388
rect 25280 30348 30288 30376
rect 25280 30336 25286 30348
rect 30282 30336 30288 30348
rect 30340 30336 30346 30388
rect 30374 30336 30380 30388
rect 30432 30376 30438 30388
rect 69106 30376 69112 30388
rect 30432 30348 69112 30376
rect 30432 30336 30438 30348
rect 69106 30336 69112 30348
rect 69164 30376 69170 30388
rect 70210 30376 70216 30388
rect 69164 30348 70216 30376
rect 69164 30336 69170 30348
rect 70210 30336 70216 30348
rect 70268 30336 70274 30388
rect 70949 30379 71007 30385
rect 70949 30345 70961 30379
rect 70995 30376 71007 30379
rect 71314 30376 71320 30388
rect 70995 30348 71320 30376
rect 70995 30345 71007 30348
rect 70949 30339 71007 30345
rect 71314 30336 71320 30348
rect 71372 30336 71378 30388
rect 17126 30268 17132 30320
rect 17184 30308 17190 30320
rect 54202 30308 54208 30320
rect 17184 30280 54208 30308
rect 17184 30268 17190 30280
rect 54202 30268 54208 30280
rect 54260 30268 54266 30320
rect 55122 30268 55128 30320
rect 55180 30308 55186 30320
rect 59538 30308 59544 30320
rect 55180 30280 59544 30308
rect 55180 30268 55186 30280
rect 59538 30268 59544 30280
rect 59596 30268 59602 30320
rect 60752 30280 65472 30308
rect 6086 30200 6092 30252
rect 6144 30240 6150 30252
rect 10134 30240 10140 30252
rect 6144 30212 10140 30240
rect 6144 30200 6150 30212
rect 10134 30200 10140 30212
rect 10192 30200 10198 30252
rect 10778 30200 10784 30252
rect 10836 30240 10842 30252
rect 12345 30243 12403 30249
rect 12345 30240 12357 30243
rect 10836 30212 12357 30240
rect 10836 30200 10842 30212
rect 12345 30209 12357 30212
rect 12391 30209 12403 30243
rect 12345 30203 12403 30209
rect 13998 30200 14004 30252
rect 14056 30240 14062 30252
rect 37642 30240 37648 30252
rect 14056 30212 37648 30240
rect 14056 30200 14062 30212
rect 37642 30200 37648 30212
rect 37700 30200 37706 30252
rect 43714 30200 43720 30252
rect 43772 30240 43778 30252
rect 60752 30240 60780 30280
rect 43772 30212 60780 30240
rect 65444 30240 65472 30280
rect 65610 30268 65616 30320
rect 65668 30308 65674 30320
rect 73614 30308 73620 30320
rect 65668 30280 73620 30308
rect 65668 30268 65674 30280
rect 73614 30268 73620 30280
rect 73672 30268 73678 30320
rect 71038 30240 71044 30252
rect 65444 30212 71044 30240
rect 43772 30200 43778 30212
rect 71038 30200 71044 30212
rect 71096 30200 71102 30252
rect 87877 30243 87935 30249
rect 87877 30240 87889 30243
rect 71148 30212 87889 30240
rect 9953 30175 10011 30181
rect 9953 30141 9965 30175
rect 9999 30172 10011 30175
rect 10870 30172 10876 30184
rect 9999 30144 10876 30172
rect 9999 30141 10011 30144
rect 9953 30135 10011 30141
rect 10870 30132 10876 30144
rect 10928 30132 10934 30184
rect 12066 30172 12072 30184
rect 12027 30144 12072 30172
rect 12066 30132 12072 30144
rect 12124 30132 12130 30184
rect 17218 30132 17224 30184
rect 17276 30172 17282 30184
rect 17862 30172 17868 30184
rect 17276 30144 17868 30172
rect 17276 30132 17282 30144
rect 17862 30132 17868 30144
rect 17920 30132 17926 30184
rect 24121 30175 24179 30181
rect 24121 30141 24133 30175
rect 24167 30172 24179 30175
rect 33226 30172 33232 30184
rect 24167 30144 33232 30172
rect 24167 30141 24179 30144
rect 24121 30135 24179 30141
rect 33226 30132 33232 30144
rect 33284 30172 33290 30184
rect 43625 30175 43683 30181
rect 43625 30172 43637 30175
rect 33284 30144 43637 30172
rect 33284 30132 33290 30144
rect 43625 30141 43637 30144
rect 43671 30172 43683 30175
rect 54662 30172 54668 30184
rect 43671 30144 54668 30172
rect 43671 30141 43683 30144
rect 43625 30135 43683 30141
rect 54662 30132 54668 30144
rect 54720 30132 54726 30184
rect 55122 30172 55128 30184
rect 54772 30144 55128 30172
rect 13725 30107 13783 30113
rect 13725 30073 13737 30107
rect 13771 30104 13783 30107
rect 15470 30104 15476 30116
rect 13771 30076 15476 30104
rect 13771 30073 13783 30076
rect 13725 30067 13783 30073
rect 15470 30064 15476 30076
rect 15528 30064 15534 30116
rect 24670 30104 24676 30116
rect 24631 30076 24676 30104
rect 24670 30064 24676 30076
rect 24728 30064 24734 30116
rect 25958 30064 25964 30116
rect 26016 30104 26022 30116
rect 30374 30104 30380 30116
rect 26016 30076 30380 30104
rect 26016 30064 26022 30076
rect 30374 30064 30380 30076
rect 30432 30064 30438 30116
rect 35618 30064 35624 30116
rect 35676 30104 35682 30116
rect 36354 30104 36360 30116
rect 35676 30076 36360 30104
rect 35676 30064 35682 30076
rect 36354 30064 36360 30076
rect 36412 30104 36418 30116
rect 40034 30104 40040 30116
rect 36412 30076 40040 30104
rect 36412 30064 36418 30076
rect 40034 30064 40040 30076
rect 40092 30104 40098 30116
rect 40678 30104 40684 30116
rect 40092 30076 40684 30104
rect 40092 30064 40098 30076
rect 40678 30064 40684 30076
rect 40736 30064 40742 30116
rect 42978 30064 42984 30116
rect 43036 30104 43042 30116
rect 43438 30104 43444 30116
rect 43036 30076 43444 30104
rect 43036 30064 43042 30076
rect 43438 30064 43444 30076
rect 43496 30104 43502 30116
rect 43993 30107 44051 30113
rect 43993 30104 44005 30107
rect 43496 30076 44005 30104
rect 43496 30064 43502 30076
rect 43993 30073 44005 30076
rect 44039 30073 44051 30107
rect 54772 30104 54800 30144
rect 55122 30132 55128 30144
rect 55180 30132 55186 30184
rect 55214 30132 55220 30184
rect 55272 30172 55278 30184
rect 62485 30175 62543 30181
rect 62485 30172 62497 30175
rect 55272 30144 58204 30172
rect 55272 30132 55278 30144
rect 43993 30067 44051 30073
rect 44652 30076 54800 30104
rect 12066 29996 12072 30048
rect 12124 30036 12130 30048
rect 15838 30036 15844 30048
rect 12124 30008 15844 30036
rect 12124 29996 12130 30008
rect 15838 29996 15844 30008
rect 15896 29996 15902 30048
rect 17218 29996 17224 30048
rect 17276 30036 17282 30048
rect 44652 30036 44680 30076
rect 55030 30064 55036 30116
rect 55088 30104 55094 30116
rect 58066 30104 58072 30116
rect 55088 30076 58072 30104
rect 55088 30064 55094 30076
rect 58066 30064 58072 30076
rect 58124 30064 58130 30116
rect 58176 30104 58204 30144
rect 60936 30144 62497 30172
rect 60936 30104 60964 30144
rect 62485 30141 62497 30144
rect 62531 30172 62543 30175
rect 62669 30175 62727 30181
rect 62669 30172 62681 30175
rect 62531 30144 62681 30172
rect 62531 30141 62543 30144
rect 62485 30135 62543 30141
rect 62669 30141 62681 30144
rect 62715 30141 62727 30175
rect 62669 30135 62727 30141
rect 62758 30132 62764 30184
rect 62816 30172 62822 30184
rect 68462 30172 68468 30184
rect 62816 30144 68468 30172
rect 62816 30132 62822 30144
rect 68462 30132 68468 30144
rect 68520 30132 68526 30184
rect 68554 30132 68560 30184
rect 68612 30172 68618 30184
rect 71148 30172 71176 30212
rect 87877 30209 87889 30212
rect 87923 30209 87935 30243
rect 94682 30240 94688 30252
rect 87877 30203 87935 30209
rect 91020 30212 94688 30240
rect 68612 30144 71176 30172
rect 71225 30175 71283 30181
rect 68612 30132 68618 30144
rect 71225 30141 71237 30175
rect 71271 30172 71283 30175
rect 71314 30172 71320 30184
rect 71271 30144 71320 30172
rect 71271 30141 71283 30144
rect 71225 30135 71283 30141
rect 71314 30132 71320 30144
rect 71372 30132 71378 30184
rect 80241 30175 80299 30181
rect 80241 30141 80253 30175
rect 80287 30141 80299 30175
rect 80514 30172 80520 30184
rect 80475 30144 80520 30172
rect 80241 30135 80299 30141
rect 79870 30104 79876 30116
rect 58176 30076 60964 30104
rect 61028 30076 79876 30104
rect 17276 30008 44680 30036
rect 17276 29996 17282 30008
rect 45278 29996 45284 30048
rect 45336 30036 45342 30048
rect 47210 30036 47216 30048
rect 45336 30008 47216 30036
rect 45336 29996 45342 30008
rect 47210 29996 47216 30008
rect 47268 29996 47274 30048
rect 47302 29996 47308 30048
rect 47360 30036 47366 30048
rect 48130 30036 48136 30048
rect 47360 30008 48136 30036
rect 47360 29996 47366 30008
rect 48130 29996 48136 30008
rect 48188 29996 48194 30048
rect 49326 29996 49332 30048
rect 49384 30036 49390 30048
rect 55674 30036 55680 30048
rect 49384 30008 55680 30036
rect 49384 29996 49390 30008
rect 55674 29996 55680 30008
rect 55732 29996 55738 30048
rect 59998 29996 60004 30048
rect 60056 30036 60062 30048
rect 61028 30036 61056 30076
rect 79870 30064 79876 30076
rect 79928 30064 79934 30116
rect 60056 30008 61056 30036
rect 60056 29996 60062 30008
rect 62022 29996 62028 30048
rect 62080 30036 62086 30048
rect 68278 30036 68284 30048
rect 62080 30008 68284 30036
rect 62080 29996 62086 30008
rect 68278 29996 68284 30008
rect 68336 29996 68342 30048
rect 70762 29996 70768 30048
rect 70820 30036 70826 30048
rect 73982 30036 73988 30048
rect 70820 30008 73988 30036
rect 70820 29996 70826 30008
rect 73982 29996 73988 30008
rect 74040 29996 74046 30048
rect 80256 30036 80284 30135
rect 80514 30132 80520 30144
rect 80572 30132 80578 30184
rect 86218 30132 86224 30184
rect 86276 30172 86282 30184
rect 87601 30175 87659 30181
rect 87601 30172 87613 30175
rect 86276 30144 87613 30172
rect 86276 30132 86282 30144
rect 87601 30141 87613 30144
rect 87647 30172 87659 30175
rect 89622 30172 89628 30184
rect 87647 30144 89628 30172
rect 87647 30141 87659 30144
rect 87601 30135 87659 30141
rect 89622 30132 89628 30144
rect 89680 30172 89686 30184
rect 91020 30181 91048 30212
rect 94682 30200 94688 30212
rect 94740 30240 94746 30252
rect 95142 30240 95148 30252
rect 94740 30212 95148 30240
rect 94740 30200 94746 30212
rect 95142 30200 95148 30212
rect 95200 30200 95206 30252
rect 91005 30175 91063 30181
rect 91005 30172 91017 30175
rect 89680 30144 91017 30172
rect 89680 30132 89686 30144
rect 91005 30141 91017 30144
rect 91051 30141 91063 30175
rect 91005 30135 91063 30141
rect 91281 30175 91339 30181
rect 91281 30141 91293 30175
rect 91327 30172 91339 30175
rect 93302 30172 93308 30184
rect 91327 30144 93308 30172
rect 91327 30141 91339 30144
rect 91281 30135 91339 30141
rect 93302 30132 93308 30144
rect 93360 30132 93366 30184
rect 81618 30064 81624 30116
rect 81676 30104 81682 30116
rect 81894 30104 81900 30116
rect 81676 30076 81900 30104
rect 81676 30064 81682 30076
rect 81894 30064 81900 30076
rect 81952 30064 81958 30116
rect 92658 30104 92664 30116
rect 92619 30076 92664 30104
rect 92658 30064 92664 30076
rect 92716 30064 92722 30116
rect 80882 30036 80888 30048
rect 80256 30008 80888 30036
rect 80882 29996 80888 30008
rect 80940 29996 80946 30048
rect 84470 29996 84476 30048
rect 84528 30036 84534 30048
rect 88981 30039 89039 30045
rect 88981 30036 88993 30039
rect 84528 30008 88993 30036
rect 84528 29996 84534 30008
rect 88981 30005 88993 30008
rect 89027 30005 89039 30039
rect 88981 29999 89039 30005
rect 1104 29946 98808 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 50326 29946
rect 50378 29894 50390 29946
rect 50442 29894 50454 29946
rect 50506 29894 50518 29946
rect 50570 29894 81046 29946
rect 81098 29894 81110 29946
rect 81162 29894 81174 29946
rect 81226 29894 81238 29946
rect 81290 29894 98808 29946
rect 1104 29872 98808 29894
rect 15470 29792 15476 29844
rect 15528 29832 15534 29844
rect 16390 29832 16396 29844
rect 15528 29804 16396 29832
rect 15528 29792 15534 29804
rect 16390 29792 16396 29804
rect 16448 29832 16454 29844
rect 43346 29832 43352 29844
rect 16448 29804 43352 29832
rect 16448 29792 16454 29804
rect 43346 29792 43352 29804
rect 43404 29792 43410 29844
rect 46566 29832 46572 29844
rect 46492 29804 46572 29832
rect 13446 29724 13452 29776
rect 13504 29764 13510 29776
rect 13504 29736 38240 29764
rect 13504 29724 13510 29736
rect 26142 29656 26148 29708
rect 26200 29696 26206 29708
rect 38212 29705 38240 29736
rect 38286 29724 38292 29776
rect 38344 29764 38350 29776
rect 39114 29764 39120 29776
rect 38344 29736 38424 29764
rect 39075 29736 39120 29764
rect 38344 29724 38350 29736
rect 38396 29705 38424 29736
rect 39114 29724 39120 29736
rect 39172 29764 39178 29776
rect 39172 29736 39436 29764
rect 39172 29724 39178 29736
rect 39408 29705 39436 29736
rect 43162 29724 43168 29776
rect 43220 29764 43226 29776
rect 45646 29764 45652 29776
rect 43220 29736 45652 29764
rect 43220 29724 43226 29736
rect 45646 29724 45652 29736
rect 45704 29724 45710 29776
rect 36357 29699 36415 29705
rect 36357 29696 36369 29699
rect 26200 29668 36369 29696
rect 26200 29656 26206 29668
rect 36357 29665 36369 29668
rect 36403 29665 36415 29699
rect 36357 29659 36415 29665
rect 38013 29699 38071 29705
rect 38013 29665 38025 29699
rect 38059 29665 38071 29699
rect 38013 29659 38071 29665
rect 38197 29699 38255 29705
rect 38197 29665 38209 29699
rect 38243 29665 38255 29699
rect 38197 29659 38255 29665
rect 38381 29699 38439 29705
rect 38381 29665 38393 29699
rect 38427 29665 38439 29699
rect 38381 29659 38439 29665
rect 38565 29699 38623 29705
rect 38565 29665 38577 29699
rect 38611 29665 38623 29699
rect 38565 29659 38623 29665
rect 39393 29699 39451 29705
rect 39393 29665 39405 29699
rect 39439 29665 39451 29699
rect 45738 29696 45744 29708
rect 39393 29659 39451 29665
rect 40052 29668 45744 29696
rect 20809 29631 20867 29637
rect 20809 29597 20821 29631
rect 20855 29628 20867 29631
rect 21085 29631 21143 29637
rect 21085 29628 21097 29631
rect 20855 29600 21097 29628
rect 20855 29597 20867 29600
rect 20809 29591 20867 29597
rect 21085 29597 21097 29600
rect 21131 29628 21143 29631
rect 34422 29628 34428 29640
rect 21131 29600 34428 29628
rect 21131 29597 21143 29600
rect 21085 29591 21143 29597
rect 34422 29588 34428 29600
rect 34480 29588 34486 29640
rect 35526 29588 35532 29640
rect 35584 29628 35590 29640
rect 38028 29628 38056 29659
rect 38286 29628 38292 29640
rect 35584 29600 38056 29628
rect 38247 29600 38292 29628
rect 35584 29588 35590 29600
rect 2225 29563 2283 29569
rect 2225 29529 2237 29563
rect 2271 29560 2283 29563
rect 2498 29560 2504 29572
rect 2271 29532 2504 29560
rect 2271 29529 2283 29532
rect 2225 29523 2283 29529
rect 2498 29520 2504 29532
rect 2556 29520 2562 29572
rect 6454 29520 6460 29572
rect 6512 29560 6518 29572
rect 35710 29560 35716 29572
rect 6512 29532 35716 29560
rect 6512 29520 6518 29532
rect 35710 29520 35716 29532
rect 35768 29520 35774 29572
rect 36173 29563 36231 29569
rect 36173 29529 36185 29563
rect 36219 29560 36231 29563
rect 36354 29560 36360 29572
rect 36219 29532 36360 29560
rect 36219 29529 36231 29532
rect 36173 29523 36231 29529
rect 36354 29520 36360 29532
rect 36412 29520 36418 29572
rect 15194 29452 15200 29504
rect 15252 29492 15258 29504
rect 18966 29492 18972 29504
rect 15252 29464 18972 29492
rect 15252 29452 15258 29464
rect 18966 29452 18972 29464
rect 19024 29452 19030 29504
rect 22186 29452 22192 29504
rect 22244 29492 22250 29504
rect 27706 29492 27712 29504
rect 22244 29464 27712 29492
rect 22244 29452 22250 29464
rect 27706 29452 27712 29464
rect 27764 29452 27770 29504
rect 29822 29452 29828 29504
rect 29880 29492 29886 29504
rect 30650 29492 30656 29504
rect 29880 29464 30656 29492
rect 29880 29452 29886 29464
rect 30650 29452 30656 29464
rect 30708 29452 30714 29504
rect 36909 29495 36967 29501
rect 36909 29461 36921 29495
rect 36955 29492 36967 29495
rect 37182 29492 37188 29504
rect 36955 29464 37188 29492
rect 36955 29461 36967 29464
rect 36909 29455 36967 29461
rect 37182 29452 37188 29464
rect 37240 29452 37246 29504
rect 37936 29492 37964 29600
rect 38286 29588 38292 29600
rect 38344 29588 38350 29640
rect 38580 29628 38608 29659
rect 38488 29600 38608 29628
rect 38749 29631 38807 29637
rect 38488 29572 38516 29600
rect 38749 29597 38761 29631
rect 38795 29628 38807 29631
rect 40052 29628 40080 29668
rect 45738 29656 45744 29668
rect 45796 29656 45802 29708
rect 46492 29705 46520 29804
rect 46566 29792 46572 29804
rect 46624 29792 46630 29844
rect 46934 29792 46940 29844
rect 46992 29832 46998 29844
rect 55030 29832 55036 29844
rect 46992 29804 55036 29832
rect 46992 29792 46998 29804
rect 55030 29792 55036 29804
rect 55088 29792 55094 29844
rect 55692 29804 57974 29832
rect 46658 29764 46664 29776
rect 46619 29736 46664 29764
rect 46658 29724 46664 29736
rect 46716 29724 46722 29776
rect 47210 29724 47216 29776
rect 47268 29764 47274 29776
rect 55692 29764 55720 29804
rect 47268 29736 55720 29764
rect 57946 29764 57974 29804
rect 65426 29792 65432 29844
rect 65484 29832 65490 29844
rect 65484 29804 68140 29832
rect 65484 29792 65490 29804
rect 61378 29764 61384 29776
rect 57946 29736 61384 29764
rect 47268 29724 47274 29736
rect 61378 29724 61384 29736
rect 61436 29764 61442 29776
rect 62022 29764 62028 29776
rect 61436 29736 62028 29764
rect 61436 29724 61442 29736
rect 62022 29724 62028 29736
rect 62080 29724 62086 29776
rect 68112 29764 68140 29804
rect 68278 29792 68284 29844
rect 68336 29832 68342 29844
rect 92198 29832 92204 29844
rect 68336 29804 92204 29832
rect 68336 29792 68342 29804
rect 92198 29792 92204 29804
rect 92256 29792 92262 29844
rect 70762 29764 70768 29776
rect 68112 29736 70768 29764
rect 70762 29724 70768 29736
rect 70820 29724 70826 29776
rect 88334 29764 88340 29776
rect 88295 29736 88340 29764
rect 88334 29724 88340 29736
rect 88392 29724 88398 29776
rect 46477 29699 46535 29705
rect 46477 29665 46489 29699
rect 46523 29665 46535 29699
rect 46477 29659 46535 29665
rect 46753 29699 46811 29705
rect 46753 29665 46765 29699
rect 46799 29665 46811 29699
rect 46753 29659 46811 29665
rect 38795 29600 40080 29628
rect 38795 29597 38807 29600
rect 38749 29591 38807 29597
rect 40126 29588 40132 29640
rect 40184 29628 40190 29640
rect 46198 29628 46204 29640
rect 40184 29600 46204 29628
rect 40184 29588 40190 29600
rect 46198 29588 46204 29600
rect 46256 29588 46262 29640
rect 46658 29588 46664 29640
rect 46716 29628 46722 29640
rect 46768 29628 46796 29659
rect 46934 29656 46940 29708
rect 46992 29696 46998 29708
rect 46992 29668 93854 29696
rect 46992 29656 46998 29668
rect 46716 29600 46796 29628
rect 46716 29588 46722 29600
rect 47302 29588 47308 29640
rect 47360 29628 47366 29640
rect 47360 29600 48728 29628
rect 47360 29588 47366 29600
rect 38470 29520 38476 29572
rect 38528 29520 38534 29572
rect 38562 29520 38568 29572
rect 38620 29560 38626 29572
rect 43346 29560 43352 29572
rect 38620 29532 43352 29560
rect 38620 29520 38626 29532
rect 43346 29520 43352 29532
rect 43404 29520 43410 29572
rect 45830 29520 45836 29572
rect 45888 29560 45894 29572
rect 46293 29563 46351 29569
rect 46293 29560 46305 29563
rect 45888 29532 46305 29560
rect 45888 29520 45894 29532
rect 46293 29529 46305 29532
rect 46339 29529 46351 29563
rect 48700 29560 48728 29600
rect 48774 29588 48780 29640
rect 48832 29628 48838 29640
rect 55490 29628 55496 29640
rect 48832 29600 55496 29628
rect 48832 29588 48838 29600
rect 55490 29588 55496 29600
rect 55548 29588 55554 29640
rect 55674 29588 55680 29640
rect 55732 29628 55738 29640
rect 66530 29628 66536 29640
rect 55732 29600 66536 29628
rect 55732 29588 55738 29600
rect 66530 29588 66536 29600
rect 66588 29628 66594 29640
rect 66993 29631 67051 29637
rect 66993 29628 67005 29631
rect 66588 29600 67005 29628
rect 66588 29588 66594 29600
rect 66993 29597 67005 29600
rect 67039 29597 67051 29631
rect 67174 29628 67180 29640
rect 67135 29600 67180 29628
rect 66993 29591 67051 29597
rect 67174 29588 67180 29600
rect 67232 29588 67238 29640
rect 67450 29628 67456 29640
rect 67411 29600 67456 29628
rect 67450 29588 67456 29600
rect 67508 29588 67514 29640
rect 67542 29588 67548 29640
rect 67600 29628 67606 29640
rect 68554 29628 68560 29640
rect 67600 29600 68560 29628
rect 67600 29588 67606 29600
rect 68554 29588 68560 29600
rect 68612 29588 68618 29640
rect 68646 29588 68652 29640
rect 68704 29628 68710 29640
rect 68704 29600 68876 29628
rect 68704 29588 68710 29600
rect 61010 29560 61016 29572
rect 48700 29532 61016 29560
rect 46293 29523 46351 29529
rect 61010 29520 61016 29532
rect 61068 29520 61074 29572
rect 68848 29560 68876 29600
rect 68922 29588 68928 29640
rect 68980 29628 68986 29640
rect 84470 29628 84476 29640
rect 68980 29600 84476 29628
rect 68980 29588 68986 29600
rect 84470 29588 84476 29600
rect 84528 29588 84534 29640
rect 89717 29631 89775 29637
rect 89717 29628 89729 29631
rect 88812 29600 89729 29628
rect 82906 29560 82912 29572
rect 64432 29532 67128 29560
rect 39942 29492 39948 29504
rect 37936 29464 39948 29492
rect 39942 29452 39948 29464
rect 40000 29452 40006 29504
rect 41598 29452 41604 29504
rect 41656 29492 41662 29504
rect 42610 29492 42616 29504
rect 41656 29464 42616 29492
rect 41656 29452 41662 29464
rect 42610 29452 42616 29464
rect 42668 29492 42674 29504
rect 46658 29492 46664 29504
rect 42668 29464 46664 29492
rect 42668 29452 42674 29464
rect 46658 29452 46664 29464
rect 46716 29452 46722 29504
rect 47210 29452 47216 29504
rect 47268 29492 47274 29504
rect 64432 29492 64460 29532
rect 47268 29464 64460 29492
rect 67100 29492 67128 29532
rect 68112 29532 68692 29560
rect 68848 29532 82912 29560
rect 68112 29492 68140 29532
rect 68554 29492 68560 29504
rect 67100 29464 68140 29492
rect 68515 29464 68560 29492
rect 47268 29452 47274 29464
rect 68554 29452 68560 29464
rect 68612 29452 68618 29504
rect 68664 29492 68692 29532
rect 82906 29520 82912 29532
rect 82964 29520 82970 29572
rect 84102 29520 84108 29572
rect 84160 29560 84166 29572
rect 88702 29560 88708 29572
rect 84160 29532 88708 29560
rect 84160 29520 84166 29532
rect 88702 29520 88708 29532
rect 88760 29520 88766 29572
rect 88153 29495 88211 29501
rect 88153 29492 88165 29495
rect 68664 29464 88165 29492
rect 88153 29461 88165 29464
rect 88199 29492 88211 29495
rect 88812 29492 88840 29600
rect 89717 29597 89729 29600
rect 89763 29597 89775 29631
rect 89717 29591 89775 29597
rect 89993 29631 90051 29637
rect 89993 29597 90005 29631
rect 90039 29597 90051 29631
rect 93826 29628 93854 29668
rect 94038 29628 94044 29640
rect 93826 29600 94044 29628
rect 89993 29591 90051 29597
rect 88199 29464 88840 29492
rect 88199 29461 88211 29464
rect 88153 29455 88211 29461
rect 89622 29452 89628 29504
rect 89680 29492 89686 29504
rect 90008 29492 90036 29591
rect 94038 29588 94044 29600
rect 94096 29628 94102 29640
rect 95142 29628 95148 29640
rect 94096 29600 95148 29628
rect 94096 29588 94102 29600
rect 95142 29588 95148 29600
rect 95200 29588 95206 29640
rect 89680 29464 90036 29492
rect 89680 29452 89686 29464
rect 1104 29402 98808 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 65686 29402
rect 65738 29350 65750 29402
rect 65802 29350 65814 29402
rect 65866 29350 65878 29402
rect 65930 29350 96406 29402
rect 96458 29350 96470 29402
rect 96522 29350 96534 29402
rect 96586 29350 96598 29402
rect 96650 29350 98808 29402
rect 1104 29328 98808 29350
rect 9677 29291 9735 29297
rect 9677 29257 9689 29291
rect 9723 29288 9735 29291
rect 17126 29288 17132 29300
rect 9723 29260 17132 29288
rect 9723 29257 9735 29260
rect 9677 29251 9735 29257
rect 17126 29248 17132 29260
rect 17184 29248 17190 29300
rect 17313 29291 17371 29297
rect 17313 29288 17325 29291
rect 17236 29260 17325 29288
rect 15838 29180 15844 29232
rect 15896 29220 15902 29232
rect 17236 29220 17264 29260
rect 17313 29257 17325 29260
rect 17359 29288 17371 29291
rect 19058 29288 19064 29300
rect 17359 29260 19064 29288
rect 17359 29257 17371 29260
rect 17313 29251 17371 29257
rect 19058 29248 19064 29260
rect 19116 29248 19122 29300
rect 21818 29248 21824 29300
rect 21876 29288 21882 29300
rect 68189 29291 68247 29297
rect 68189 29288 68201 29291
rect 21876 29260 68201 29288
rect 21876 29248 21882 29260
rect 68189 29257 68201 29260
rect 68235 29257 68247 29291
rect 68189 29251 68247 29257
rect 71038 29248 71044 29300
rect 71096 29288 71102 29300
rect 79689 29291 79747 29297
rect 71096 29260 76236 29288
rect 71096 29248 71102 29260
rect 26142 29220 26148 29232
rect 15896 29192 17264 29220
rect 22066 29192 26148 29220
rect 15896 29180 15902 29192
rect 8389 29155 8447 29161
rect 8389 29121 8401 29155
rect 8435 29152 8447 29155
rect 17218 29152 17224 29164
rect 8435 29124 17224 29152
rect 8435 29121 8447 29124
rect 8389 29115 8447 29121
rect 17218 29112 17224 29124
rect 17276 29112 17282 29164
rect 3510 29044 3516 29096
rect 3568 29084 3574 29096
rect 8113 29087 8171 29093
rect 8113 29084 8125 29087
rect 3568 29056 8125 29084
rect 3568 29044 3574 29056
rect 8113 29053 8125 29056
rect 8159 29084 8171 29087
rect 9398 29084 9404 29096
rect 8159 29056 9404 29084
rect 8159 29053 8171 29056
rect 8113 29047 8171 29053
rect 9398 29044 9404 29056
rect 9456 29084 9462 29096
rect 12066 29084 12072 29096
rect 9456 29056 12072 29084
rect 9456 29044 9462 29056
rect 12066 29044 12072 29056
rect 12124 29044 12130 29096
rect 13998 29084 14004 29096
rect 13959 29056 14004 29084
rect 13998 29044 14004 29056
rect 14056 29044 14062 29096
rect 15562 29084 15568 29096
rect 15523 29056 15568 29084
rect 15562 29044 15568 29056
rect 15620 29084 15626 29096
rect 15841 29087 15899 29093
rect 15841 29084 15853 29087
rect 15620 29056 15853 29084
rect 15620 29044 15626 29056
rect 15841 29053 15853 29056
rect 15887 29053 15899 29087
rect 15841 29047 15899 29053
rect 17497 29087 17555 29093
rect 17497 29053 17509 29087
rect 17543 29084 17555 29087
rect 22066 29084 22094 29192
rect 26142 29180 26148 29192
rect 26200 29180 26206 29232
rect 26326 29180 26332 29232
rect 26384 29220 26390 29232
rect 27154 29220 27160 29232
rect 26384 29192 27160 29220
rect 26384 29180 26390 29192
rect 27154 29180 27160 29192
rect 27212 29180 27218 29232
rect 36998 29220 37004 29232
rect 36959 29192 37004 29220
rect 36998 29180 37004 29192
rect 37056 29180 37062 29232
rect 37182 29180 37188 29232
rect 37240 29220 37246 29232
rect 42058 29220 42064 29232
rect 37240 29192 42064 29220
rect 37240 29180 37246 29192
rect 42058 29180 42064 29192
rect 42116 29180 42122 29232
rect 42153 29223 42211 29229
rect 42153 29189 42165 29223
rect 42199 29220 42211 29223
rect 42429 29223 42487 29229
rect 42429 29220 42441 29223
rect 42199 29192 42441 29220
rect 42199 29189 42211 29192
rect 42153 29183 42211 29189
rect 42429 29189 42441 29192
rect 42475 29220 42487 29223
rect 42794 29220 42800 29232
rect 42475 29192 42800 29220
rect 42475 29189 42487 29192
rect 42429 29183 42487 29189
rect 42794 29180 42800 29192
rect 42852 29180 42858 29232
rect 46198 29180 46204 29232
rect 46256 29220 46262 29232
rect 46934 29220 46940 29232
rect 46256 29192 46940 29220
rect 46256 29180 46262 29192
rect 46934 29180 46940 29192
rect 46992 29180 46998 29232
rect 53742 29180 53748 29232
rect 53800 29220 53806 29232
rect 56502 29220 56508 29232
rect 53800 29192 56508 29220
rect 53800 29180 53806 29192
rect 56502 29180 56508 29192
rect 56560 29180 56566 29232
rect 57146 29180 57152 29232
rect 57204 29220 57210 29232
rect 57330 29220 57336 29232
rect 57204 29192 57336 29220
rect 57204 29180 57210 29192
rect 57330 29180 57336 29192
rect 57388 29180 57394 29232
rect 57514 29180 57520 29232
rect 57572 29220 57578 29232
rect 65426 29220 65432 29232
rect 57572 29192 65432 29220
rect 57572 29180 57578 29192
rect 65426 29180 65432 29192
rect 65484 29180 65490 29232
rect 67818 29180 67824 29232
rect 67876 29220 67882 29232
rect 67913 29223 67971 29229
rect 67913 29220 67925 29223
rect 67876 29192 67925 29220
rect 67876 29180 67882 29192
rect 67913 29189 67925 29192
rect 67959 29220 67971 29223
rect 68646 29220 68652 29232
rect 67959 29192 68652 29220
rect 67959 29189 67971 29192
rect 67913 29183 67971 29189
rect 68646 29180 68652 29192
rect 68704 29180 68710 29232
rect 68830 29180 68836 29232
rect 68888 29220 68894 29232
rect 75917 29223 75975 29229
rect 75917 29220 75929 29223
rect 68888 29192 75929 29220
rect 68888 29180 68894 29192
rect 75917 29189 75929 29192
rect 75963 29220 75975 29223
rect 76101 29223 76159 29229
rect 76101 29220 76113 29223
rect 75963 29192 76113 29220
rect 75963 29189 75975 29192
rect 75917 29183 75975 29189
rect 76101 29189 76113 29192
rect 76147 29189 76159 29223
rect 76208 29220 76236 29260
rect 79689 29257 79701 29291
rect 79735 29288 79747 29291
rect 79735 29260 93854 29288
rect 79735 29257 79747 29260
rect 79689 29251 79747 29257
rect 83918 29220 83924 29232
rect 76208 29192 83924 29220
rect 76101 29183 76159 29189
rect 83918 29180 83924 29192
rect 83976 29220 83982 29232
rect 84102 29220 84108 29232
rect 83976 29192 84108 29220
rect 83976 29180 83982 29192
rect 84102 29180 84108 29192
rect 84160 29180 84166 29232
rect 86218 29180 86224 29232
rect 86276 29220 86282 29232
rect 93826 29220 93854 29260
rect 95878 29248 95884 29300
rect 95936 29288 95942 29300
rect 95936 29260 97304 29288
rect 95936 29248 95942 29260
rect 86276 29192 87092 29220
rect 93826 29192 97212 29220
rect 86276 29180 86282 29192
rect 24302 29112 24308 29164
rect 24360 29152 24366 29164
rect 24762 29152 24768 29164
rect 24360 29124 24768 29152
rect 24360 29112 24366 29124
rect 24762 29112 24768 29124
rect 24820 29152 24826 29164
rect 68557 29155 68615 29161
rect 24820 29124 35756 29152
rect 24820 29112 24826 29124
rect 17543 29056 22094 29084
rect 23937 29087 23995 29093
rect 17543 29053 17555 29056
rect 17497 29047 17555 29053
rect 23937 29053 23949 29087
rect 23983 29084 23995 29087
rect 24210 29084 24216 29096
rect 23983 29056 24216 29084
rect 23983 29053 23995 29056
rect 23937 29047 23995 29053
rect 24210 29044 24216 29056
rect 24268 29044 24274 29096
rect 26329 29087 26387 29093
rect 26329 29053 26341 29087
rect 26375 29084 26387 29087
rect 26602 29084 26608 29096
rect 26375 29056 26608 29084
rect 26375 29053 26387 29056
rect 26329 29047 26387 29053
rect 26602 29044 26608 29056
rect 26660 29044 26666 29096
rect 33410 29044 33416 29096
rect 33468 29084 33474 29096
rect 35618 29084 35624 29096
rect 33468 29056 35624 29084
rect 33468 29044 33474 29056
rect 35618 29044 35624 29056
rect 35676 29044 35682 29096
rect 35728 29084 35756 29124
rect 36648 29124 68140 29152
rect 36648 29084 36676 29124
rect 35728 29056 36676 29084
rect 38102 29044 38108 29096
rect 38160 29084 38166 29096
rect 38286 29084 38292 29096
rect 38160 29056 38292 29084
rect 38160 29044 38166 29056
rect 38286 29044 38292 29056
rect 38344 29044 38350 29096
rect 38470 29044 38476 29096
rect 38528 29084 38534 29096
rect 38528 29056 45692 29084
rect 38528 29044 38534 29056
rect 14550 29016 14556 29028
rect 14511 28988 14556 29016
rect 14550 28976 14556 28988
rect 14608 28976 14614 29028
rect 35888 29019 35946 29025
rect 23768 28988 23980 29016
rect 9030 28908 9036 28960
rect 9088 28948 9094 28960
rect 23768 28948 23796 28988
rect 9088 28920 23796 28948
rect 23952 28948 23980 28988
rect 26068 28988 26280 29016
rect 26068 28948 26096 28988
rect 23952 28920 26096 28948
rect 26252 28948 26280 28988
rect 35888 28985 35900 29019
rect 35934 29016 35946 29019
rect 36722 29016 36728 29028
rect 35934 28988 36728 29016
rect 35934 28985 35946 28988
rect 35888 28979 35946 28985
rect 36722 28976 36728 28988
rect 36780 28976 36786 29028
rect 45664 29016 45692 29056
rect 45830 29044 45836 29096
rect 45888 29084 45894 29096
rect 68112 29084 68140 29124
rect 68557 29121 68569 29155
rect 68603 29152 68615 29155
rect 79042 29152 79048 29164
rect 68603 29124 79048 29152
rect 68603 29121 68615 29124
rect 68557 29115 68615 29121
rect 79042 29112 79048 29124
rect 79100 29112 79106 29164
rect 86954 29152 86960 29164
rect 86915 29124 86960 29152
rect 86954 29112 86960 29124
rect 87012 29112 87018 29164
rect 87064 29152 87092 29192
rect 88521 29155 88579 29161
rect 88521 29152 88533 29155
rect 87064 29124 88533 29152
rect 88521 29121 88533 29124
rect 88567 29121 88579 29155
rect 88521 29115 88579 29121
rect 88702 29112 88708 29164
rect 88760 29152 88766 29164
rect 97184 29161 97212 29192
rect 96893 29155 96951 29161
rect 96893 29152 96905 29155
rect 88760 29124 96905 29152
rect 88760 29112 88766 29124
rect 96893 29121 96905 29124
rect 96939 29121 96951 29155
rect 96893 29115 96951 29121
rect 97169 29155 97227 29161
rect 97169 29121 97181 29155
rect 97215 29121 97227 29155
rect 97169 29115 97227 29121
rect 68281 29087 68339 29093
rect 68281 29084 68293 29087
rect 45888 29056 68048 29084
rect 68112 29056 68293 29084
rect 45888 29044 45894 29056
rect 46106 29016 46112 29028
rect 36924 28988 37136 29016
rect 36924 28948 36952 28988
rect 26252 28920 36952 28948
rect 37108 28948 37136 28988
rect 41984 28988 42196 29016
rect 45664 28988 46112 29016
rect 41984 28948 42012 28988
rect 37108 28920 42012 28948
rect 42168 28948 42196 28988
rect 46106 28976 46112 28988
rect 46164 28976 46170 29028
rect 46198 28976 46204 29028
rect 46256 29016 46262 29028
rect 55306 29016 55312 29028
rect 46256 28988 55312 29016
rect 46256 28976 46262 28988
rect 55306 28976 55312 28988
rect 55364 28976 55370 29028
rect 55490 28976 55496 29028
rect 55548 29016 55554 29028
rect 67910 29016 67916 29028
rect 55548 28988 67916 29016
rect 55548 28976 55554 28988
rect 67910 28976 67916 28988
rect 67968 28976 67974 29028
rect 53834 28948 53840 28960
rect 42168 28920 53840 28948
rect 9088 28908 9094 28920
rect 53834 28908 53840 28920
rect 53892 28908 53898 28960
rect 55674 28908 55680 28960
rect 55732 28948 55738 28960
rect 59630 28948 59636 28960
rect 55732 28920 59636 28948
rect 55732 28908 55738 28920
rect 59630 28908 59636 28920
rect 59688 28908 59694 28960
rect 59722 28908 59728 28960
rect 59780 28948 59786 28960
rect 63034 28948 63040 28960
rect 59780 28920 63040 28948
rect 59780 28908 59786 28920
rect 63034 28908 63040 28920
rect 63092 28908 63098 28960
rect 63126 28908 63132 28960
rect 63184 28948 63190 28960
rect 67174 28948 67180 28960
rect 63184 28920 67180 28948
rect 63184 28908 63190 28920
rect 67174 28908 67180 28920
rect 67232 28908 67238 28960
rect 68020 28948 68048 29056
rect 68281 29053 68293 29056
rect 68327 29053 68339 29087
rect 68462 29084 68468 29096
rect 68423 29056 68468 29084
rect 68281 29047 68339 29053
rect 68462 29044 68468 29056
rect 68520 29044 68526 29096
rect 68646 29044 68652 29096
rect 68704 29084 68710 29096
rect 68833 29087 68891 29093
rect 68704 29056 68749 29084
rect 68704 29044 68710 29056
rect 68833 29053 68845 29087
rect 68879 29084 68891 29087
rect 68922 29084 68928 29096
rect 68879 29056 68928 29084
rect 68879 29053 68891 29056
rect 68833 29047 68891 29053
rect 68922 29044 68928 29056
rect 68980 29044 68986 29096
rect 71130 29044 71136 29096
rect 71188 29084 71194 29096
rect 71225 29087 71283 29093
rect 71225 29084 71237 29087
rect 71188 29056 71237 29084
rect 71188 29044 71194 29056
rect 71225 29053 71237 29056
rect 71271 29053 71283 29087
rect 71225 29047 71283 29053
rect 73982 29044 73988 29096
rect 74040 29084 74046 29096
rect 79689 29087 79747 29093
rect 79689 29084 79701 29087
rect 74040 29056 79701 29084
rect 74040 29044 74046 29056
rect 79689 29053 79701 29056
rect 79735 29053 79747 29087
rect 79689 29047 79747 29053
rect 86586 29044 86592 29096
rect 86644 29084 86650 29096
rect 86681 29087 86739 29093
rect 86681 29084 86693 29087
rect 86644 29056 86693 29084
rect 86644 29044 86650 29056
rect 86681 29053 86693 29056
rect 86727 29084 86739 29087
rect 88245 29087 88303 29093
rect 88245 29084 88257 29087
rect 86727 29056 88257 29084
rect 86727 29053 86739 29056
rect 86681 29047 86739 29053
rect 88245 29053 88257 29056
rect 88291 29053 88303 29087
rect 88245 29047 88303 29053
rect 69382 28976 69388 29028
rect 69440 29016 69446 29028
rect 79594 29016 79600 29028
rect 69440 28988 79600 29016
rect 69440 28976 69446 28988
rect 79594 28976 79600 28988
rect 79652 28976 79658 29028
rect 96908 29016 96936 29115
rect 97276 29093 97304 29260
rect 97261 29087 97319 29093
rect 97261 29053 97273 29087
rect 97307 29053 97319 29087
rect 97261 29047 97319 29053
rect 97629 29087 97687 29093
rect 97629 29053 97641 29087
rect 97675 29053 97687 29087
rect 97629 29047 97687 29053
rect 97644 29016 97672 29047
rect 98086 29016 98092 29028
rect 86604 28988 86816 29016
rect 96908 28988 97672 29016
rect 98047 28988 98092 29016
rect 68278 28948 68284 28960
rect 68020 28920 68284 28948
rect 68278 28908 68284 28920
rect 68336 28908 68342 28960
rect 71038 28948 71044 28960
rect 70999 28920 71044 28948
rect 71038 28908 71044 28920
rect 71096 28908 71102 28960
rect 74718 28908 74724 28960
rect 74776 28948 74782 28960
rect 86604 28948 86632 28988
rect 74776 28920 86632 28948
rect 86788 28948 86816 28988
rect 98086 28976 98092 28988
rect 98144 28976 98150 29028
rect 92658 28948 92664 28960
rect 86788 28920 92664 28948
rect 74776 28908 74782 28920
rect 92658 28908 92664 28920
rect 92716 28908 92722 28960
rect 1104 28858 98808 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 50326 28858
rect 50378 28806 50390 28858
rect 50442 28806 50454 28858
rect 50506 28806 50518 28858
rect 50570 28806 81046 28858
rect 81098 28806 81110 28858
rect 81162 28806 81174 28858
rect 81226 28806 81238 28858
rect 81290 28806 98808 28858
rect 1104 28784 98808 28806
rect 4062 28704 4068 28756
rect 4120 28744 4126 28756
rect 22554 28744 22560 28756
rect 4120 28716 22560 28744
rect 4120 28704 4126 28716
rect 22554 28704 22560 28716
rect 22612 28704 22618 28756
rect 26786 28704 26792 28756
rect 26844 28744 26850 28756
rect 26844 28716 26924 28744
rect 26844 28704 26850 28716
rect 26896 28676 26924 28716
rect 28074 28704 28080 28756
rect 28132 28744 28138 28756
rect 37001 28747 37059 28753
rect 28132 28716 35848 28744
rect 28132 28704 28138 28716
rect 33229 28679 33287 28685
rect 9646 28648 15792 28676
rect 1673 28611 1731 28617
rect 1673 28577 1685 28611
rect 1719 28608 1731 28611
rect 3510 28608 3516 28620
rect 1719 28580 3516 28608
rect 1719 28577 1731 28580
rect 1673 28571 1731 28577
rect 3510 28568 3516 28580
rect 3568 28568 3574 28620
rect 6730 28568 6736 28620
rect 6788 28608 6794 28620
rect 9646 28608 9674 28648
rect 15654 28608 15660 28620
rect 6788 28580 9674 28608
rect 15615 28580 15660 28608
rect 6788 28568 6794 28580
rect 15654 28568 15660 28580
rect 15712 28568 15718 28620
rect 15764 28608 15792 28648
rect 16592 28648 26372 28676
rect 26896 28648 31754 28676
rect 16592 28608 16620 28648
rect 15764 28580 16620 28608
rect 17034 28568 17040 28620
rect 17092 28608 17098 28620
rect 20530 28608 20536 28620
rect 17092 28580 20536 28608
rect 17092 28568 17098 28580
rect 20530 28568 20536 28580
rect 20588 28568 20594 28620
rect 20806 28608 20812 28620
rect 20767 28580 20812 28608
rect 20806 28568 20812 28580
rect 20864 28568 20870 28620
rect 20916 28580 21220 28608
rect 1949 28543 2007 28549
rect 1949 28509 1961 28543
rect 1995 28540 2007 28543
rect 15197 28543 15255 28549
rect 1995 28512 12434 28540
rect 1995 28509 2007 28512
rect 1949 28503 2007 28509
rect 3237 28407 3295 28413
rect 3237 28373 3249 28407
rect 3283 28404 3295 28407
rect 5350 28404 5356 28416
rect 3283 28376 5356 28404
rect 3283 28373 3295 28376
rect 3237 28367 3295 28373
rect 5350 28364 5356 28376
rect 5408 28364 5414 28416
rect 5445 28407 5503 28413
rect 5445 28373 5457 28407
rect 5491 28404 5503 28407
rect 5721 28407 5779 28413
rect 5721 28404 5733 28407
rect 5491 28376 5733 28404
rect 5491 28373 5503 28376
rect 5445 28367 5503 28373
rect 5721 28373 5733 28376
rect 5767 28404 5779 28407
rect 5994 28404 6000 28416
rect 5767 28376 6000 28404
rect 5767 28373 5779 28376
rect 5721 28367 5779 28373
rect 5994 28364 6000 28376
rect 6052 28364 6058 28416
rect 12406 28404 12434 28512
rect 15197 28509 15209 28543
rect 15243 28540 15255 28543
rect 15381 28543 15439 28549
rect 15381 28540 15393 28543
rect 15243 28512 15393 28540
rect 15243 28509 15255 28512
rect 15197 28503 15255 28509
rect 15381 28509 15393 28512
rect 15427 28540 15439 28543
rect 15565 28543 15623 28549
rect 15565 28540 15577 28543
rect 15427 28512 15577 28540
rect 15427 28509 15439 28512
rect 15381 28503 15439 28509
rect 15565 28509 15577 28512
rect 15611 28540 15623 28543
rect 15933 28543 15991 28549
rect 15933 28540 15945 28543
rect 15611 28512 15945 28540
rect 15611 28509 15623 28512
rect 15565 28503 15623 28509
rect 15933 28509 15945 28512
rect 15979 28540 15991 28543
rect 16574 28540 16580 28552
rect 15979 28512 16580 28540
rect 15979 28509 15991 28512
rect 15933 28503 15991 28509
rect 16574 28500 16580 28512
rect 16632 28500 16638 28552
rect 16758 28500 16764 28552
rect 16816 28540 16822 28552
rect 20916 28540 20944 28580
rect 16816 28512 20944 28540
rect 16816 28500 16822 28512
rect 20990 28500 20996 28552
rect 21048 28540 21054 28552
rect 21085 28543 21143 28549
rect 21085 28540 21097 28543
rect 21048 28512 21097 28540
rect 21048 28500 21054 28512
rect 21085 28509 21097 28512
rect 21131 28509 21143 28543
rect 21192 28540 21220 28580
rect 26234 28540 26240 28552
rect 21192 28512 26240 28540
rect 21085 28503 21143 28509
rect 26234 28500 26240 28512
rect 26292 28500 26298 28552
rect 14274 28432 14280 28484
rect 14332 28472 14338 28484
rect 22094 28472 22100 28484
rect 14332 28444 15608 28472
rect 14332 28432 14338 28444
rect 15102 28404 15108 28416
rect 12406 28376 15108 28404
rect 15102 28364 15108 28376
rect 15160 28364 15166 28416
rect 15580 28404 15608 28444
rect 16592 28444 22100 28472
rect 16592 28404 16620 28444
rect 22094 28432 22100 28444
rect 22152 28472 22158 28484
rect 23382 28472 23388 28484
rect 22152 28444 23388 28472
rect 22152 28432 22158 28444
rect 23382 28432 23388 28444
rect 23440 28432 23446 28484
rect 26344 28472 26372 28648
rect 31726 28608 31754 28648
rect 33229 28645 33241 28679
rect 33275 28676 33287 28679
rect 33597 28679 33655 28685
rect 33597 28676 33609 28679
rect 33275 28648 33609 28676
rect 33275 28645 33287 28648
rect 33229 28639 33287 28645
rect 33597 28645 33609 28648
rect 33643 28676 33655 28679
rect 35820 28676 35848 28716
rect 37001 28713 37013 28747
rect 37047 28744 37059 28747
rect 37366 28744 37372 28756
rect 37047 28716 37372 28744
rect 37047 28713 37059 28716
rect 37001 28707 37059 28713
rect 37366 28704 37372 28716
rect 37424 28704 37430 28756
rect 46198 28744 46204 28756
rect 37476 28716 46204 28744
rect 37476 28676 37504 28716
rect 46198 28704 46204 28716
rect 46256 28704 46262 28756
rect 47026 28704 47032 28756
rect 47084 28744 47090 28756
rect 47084 28716 52316 28744
rect 47084 28704 47090 28716
rect 37734 28676 37740 28688
rect 33643 28648 35756 28676
rect 35820 28648 37504 28676
rect 37695 28648 37740 28676
rect 33643 28645 33655 28648
rect 33597 28639 33655 28645
rect 33321 28611 33379 28617
rect 33321 28608 33333 28611
rect 31726 28580 33333 28608
rect 33321 28577 33333 28580
rect 33367 28577 33379 28611
rect 33502 28608 33508 28620
rect 33463 28580 33508 28608
rect 33321 28571 33379 28577
rect 33502 28568 33508 28580
rect 33560 28568 33566 28620
rect 33689 28611 33747 28617
rect 33689 28577 33701 28611
rect 33735 28577 33747 28611
rect 35728 28608 35756 28648
rect 37734 28636 37740 28648
rect 37792 28636 37798 28688
rect 39666 28636 39672 28688
rect 39724 28676 39730 28688
rect 48038 28676 48044 28688
rect 39724 28648 48044 28676
rect 39724 28636 39730 28648
rect 48038 28636 48044 28648
rect 48096 28636 48102 28688
rect 52288 28676 52316 28716
rect 52362 28704 52368 28756
rect 52420 28744 52426 28756
rect 97902 28744 97908 28756
rect 52420 28716 97908 28744
rect 52420 28704 52426 28716
rect 97902 28704 97908 28716
rect 97960 28704 97966 28756
rect 52288 28648 55812 28676
rect 36998 28608 37004 28620
rect 35728 28580 37004 28608
rect 33689 28571 33747 28577
rect 27154 28500 27160 28552
rect 27212 28540 27218 28552
rect 33704 28540 33732 28571
rect 36998 28568 37004 28580
rect 37056 28568 37062 28620
rect 37274 28608 37280 28620
rect 37235 28580 37280 28608
rect 37274 28568 37280 28580
rect 37332 28568 37338 28620
rect 37550 28608 37556 28620
rect 37511 28580 37556 28608
rect 37550 28568 37556 28580
rect 37608 28568 37614 28620
rect 55674 28608 55680 28620
rect 37660 28580 55680 28608
rect 37660 28540 37688 28580
rect 55674 28568 55680 28580
rect 55732 28568 55738 28620
rect 27212 28512 37688 28540
rect 27212 28500 27218 28512
rect 37734 28500 37740 28552
rect 37792 28540 37798 28552
rect 42426 28540 42432 28552
rect 37792 28512 42432 28540
rect 37792 28500 37798 28512
rect 42426 28500 42432 28512
rect 42484 28500 42490 28552
rect 42518 28500 42524 28552
rect 42576 28540 42582 28552
rect 46290 28540 46296 28552
rect 42576 28512 46296 28540
rect 42576 28500 42582 28512
rect 46290 28500 46296 28512
rect 46348 28500 46354 28552
rect 49145 28543 49203 28549
rect 49145 28540 49157 28543
rect 47964 28512 49157 28540
rect 31754 28472 31760 28484
rect 26344 28444 31760 28472
rect 31754 28432 31760 28444
rect 31812 28432 31818 28484
rect 47857 28475 47915 28481
rect 47857 28472 47869 28475
rect 31864 28444 47869 28472
rect 17218 28404 17224 28416
rect 15580 28376 16620 28404
rect 17179 28376 17224 28404
rect 17218 28364 17224 28376
rect 17276 28364 17282 28416
rect 17497 28407 17555 28413
rect 17497 28373 17509 28407
rect 17543 28404 17555 28407
rect 17681 28407 17739 28413
rect 17681 28404 17693 28407
rect 17543 28376 17693 28404
rect 17543 28373 17555 28376
rect 17497 28367 17555 28373
rect 17681 28373 17693 28376
rect 17727 28404 17739 28407
rect 17770 28404 17776 28416
rect 17727 28376 17776 28404
rect 17727 28373 17739 28376
rect 17681 28367 17739 28373
rect 17770 28364 17776 28376
rect 17828 28364 17834 28416
rect 18782 28364 18788 28416
rect 18840 28404 18846 28416
rect 19242 28404 19248 28416
rect 18840 28376 19248 28404
rect 18840 28364 18846 28376
rect 19242 28364 19248 28376
rect 19300 28364 19306 28416
rect 19886 28364 19892 28416
rect 19944 28404 19950 28416
rect 20162 28404 20168 28416
rect 19944 28376 20168 28404
rect 19944 28364 19950 28376
rect 20162 28364 20168 28376
rect 20220 28364 20226 28416
rect 20530 28364 20536 28416
rect 20588 28404 20594 28416
rect 27154 28404 27160 28416
rect 20588 28376 27160 28404
rect 20588 28364 20594 28376
rect 27154 28364 27160 28376
rect 27212 28364 27218 28416
rect 30282 28364 30288 28416
rect 30340 28404 30346 28416
rect 31864 28404 31892 28444
rect 47857 28441 47869 28444
rect 47903 28441 47915 28475
rect 47857 28435 47915 28441
rect 33870 28404 33876 28416
rect 30340 28376 31892 28404
rect 33831 28376 33876 28404
rect 30340 28364 30346 28376
rect 33870 28364 33876 28376
rect 33928 28364 33934 28416
rect 36998 28404 37004 28416
rect 36911 28376 37004 28404
rect 36998 28364 37004 28376
rect 37056 28404 37062 28416
rect 37093 28407 37151 28413
rect 37093 28404 37105 28407
rect 37056 28376 37105 28404
rect 37056 28364 37062 28376
rect 37093 28373 37105 28376
rect 37139 28373 37151 28407
rect 37093 28367 37151 28373
rect 38286 28364 38292 28416
rect 38344 28404 38350 28416
rect 47581 28407 47639 28413
rect 47581 28404 47593 28407
rect 38344 28376 47593 28404
rect 38344 28364 38350 28376
rect 47581 28373 47593 28376
rect 47627 28404 47639 28407
rect 47964 28404 47992 28512
rect 49145 28509 49157 28512
rect 49191 28509 49203 28543
rect 49418 28540 49424 28552
rect 49379 28512 49424 28540
rect 49145 28503 49203 28509
rect 49418 28500 49424 28512
rect 49476 28500 49482 28552
rect 49786 28500 49792 28552
rect 49844 28540 49850 28552
rect 52454 28540 52460 28552
rect 49844 28512 52460 28540
rect 49844 28500 49850 28512
rect 52454 28500 52460 28512
rect 52512 28500 52518 28552
rect 53650 28500 53656 28552
rect 53708 28540 53714 28552
rect 53834 28540 53840 28552
rect 53708 28512 53840 28540
rect 53708 28500 53714 28512
rect 53834 28500 53840 28512
rect 53892 28500 53898 28552
rect 55784 28540 55812 28648
rect 60366 28636 60372 28688
rect 60424 28676 60430 28688
rect 71038 28676 71044 28688
rect 60424 28648 62068 28676
rect 60424 28636 60430 28648
rect 56318 28568 56324 28620
rect 56376 28608 56382 28620
rect 61930 28608 61936 28620
rect 56376 28580 61936 28608
rect 56376 28568 56382 28580
rect 61930 28568 61936 28580
rect 61988 28568 61994 28620
rect 61838 28540 61844 28552
rect 55784 28512 61844 28540
rect 61838 28500 61844 28512
rect 61896 28500 61902 28552
rect 62040 28540 62068 28648
rect 62132 28648 71044 28676
rect 62132 28617 62160 28648
rect 71038 28636 71044 28648
rect 71096 28676 71102 28688
rect 71096 28648 80054 28676
rect 71096 28636 71102 28648
rect 62117 28611 62175 28617
rect 62117 28577 62129 28611
rect 62163 28577 62175 28611
rect 62117 28571 62175 28577
rect 62666 28568 62672 28620
rect 62724 28608 62730 28620
rect 78401 28611 78459 28617
rect 78401 28608 78413 28611
rect 62724 28580 78413 28608
rect 62724 28568 62730 28580
rect 78401 28577 78413 28580
rect 78447 28577 78459 28611
rect 78401 28571 78459 28577
rect 78670 28611 78728 28617
rect 78670 28577 78682 28611
rect 78716 28577 78728 28611
rect 78670 28571 78728 28577
rect 78770 28611 78828 28617
rect 78770 28577 78782 28611
rect 78816 28577 78828 28611
rect 78950 28608 78956 28620
rect 78911 28580 78956 28608
rect 78770 28571 78828 28577
rect 78033 28543 78091 28549
rect 78033 28540 78045 28543
rect 62040 28512 78045 28540
rect 78033 28509 78045 28512
rect 78079 28540 78091 28543
rect 78585 28543 78643 28549
rect 78585 28540 78597 28543
rect 78079 28512 78352 28540
rect 78079 28509 78091 28512
rect 78033 28503 78091 28509
rect 49510 28432 49516 28484
rect 49568 28472 49574 28484
rect 56318 28472 56324 28484
rect 49568 28444 56324 28472
rect 49568 28432 49574 28444
rect 56318 28432 56324 28444
rect 56376 28432 56382 28484
rect 56962 28432 56968 28484
rect 57020 28472 57026 28484
rect 59722 28472 59728 28484
rect 57020 28444 59728 28472
rect 57020 28432 57026 28444
rect 59722 28432 59728 28444
rect 59780 28432 59786 28484
rect 78217 28475 78275 28481
rect 78217 28472 78229 28475
rect 60706 28444 70394 28472
rect 47627 28376 47992 28404
rect 47627 28373 47639 28376
rect 47581 28367 47639 28373
rect 48038 28364 48044 28416
rect 48096 28404 48102 28416
rect 60706 28404 60734 28444
rect 48096 28376 60734 28404
rect 61933 28407 61991 28413
rect 48096 28364 48102 28376
rect 61933 28373 61945 28407
rect 61979 28404 61991 28407
rect 63126 28404 63132 28416
rect 61979 28376 63132 28404
rect 61979 28373 61991 28376
rect 61933 28367 61991 28373
rect 63126 28364 63132 28376
rect 63184 28364 63190 28416
rect 63218 28364 63224 28416
rect 63276 28404 63282 28416
rect 69474 28404 69480 28416
rect 63276 28376 69480 28404
rect 63276 28364 63282 28376
rect 69474 28364 69480 28376
rect 69532 28364 69538 28416
rect 70366 28404 70394 28444
rect 74368 28444 78229 28472
rect 74368 28404 74396 28444
rect 78217 28441 78229 28444
rect 78263 28441 78275 28475
rect 78217 28435 78275 28441
rect 70366 28376 74396 28404
rect 78324 28404 78352 28512
rect 78416 28512 78597 28540
rect 78416 28484 78444 28512
rect 78585 28509 78597 28512
rect 78631 28509 78643 28543
rect 78585 28503 78643 28509
rect 78692 28484 78720 28571
rect 78784 28540 78812 28571
rect 78950 28568 78956 28580
rect 79008 28568 79014 28620
rect 80026 28608 80054 28648
rect 81069 28611 81127 28617
rect 81069 28608 81081 28611
rect 80026 28580 81081 28608
rect 81069 28577 81081 28580
rect 81115 28577 81127 28611
rect 81069 28571 81127 28577
rect 78784 28512 78904 28540
rect 78398 28432 78404 28484
rect 78456 28432 78462 28484
rect 78674 28432 78680 28484
rect 78732 28432 78738 28484
rect 78876 28404 78904 28512
rect 79042 28432 79048 28484
rect 79100 28472 79106 28484
rect 94774 28472 94780 28484
rect 79100 28444 94780 28472
rect 79100 28432 79106 28444
rect 94774 28432 94780 28444
rect 94832 28432 94838 28484
rect 80882 28404 80888 28416
rect 78324 28376 78904 28404
rect 80843 28376 80888 28404
rect 80882 28364 80888 28376
rect 80940 28364 80946 28416
rect 1104 28314 98808 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 65686 28314
rect 65738 28262 65750 28314
rect 65802 28262 65814 28314
rect 65866 28262 65878 28314
rect 65930 28262 96406 28314
rect 96458 28262 96470 28314
rect 96522 28262 96534 28314
rect 96586 28262 96598 28314
rect 96650 28262 98808 28314
rect 1104 28240 98808 28262
rect 3602 28200 3608 28212
rect 3563 28172 3608 28200
rect 3602 28160 3608 28172
rect 3660 28160 3666 28212
rect 3786 28160 3792 28212
rect 3844 28200 3850 28212
rect 14274 28200 14280 28212
rect 3844 28172 14280 28200
rect 3844 28160 3850 28172
rect 14274 28160 14280 28172
rect 14332 28160 14338 28212
rect 14458 28200 14464 28212
rect 14419 28172 14464 28200
rect 14458 28160 14464 28172
rect 14516 28160 14522 28212
rect 14568 28172 22094 28200
rect 2498 28092 2504 28144
rect 2556 28132 2562 28144
rect 2556 28104 4016 28132
rect 2556 28092 2562 28104
rect 3988 28064 4016 28104
rect 5350 28092 5356 28144
rect 5408 28132 5414 28144
rect 13814 28132 13820 28144
rect 5408 28104 13820 28132
rect 5408 28092 5414 28104
rect 13814 28092 13820 28104
rect 13872 28092 13878 28144
rect 14568 28132 14596 28172
rect 14200 28104 14596 28132
rect 14200 28064 14228 28104
rect 16574 28092 16580 28144
rect 16632 28132 16638 28144
rect 17770 28132 17776 28144
rect 16632 28104 17776 28132
rect 16632 28092 16638 28104
rect 17770 28092 17776 28104
rect 17828 28092 17834 28144
rect 19886 28092 19892 28144
rect 19944 28141 19950 28144
rect 19944 28135 19993 28141
rect 19944 28101 19947 28135
rect 19981 28101 19993 28135
rect 20070 28132 20076 28144
rect 20031 28104 20076 28132
rect 19944 28095 19993 28101
rect 19944 28092 19950 28095
rect 20070 28092 20076 28104
rect 20128 28092 20134 28144
rect 22066 28132 22094 28172
rect 23382 28160 23388 28212
rect 23440 28200 23446 28212
rect 30006 28200 30012 28212
rect 23440 28172 30012 28200
rect 23440 28160 23446 28172
rect 30006 28160 30012 28172
rect 30064 28160 30070 28212
rect 30374 28160 30380 28212
rect 30432 28200 30438 28212
rect 38286 28200 38292 28212
rect 30432 28172 38292 28200
rect 30432 28160 30438 28172
rect 38286 28160 38292 28172
rect 38344 28160 38350 28212
rect 38933 28203 38991 28209
rect 38933 28169 38945 28203
rect 38979 28200 38991 28203
rect 39209 28203 39267 28209
rect 39209 28200 39221 28203
rect 38979 28172 39221 28200
rect 38979 28169 38991 28172
rect 38933 28163 38991 28169
rect 39209 28169 39221 28172
rect 39255 28200 39267 28203
rect 49510 28200 49516 28212
rect 39255 28172 49516 28200
rect 39255 28169 39267 28172
rect 39209 28163 39267 28169
rect 49510 28160 49516 28172
rect 49568 28160 49574 28212
rect 49694 28160 49700 28212
rect 49752 28200 49758 28212
rect 88610 28200 88616 28212
rect 49752 28172 88616 28200
rect 49752 28160 49758 28172
rect 88610 28160 88616 28172
rect 88668 28160 88674 28212
rect 39298 28132 39304 28144
rect 22066 28104 39304 28132
rect 39298 28092 39304 28104
rect 39356 28092 39362 28144
rect 39390 28092 39396 28144
rect 39448 28132 39454 28144
rect 46198 28132 46204 28144
rect 39448 28104 46204 28132
rect 39448 28092 39454 28104
rect 46198 28092 46204 28104
rect 46256 28092 46262 28144
rect 46290 28092 46296 28144
rect 46348 28132 46354 28144
rect 49786 28132 49792 28144
rect 46348 28104 49792 28132
rect 46348 28092 46354 28104
rect 49786 28092 49792 28104
rect 49844 28092 49850 28144
rect 49970 28092 49976 28144
rect 50028 28132 50034 28144
rect 62942 28132 62948 28144
rect 50028 28104 62948 28132
rect 50028 28092 50034 28104
rect 62942 28092 62948 28104
rect 63000 28092 63006 28144
rect 63034 28092 63040 28144
rect 63092 28132 63098 28144
rect 68370 28132 68376 28144
rect 63092 28104 68376 28132
rect 63092 28092 63098 28104
rect 68370 28092 68376 28104
rect 68428 28132 68434 28144
rect 68922 28132 68928 28144
rect 68428 28104 68928 28132
rect 68428 28092 68434 28104
rect 68922 28092 68928 28104
rect 68980 28092 68986 28144
rect 92566 28132 92572 28144
rect 87432 28104 92572 28132
rect 17402 28064 17408 28076
rect 3988 28036 14228 28064
rect 14292 28036 17264 28064
rect 17363 28036 17408 28064
rect 3786 27996 3792 28008
rect 3747 27968 3792 27996
rect 3786 27956 3792 27968
rect 3844 27956 3850 28008
rect 4062 27996 4068 28008
rect 4023 27968 4068 27996
rect 4062 27956 4068 27968
rect 4120 27956 4126 28008
rect 11790 27956 11796 28008
rect 11848 27996 11854 28008
rect 14292 28005 14320 28036
rect 14277 27999 14335 28005
rect 11848 27968 14228 27996
rect 11848 27956 11854 27968
rect 3513 27931 3571 27937
rect 3513 27897 3525 27931
rect 3559 27928 3571 27931
rect 13998 27928 14004 27940
rect 3559 27900 4016 27928
rect 13959 27900 14004 27928
rect 3559 27897 3571 27900
rect 3513 27891 3571 27897
rect 3988 27872 4016 27900
rect 13998 27888 14004 27900
rect 14056 27888 14062 27940
rect 3970 27860 3976 27872
rect 3931 27832 3976 27860
rect 3970 27820 3976 27832
rect 4028 27820 4034 27872
rect 13909 27863 13967 27869
rect 13909 27829 13921 27863
rect 13955 27860 13967 27863
rect 14090 27860 14096 27872
rect 13955 27832 14096 27860
rect 13955 27829 13967 27832
rect 13909 27823 13967 27829
rect 14090 27820 14096 27832
rect 14148 27820 14154 27872
rect 14200 27860 14228 27968
rect 14277 27965 14289 27999
rect 14323 27965 14335 27999
rect 14277 27959 14335 27965
rect 15102 27956 15108 28008
rect 15160 27996 15166 28008
rect 16758 27996 16764 28008
rect 15160 27968 16764 27996
rect 15160 27956 15166 27968
rect 16758 27956 16764 27968
rect 16816 27956 16822 28008
rect 17037 27999 17095 28005
rect 17037 27965 17049 27999
rect 17083 27996 17095 27999
rect 17126 27996 17132 28008
rect 17083 27968 17132 27996
rect 17083 27965 17095 27968
rect 17037 27959 17095 27965
rect 17126 27956 17132 27968
rect 17184 27956 17190 28008
rect 17236 27996 17264 28036
rect 17402 28024 17408 28036
rect 17460 28024 17466 28076
rect 20165 28067 20223 28073
rect 17512 28036 20116 28064
rect 17512 27996 17540 28036
rect 17236 27968 17540 27996
rect 18598 27956 18604 28008
rect 18656 27996 18662 28008
rect 18693 27999 18751 28005
rect 18693 27996 18705 27999
rect 18656 27968 18705 27996
rect 18656 27956 18662 27968
rect 18693 27965 18705 27968
rect 18739 27965 18751 27999
rect 18693 27959 18751 27965
rect 18874 27956 18880 28008
rect 18932 27996 18938 28008
rect 18969 27999 19027 28005
rect 18969 27996 18981 27999
rect 18932 27968 18981 27996
rect 18932 27956 18938 27968
rect 18969 27965 18981 27968
rect 19015 27965 19027 27999
rect 18969 27959 19027 27965
rect 19058 27956 19064 28008
rect 19116 27996 19122 28008
rect 20088 27996 20116 28036
rect 20165 28033 20177 28067
rect 20211 28064 20223 28067
rect 20254 28064 20260 28076
rect 20211 28036 20260 28064
rect 20211 28033 20223 28036
rect 20165 28027 20223 28033
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 24210 28024 24216 28076
rect 24268 28064 24274 28076
rect 64322 28064 64328 28076
rect 24268 28036 64328 28064
rect 24268 28024 24274 28036
rect 64322 28024 64328 28036
rect 64380 28024 64386 28076
rect 84194 28024 84200 28076
rect 84252 28064 84258 28076
rect 87432 28073 87460 28104
rect 92566 28092 92572 28104
rect 92624 28092 92630 28144
rect 87049 28067 87107 28073
rect 87049 28064 87061 28067
rect 84252 28036 87061 28064
rect 84252 28024 84258 28036
rect 87049 28033 87061 28036
rect 87095 28033 87107 28067
rect 87049 28027 87107 28033
rect 87417 28067 87475 28073
rect 87417 28033 87429 28067
rect 87463 28033 87475 28067
rect 87417 28027 87475 28033
rect 87509 28067 87567 28073
rect 87509 28033 87521 28067
rect 87555 28064 87567 28067
rect 92474 28064 92480 28076
rect 87555 28036 92480 28064
rect 87555 28033 87567 28036
rect 87509 28027 87567 28033
rect 92474 28024 92480 28036
rect 92532 28024 92538 28076
rect 22370 27996 22376 28008
rect 19116 27968 19932 27996
rect 20088 27968 22376 27996
rect 19116 27956 19122 27968
rect 19334 27888 19340 27940
rect 19392 27928 19398 27940
rect 19797 27931 19855 27937
rect 19797 27928 19809 27931
rect 19392 27900 19809 27928
rect 19392 27888 19398 27900
rect 19797 27897 19809 27900
rect 19843 27897 19855 27931
rect 19904 27928 19932 27968
rect 22370 27956 22376 27968
rect 22428 27996 22434 28008
rect 23290 27996 23296 28008
rect 22428 27968 23296 27996
rect 22428 27956 22434 27968
rect 23290 27956 23296 27968
rect 23348 27956 23354 28008
rect 26234 27956 26240 28008
rect 26292 27996 26298 28008
rect 32122 27996 32128 28008
rect 26292 27968 32128 27996
rect 26292 27956 26298 27968
rect 32122 27956 32128 27968
rect 32180 27956 32186 28008
rect 33134 27996 33140 28008
rect 33095 27968 33140 27996
rect 33134 27956 33140 27968
rect 33192 27956 33198 28008
rect 33520 27968 33778 27996
rect 33520 27928 33548 27968
rect 19904 27900 33548 27928
rect 19797 27891 19855 27897
rect 33594 27888 33600 27940
rect 33652 27928 33658 27940
rect 33750 27928 33778 27968
rect 34790 27956 34796 28008
rect 34848 27996 34854 28008
rect 38930 27996 38936 28008
rect 34848 27968 38936 27996
rect 34848 27956 34854 27968
rect 38930 27956 38936 27968
rect 38988 27956 38994 28008
rect 41506 27956 41512 28008
rect 41564 27996 41570 28008
rect 73798 27996 73804 28008
rect 41564 27968 73804 27996
rect 41564 27956 41570 27968
rect 73798 27956 73804 27968
rect 73856 27996 73862 28008
rect 74350 27996 74356 28008
rect 73856 27968 74356 27996
rect 73856 27956 73862 27968
rect 74350 27956 74356 27968
rect 74408 27956 74414 28008
rect 87233 27999 87291 28005
rect 87233 27996 87245 27999
rect 86972 27968 87245 27996
rect 51074 27928 51080 27940
rect 33652 27900 33697 27928
rect 33750 27900 51080 27928
rect 33652 27888 33658 27900
rect 51074 27888 51080 27900
rect 51132 27888 51138 27940
rect 51166 27888 51172 27940
rect 51224 27928 51230 27940
rect 69842 27928 69848 27940
rect 51224 27900 69848 27928
rect 51224 27888 51230 27900
rect 69842 27888 69848 27900
rect 69900 27888 69906 27940
rect 17954 27860 17960 27872
rect 14200 27832 17960 27860
rect 17954 27820 17960 27832
rect 18012 27820 18018 27872
rect 19150 27860 19156 27872
rect 19111 27832 19156 27860
rect 19150 27820 19156 27832
rect 19208 27820 19214 27872
rect 19242 27820 19248 27872
rect 19300 27860 19306 27872
rect 20441 27863 20499 27869
rect 20441 27860 20453 27863
rect 19300 27832 20453 27860
rect 19300 27820 19306 27832
rect 20441 27829 20453 27832
rect 20487 27829 20499 27863
rect 20441 27823 20499 27829
rect 20530 27820 20536 27872
rect 20588 27860 20594 27872
rect 74718 27860 74724 27872
rect 20588 27832 74724 27860
rect 20588 27820 20594 27832
rect 74718 27820 74724 27832
rect 74776 27820 74782 27872
rect 85574 27820 85580 27872
rect 85632 27860 85638 27872
rect 86972 27869 87000 27968
rect 87233 27965 87245 27968
rect 87279 27965 87291 27999
rect 87598 27996 87604 28008
rect 87559 27968 87604 27996
rect 87233 27959 87291 27965
rect 87598 27956 87604 27968
rect 87656 27956 87662 28008
rect 87690 27956 87696 28008
rect 87748 27996 87754 28008
rect 87785 27999 87843 28005
rect 87785 27996 87797 27999
rect 87748 27968 87797 27996
rect 87748 27956 87754 27968
rect 87785 27965 87797 27968
rect 87831 27965 87843 27999
rect 87785 27959 87843 27965
rect 86957 27863 87015 27869
rect 86957 27860 86969 27863
rect 85632 27832 86969 27860
rect 85632 27820 85638 27832
rect 86957 27829 86969 27832
rect 87003 27829 87015 27863
rect 86957 27823 87015 27829
rect 1104 27770 98808 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 50326 27770
rect 50378 27718 50390 27770
rect 50442 27718 50454 27770
rect 50506 27718 50518 27770
rect 50570 27718 81046 27770
rect 81098 27718 81110 27770
rect 81162 27718 81174 27770
rect 81226 27718 81238 27770
rect 81290 27718 98808 27770
rect 1104 27696 98808 27718
rect 3970 27616 3976 27668
rect 4028 27656 4034 27668
rect 20530 27656 20536 27668
rect 4028 27628 20536 27656
rect 4028 27616 4034 27628
rect 20530 27616 20536 27628
rect 20588 27616 20594 27668
rect 21358 27616 21364 27668
rect 21416 27656 21422 27668
rect 21542 27656 21548 27668
rect 21416 27628 21548 27656
rect 21416 27616 21422 27628
rect 21542 27616 21548 27628
rect 21600 27616 21606 27668
rect 23198 27616 23204 27668
rect 23256 27656 23262 27668
rect 28902 27656 28908 27668
rect 23256 27628 28908 27656
rect 23256 27616 23262 27628
rect 28902 27616 28908 27628
rect 28960 27616 28966 27668
rect 29086 27656 29092 27668
rect 29047 27628 29092 27656
rect 29086 27616 29092 27628
rect 29144 27616 29150 27668
rect 33502 27616 33508 27668
rect 33560 27656 33566 27668
rect 38010 27656 38016 27668
rect 33560 27628 38016 27656
rect 33560 27616 33566 27628
rect 38010 27616 38016 27628
rect 38068 27616 38074 27668
rect 38672 27628 39344 27656
rect 11790 27588 11796 27600
rect 11751 27560 11796 27588
rect 11790 27548 11796 27560
rect 11848 27548 11854 27600
rect 15194 27588 15200 27600
rect 12360 27560 15200 27588
rect 11057 27523 11115 27529
rect 11057 27489 11069 27523
rect 11103 27489 11115 27523
rect 11238 27520 11244 27532
rect 11199 27492 11244 27520
rect 11057 27483 11115 27489
rect 11072 27452 11100 27483
rect 11238 27480 11244 27492
rect 11296 27480 11302 27532
rect 11514 27520 11520 27532
rect 11475 27492 11520 27520
rect 11514 27480 11520 27492
rect 11572 27480 11578 27532
rect 11698 27520 11704 27532
rect 11659 27492 11704 27520
rect 11698 27480 11704 27492
rect 11756 27480 11762 27532
rect 12253 27523 12311 27529
rect 12253 27489 12265 27523
rect 12299 27489 12311 27523
rect 12253 27483 12311 27489
rect 11146 27452 11152 27464
rect 11072 27424 11152 27452
rect 11146 27412 11152 27424
rect 11204 27412 11210 27464
rect 12268 27316 12296 27483
rect 12360 27452 12388 27560
rect 15194 27548 15200 27560
rect 15252 27548 15258 27600
rect 26142 27588 26148 27600
rect 19076 27560 26148 27588
rect 12437 27523 12495 27529
rect 12437 27489 12449 27523
rect 12483 27520 12495 27523
rect 12483 27492 12756 27520
rect 12483 27489 12495 27492
rect 12437 27483 12495 27489
rect 12529 27455 12587 27461
rect 12529 27452 12541 27455
rect 12360 27424 12541 27452
rect 12529 27421 12541 27424
rect 12575 27421 12587 27455
rect 12529 27415 12587 27421
rect 12621 27455 12679 27461
rect 12621 27421 12633 27455
rect 12667 27421 12679 27455
rect 12728 27452 12756 27492
rect 12802 27480 12808 27532
rect 12860 27520 12866 27532
rect 16117 27523 16175 27529
rect 12860 27492 12905 27520
rect 12860 27480 12866 27492
rect 16117 27489 16129 27523
rect 16163 27520 16175 27523
rect 19076 27520 19104 27560
rect 26142 27548 26148 27560
rect 26200 27548 26206 27600
rect 33318 27588 33324 27600
rect 28828 27560 33324 27588
rect 23658 27520 23664 27532
rect 16163 27492 19104 27520
rect 23619 27492 23664 27520
rect 16163 27489 16175 27492
rect 16117 27483 16175 27489
rect 23658 27480 23664 27492
rect 23716 27480 23722 27532
rect 27798 27520 27804 27532
rect 27759 27492 27804 27520
rect 27798 27480 27804 27492
rect 27856 27480 27862 27532
rect 27890 27480 27896 27532
rect 27948 27520 27954 27532
rect 28828 27520 28856 27560
rect 33318 27548 33324 27560
rect 33376 27548 33382 27600
rect 34330 27548 34336 27600
rect 34388 27588 34394 27600
rect 35894 27588 35900 27600
rect 34388 27560 35900 27588
rect 34388 27548 34394 27560
rect 35894 27548 35900 27560
rect 35952 27548 35958 27600
rect 35986 27548 35992 27600
rect 36044 27588 36050 27600
rect 38562 27588 38568 27600
rect 36044 27560 38568 27588
rect 36044 27548 36050 27560
rect 38562 27548 38568 27560
rect 38620 27548 38626 27600
rect 27948 27492 28856 27520
rect 27948 27480 27954 27492
rect 28902 27480 28908 27532
rect 28960 27520 28966 27532
rect 30374 27520 30380 27532
rect 28960 27492 30380 27520
rect 28960 27480 28966 27492
rect 30374 27480 30380 27492
rect 30432 27480 30438 27532
rect 30466 27480 30472 27532
rect 30524 27520 30530 27532
rect 38672 27520 38700 27628
rect 38746 27548 38752 27600
rect 38804 27588 38810 27600
rect 39316 27588 39344 27628
rect 40034 27616 40040 27668
rect 40092 27656 40098 27668
rect 41230 27656 41236 27668
rect 40092 27628 41236 27656
rect 40092 27616 40098 27628
rect 41230 27616 41236 27628
rect 41288 27616 41294 27668
rect 41414 27616 41420 27668
rect 41472 27656 41478 27668
rect 41472 27628 42012 27656
rect 41472 27616 41478 27628
rect 41984 27588 42012 27628
rect 46198 27616 46204 27668
rect 46256 27656 46262 27668
rect 51074 27656 51080 27668
rect 46256 27628 51080 27656
rect 46256 27616 46262 27628
rect 51074 27616 51080 27628
rect 51132 27616 51138 27668
rect 51166 27616 51172 27668
rect 51224 27656 51230 27668
rect 53837 27659 53895 27665
rect 53837 27656 53849 27659
rect 51224 27628 53849 27656
rect 51224 27616 51230 27628
rect 53837 27625 53849 27628
rect 53883 27625 53895 27659
rect 53837 27619 53895 27625
rect 53926 27616 53932 27668
rect 53984 27656 53990 27668
rect 59354 27656 59360 27668
rect 53984 27628 59360 27656
rect 53984 27616 53990 27628
rect 59354 27616 59360 27628
rect 59412 27616 59418 27668
rect 61838 27616 61844 27668
rect 61896 27656 61902 27668
rect 69750 27656 69756 27668
rect 61896 27628 69756 27656
rect 61896 27616 61902 27628
rect 69750 27616 69756 27628
rect 69808 27656 69814 27668
rect 74258 27656 74264 27668
rect 69808 27628 74264 27656
rect 69808 27616 69814 27628
rect 74258 27616 74264 27628
rect 74316 27616 74322 27668
rect 50614 27588 50620 27600
rect 38804 27560 39252 27588
rect 39316 27560 41920 27588
rect 41984 27560 50620 27588
rect 38804 27548 38810 27560
rect 30524 27492 38700 27520
rect 38933 27523 38991 27529
rect 30524 27480 30530 27492
rect 38933 27489 38945 27523
rect 38979 27520 38991 27523
rect 39022 27520 39028 27532
rect 38979 27492 39028 27520
rect 38979 27489 38991 27492
rect 38933 27483 38991 27489
rect 39022 27480 39028 27492
rect 39080 27480 39086 27532
rect 39224 27529 39252 27560
rect 39117 27523 39175 27529
rect 39117 27489 39129 27523
rect 39163 27489 39175 27523
rect 39117 27483 39175 27489
rect 39209 27523 39267 27529
rect 39209 27489 39221 27523
rect 39255 27489 39267 27523
rect 39209 27483 39267 27489
rect 39485 27523 39543 27529
rect 39485 27489 39497 27523
rect 39531 27520 39543 27523
rect 39574 27520 39580 27532
rect 39531 27492 39580 27520
rect 39531 27489 39543 27492
rect 39485 27483 39543 27489
rect 13906 27452 13912 27464
rect 12728 27424 13912 27452
rect 12621 27415 12679 27421
rect 12636 27384 12664 27415
rect 13906 27412 13912 27424
rect 13964 27452 13970 27464
rect 14366 27452 14372 27464
rect 13964 27424 14372 27452
rect 13964 27412 13970 27424
rect 14366 27412 14372 27424
rect 14424 27412 14430 27464
rect 15838 27452 15844 27464
rect 15799 27424 15844 27452
rect 15838 27412 15844 27424
rect 15896 27412 15902 27464
rect 16022 27412 16028 27464
rect 16080 27452 16086 27464
rect 22002 27452 22008 27464
rect 16080 27424 22008 27452
rect 16080 27412 16086 27424
rect 22002 27412 22008 27424
rect 22060 27412 22066 27464
rect 27522 27452 27528 27464
rect 27483 27424 27528 27452
rect 27522 27412 27528 27424
rect 27580 27412 27586 27464
rect 32674 27452 32680 27464
rect 28552 27424 32680 27452
rect 15470 27384 15476 27396
rect 12636 27356 15476 27384
rect 15470 27344 15476 27356
rect 15528 27344 15534 27396
rect 17144 27356 22094 27384
rect 12710 27316 12716 27328
rect 12268 27288 12716 27316
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 12986 27316 12992 27328
rect 12947 27288 12992 27316
rect 12986 27276 12992 27288
rect 13044 27276 13050 27328
rect 15013 27319 15071 27325
rect 15013 27285 15025 27319
rect 15059 27316 15071 27319
rect 15289 27319 15347 27325
rect 15289 27316 15301 27319
rect 15059 27288 15301 27316
rect 15059 27285 15071 27288
rect 15013 27279 15071 27285
rect 15289 27285 15301 27288
rect 15335 27316 15347 27319
rect 17144 27316 17172 27356
rect 15335 27288 17172 27316
rect 17405 27319 17463 27325
rect 15335 27285 15347 27288
rect 15289 27279 15347 27285
rect 17405 27285 17417 27319
rect 17451 27316 17463 27319
rect 17586 27316 17592 27328
rect 17451 27288 17592 27316
rect 17451 27285 17463 27288
rect 17405 27279 17463 27285
rect 17586 27276 17592 27288
rect 17644 27316 17650 27328
rect 21910 27316 21916 27328
rect 17644 27288 21916 27316
rect 17644 27276 17650 27288
rect 21910 27276 21916 27288
rect 21968 27276 21974 27328
rect 22066 27316 22094 27356
rect 23014 27344 23020 27396
rect 23072 27384 23078 27396
rect 27154 27384 27160 27396
rect 23072 27356 27160 27384
rect 23072 27344 23078 27356
rect 27154 27344 27160 27356
rect 27212 27344 27218 27396
rect 28552 27316 28580 27424
rect 32674 27412 32680 27424
rect 32732 27412 32738 27464
rect 35250 27412 35256 27464
rect 35308 27452 35314 27464
rect 38010 27452 38016 27464
rect 35308 27424 38016 27452
rect 35308 27412 35314 27424
rect 38010 27412 38016 27424
rect 38068 27412 38074 27464
rect 38838 27412 38844 27464
rect 38896 27452 38902 27464
rect 39132 27452 39160 27483
rect 39574 27480 39580 27492
rect 39632 27520 39638 27532
rect 41233 27523 41291 27529
rect 39632 27492 41184 27520
rect 39632 27480 39638 27492
rect 39298 27452 39304 27464
rect 38896 27424 39160 27452
rect 39259 27424 39304 27452
rect 38896 27412 38902 27424
rect 39298 27412 39304 27424
rect 39356 27412 39362 27464
rect 39666 27452 39672 27464
rect 39627 27424 39672 27452
rect 39666 27412 39672 27424
rect 39724 27412 39730 27464
rect 28626 27344 28632 27396
rect 28684 27384 28690 27396
rect 40494 27384 40500 27396
rect 28684 27356 40500 27384
rect 28684 27344 28690 27356
rect 40494 27344 40500 27356
rect 40552 27344 40558 27396
rect 41156 27384 41184 27492
rect 41233 27489 41245 27523
rect 41279 27520 41291 27523
rect 41506 27520 41512 27532
rect 41279 27492 41512 27520
rect 41279 27489 41291 27492
rect 41233 27483 41291 27489
rect 41506 27480 41512 27492
rect 41564 27480 41570 27532
rect 41892 27529 41920 27560
rect 50614 27548 50620 27560
rect 50672 27548 50678 27600
rect 50706 27548 50712 27600
rect 50764 27588 50770 27600
rect 52822 27588 52828 27600
rect 50764 27560 52828 27588
rect 50764 27548 50770 27560
rect 52822 27548 52828 27560
rect 52880 27548 52886 27600
rect 53116 27560 60734 27588
rect 41785 27523 41843 27529
rect 41785 27489 41797 27523
rect 41831 27489 41843 27523
rect 41785 27483 41843 27489
rect 41877 27523 41935 27529
rect 41877 27489 41889 27523
rect 41923 27489 41935 27523
rect 42058 27520 42064 27532
rect 42019 27492 42064 27520
rect 41877 27483 41935 27489
rect 41690 27452 41696 27464
rect 41651 27424 41696 27452
rect 41690 27412 41696 27424
rect 41748 27412 41754 27464
rect 41800 27396 41828 27483
rect 42058 27480 42064 27492
rect 42116 27480 42122 27532
rect 53116 27520 53144 27560
rect 42168 27492 53144 27520
rect 53193 27523 53251 27529
rect 41156 27356 41460 27384
rect 22066 27288 28580 27316
rect 28994 27276 29000 27328
rect 29052 27316 29058 27328
rect 31018 27316 31024 27328
rect 29052 27288 31024 27316
rect 29052 27276 29058 27288
rect 31018 27276 31024 27288
rect 31076 27276 31082 27328
rect 33870 27276 33876 27328
rect 33928 27316 33934 27328
rect 37642 27316 37648 27328
rect 33928 27288 37648 27316
rect 33928 27276 33934 27288
rect 37642 27276 37648 27288
rect 37700 27276 37706 27328
rect 38010 27276 38016 27328
rect 38068 27316 38074 27328
rect 40954 27316 40960 27328
rect 38068 27288 40960 27316
rect 38068 27276 38074 27288
rect 40954 27276 40960 27288
rect 41012 27276 41018 27328
rect 41322 27316 41328 27328
rect 41283 27288 41328 27316
rect 41322 27276 41328 27288
rect 41380 27276 41386 27328
rect 41432 27316 41460 27356
rect 41782 27344 41788 27396
rect 41840 27344 41846 27396
rect 42168 27316 42196 27492
rect 53193 27489 53205 27523
rect 53239 27520 53251 27523
rect 53282 27520 53288 27532
rect 53239 27492 53288 27520
rect 53239 27489 53251 27492
rect 53193 27483 53251 27489
rect 53282 27480 53288 27492
rect 53340 27480 53346 27532
rect 53374 27480 53380 27532
rect 53432 27520 53438 27532
rect 53432 27492 53476 27520
rect 53432 27480 53438 27492
rect 53742 27480 53748 27532
rect 53800 27520 53806 27532
rect 53800 27492 53845 27520
rect 53800 27480 53806 27492
rect 53926 27480 53932 27532
rect 53984 27520 53990 27532
rect 60706 27520 60734 27560
rect 72050 27548 72056 27600
rect 72108 27588 72114 27600
rect 76742 27588 76748 27600
rect 72108 27560 76748 27588
rect 72108 27548 72114 27560
rect 76742 27548 76748 27560
rect 76800 27548 76806 27600
rect 91646 27520 91652 27532
rect 53984 27492 60596 27520
rect 60706 27492 91652 27520
rect 53984 27480 53990 27492
rect 46198 27412 46204 27464
rect 46256 27452 46262 27464
rect 53469 27455 53527 27461
rect 53469 27452 53481 27455
rect 46256 27424 53481 27452
rect 46256 27412 46262 27424
rect 53469 27421 53481 27424
rect 53515 27421 53527 27455
rect 53469 27415 53527 27421
rect 53561 27455 53619 27461
rect 53561 27421 53573 27455
rect 53607 27421 53619 27455
rect 53561 27415 53619 27421
rect 42518 27344 42524 27396
rect 42576 27384 42582 27396
rect 50706 27384 50712 27396
rect 42576 27356 50712 27384
rect 42576 27344 42582 27356
rect 50706 27344 50712 27356
rect 50764 27344 50770 27396
rect 53098 27384 53104 27396
rect 50816 27356 53104 27384
rect 41432 27288 42196 27316
rect 42794 27276 42800 27328
rect 42852 27316 42858 27328
rect 50816 27316 50844 27356
rect 53098 27344 53104 27356
rect 53156 27344 53162 27396
rect 42852 27288 50844 27316
rect 42852 27276 42858 27288
rect 52362 27276 52368 27328
rect 52420 27316 52426 27328
rect 53576 27316 53604 27415
rect 53834 27412 53840 27464
rect 53892 27452 53898 27464
rect 60458 27452 60464 27464
rect 53892 27424 60464 27452
rect 53892 27412 53898 27424
rect 60458 27412 60464 27424
rect 60516 27412 60522 27464
rect 60568 27452 60596 27492
rect 91646 27480 91652 27492
rect 91704 27480 91710 27532
rect 72142 27452 72148 27464
rect 60568 27424 72148 27452
rect 72142 27412 72148 27424
rect 72200 27412 72206 27464
rect 78306 27412 78312 27464
rect 78364 27452 78370 27464
rect 79318 27452 79324 27464
rect 78364 27424 79324 27452
rect 78364 27412 78370 27424
rect 79318 27412 79324 27424
rect 79376 27412 79382 27464
rect 79594 27452 79600 27464
rect 79555 27424 79600 27452
rect 79594 27412 79600 27424
rect 79652 27412 79658 27464
rect 83550 27412 83556 27464
rect 83608 27452 83614 27464
rect 86862 27452 86868 27464
rect 83608 27424 86868 27452
rect 83608 27412 83614 27424
rect 86862 27412 86868 27424
rect 86920 27412 86926 27464
rect 53650 27344 53656 27396
rect 53708 27384 53714 27396
rect 72602 27384 72608 27396
rect 53708 27356 72608 27384
rect 53708 27344 53714 27356
rect 72602 27344 72608 27356
rect 72660 27344 72666 27396
rect 83274 27344 83280 27396
rect 83332 27384 83338 27396
rect 87046 27384 87052 27396
rect 83332 27356 87052 27384
rect 83332 27344 83338 27356
rect 87046 27344 87052 27356
rect 87104 27344 87110 27396
rect 53926 27316 53932 27328
rect 52420 27288 53932 27316
rect 52420 27276 52426 27288
rect 53926 27276 53932 27288
rect 53984 27276 53990 27328
rect 55674 27276 55680 27328
rect 55732 27316 55738 27328
rect 60642 27316 60648 27328
rect 55732 27288 60648 27316
rect 55732 27276 55738 27288
rect 60642 27276 60648 27288
rect 60700 27276 60706 27328
rect 60918 27276 60924 27328
rect 60976 27316 60982 27328
rect 68094 27316 68100 27328
rect 60976 27288 68100 27316
rect 60976 27276 60982 27288
rect 68094 27276 68100 27288
rect 68152 27276 68158 27328
rect 74350 27276 74356 27328
rect 74408 27316 74414 27328
rect 80701 27319 80759 27325
rect 80701 27316 80713 27319
rect 74408 27288 80713 27316
rect 74408 27276 74414 27288
rect 80701 27285 80713 27288
rect 80747 27285 80759 27319
rect 80701 27279 80759 27285
rect 84838 27276 84844 27328
rect 84896 27316 84902 27328
rect 94406 27316 94412 27328
rect 84896 27288 94412 27316
rect 84896 27276 84902 27288
rect 94406 27276 94412 27288
rect 94464 27276 94470 27328
rect 1104 27226 98808 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 65686 27226
rect 65738 27174 65750 27226
rect 65802 27174 65814 27226
rect 65866 27174 65878 27226
rect 65930 27174 96406 27226
rect 96458 27174 96470 27226
rect 96522 27174 96534 27226
rect 96586 27174 96598 27226
rect 96650 27174 98808 27226
rect 1104 27152 98808 27174
rect 12710 27072 12716 27124
rect 12768 27112 12774 27124
rect 14182 27112 14188 27124
rect 12768 27084 14188 27112
rect 12768 27072 12774 27084
rect 14182 27072 14188 27084
rect 14240 27072 14246 27124
rect 15930 27072 15936 27124
rect 15988 27112 15994 27124
rect 17586 27112 17592 27124
rect 15988 27084 17592 27112
rect 15988 27072 15994 27084
rect 17586 27072 17592 27084
rect 17644 27072 17650 27124
rect 18138 27072 18144 27124
rect 18196 27112 18202 27124
rect 19886 27112 19892 27124
rect 18196 27084 19892 27112
rect 18196 27072 18202 27084
rect 19886 27072 19892 27084
rect 19944 27112 19950 27124
rect 21634 27112 21640 27124
rect 19944 27084 21640 27112
rect 19944 27072 19950 27084
rect 21634 27072 21640 27084
rect 21692 27072 21698 27124
rect 21818 27072 21824 27124
rect 21876 27112 21882 27124
rect 28626 27112 28632 27124
rect 21876 27084 28632 27112
rect 21876 27072 21882 27084
rect 28626 27072 28632 27084
rect 28684 27072 28690 27124
rect 28902 27072 28908 27124
rect 28960 27112 28966 27124
rect 35250 27112 35256 27124
rect 28960 27084 35256 27112
rect 28960 27072 28966 27084
rect 35250 27072 35256 27084
rect 35308 27072 35314 27124
rect 37642 27072 37648 27124
rect 37700 27112 37706 27124
rect 46198 27112 46204 27124
rect 37700 27084 46204 27112
rect 37700 27072 37706 27084
rect 46198 27072 46204 27084
rect 46256 27072 46262 27124
rect 46290 27072 46296 27124
rect 46348 27112 46354 27124
rect 55674 27112 55680 27124
rect 46348 27084 55680 27112
rect 46348 27072 46354 27084
rect 55674 27072 55680 27084
rect 55732 27072 55738 27124
rect 55876 27084 60596 27112
rect 7282 27004 7288 27056
rect 7340 27044 7346 27056
rect 21542 27044 21548 27056
rect 7340 27016 21548 27044
rect 7340 27004 7346 27016
rect 21542 27004 21548 27016
rect 21600 27004 21606 27056
rect 22278 27004 22284 27056
rect 22336 27044 22342 27056
rect 41414 27044 41420 27056
rect 22336 27016 41420 27044
rect 22336 27004 22342 27016
rect 41414 27004 41420 27016
rect 41472 27004 41478 27056
rect 43346 27004 43352 27056
rect 43404 27044 43410 27056
rect 55876 27044 55904 27084
rect 43404 27016 55904 27044
rect 43404 27004 43410 27016
rect 56042 27004 56048 27056
rect 56100 27044 56106 27056
rect 60568 27044 60596 27084
rect 60642 27072 60648 27124
rect 60700 27112 60706 27124
rect 84838 27112 84844 27124
rect 60700 27084 84844 27112
rect 60700 27072 60706 27084
rect 84838 27072 84844 27084
rect 84896 27072 84902 27124
rect 85040 27084 97396 27112
rect 75086 27044 75092 27056
rect 56100 27016 59676 27044
rect 60568 27016 75092 27044
rect 56100 27004 56106 27016
rect 14090 26936 14096 26988
rect 14148 26976 14154 26988
rect 21818 26976 21824 26988
rect 14148 26948 21824 26976
rect 14148 26936 14154 26948
rect 21818 26936 21824 26948
rect 21876 26936 21882 26988
rect 22002 26936 22008 26988
rect 22060 26976 22066 26988
rect 28994 26976 29000 26988
rect 22060 26948 29000 26976
rect 22060 26936 22066 26948
rect 28994 26936 29000 26948
rect 29052 26936 29058 26988
rect 29914 26936 29920 26988
rect 29972 26976 29978 26988
rect 30282 26976 30288 26988
rect 29972 26948 30288 26976
rect 29972 26936 29978 26948
rect 30282 26936 30288 26948
rect 30340 26936 30346 26988
rect 36170 26936 36176 26988
rect 36228 26976 36234 26988
rect 36630 26976 36636 26988
rect 36228 26948 36636 26976
rect 36228 26936 36234 26948
rect 36630 26936 36636 26948
rect 36688 26936 36694 26988
rect 38930 26936 38936 26988
rect 38988 26976 38994 26988
rect 39666 26976 39672 26988
rect 38988 26948 39672 26976
rect 38988 26936 38994 26948
rect 39666 26936 39672 26948
rect 39724 26936 39730 26988
rect 40402 26936 40408 26988
rect 40460 26976 40466 26988
rect 40862 26976 40868 26988
rect 40460 26948 40868 26976
rect 40460 26936 40466 26948
rect 40862 26936 40868 26948
rect 40920 26936 40926 26988
rect 40954 26936 40960 26988
rect 41012 26976 41018 26988
rect 59170 26976 59176 26988
rect 41012 26948 59176 26976
rect 41012 26936 41018 26948
rect 59170 26936 59176 26948
rect 59228 26936 59234 26988
rect 59648 26985 59676 27016
rect 75086 27004 75092 27016
rect 75144 27004 75150 27056
rect 77662 27004 77668 27056
rect 77720 27044 77726 27056
rect 78214 27044 78220 27056
rect 77720 27016 78220 27044
rect 77720 27004 77726 27016
rect 78214 27004 78220 27016
rect 78272 27044 78278 27056
rect 78493 27047 78551 27053
rect 78493 27044 78505 27047
rect 78272 27016 78505 27044
rect 78272 27004 78278 27016
rect 78493 27013 78505 27016
rect 78539 27013 78551 27047
rect 78493 27007 78551 27013
rect 79318 27004 79324 27056
rect 79376 27044 79382 27056
rect 80882 27044 80888 27056
rect 79376 27016 80888 27044
rect 79376 27004 79382 27016
rect 80882 27004 80888 27016
rect 80940 27004 80946 27056
rect 59633 26979 59691 26985
rect 59633 26945 59645 26979
rect 59679 26945 59691 26979
rect 61194 26976 61200 26988
rect 59633 26939 59691 26945
rect 59832 26948 60136 26976
rect 61155 26948 61200 26976
rect 17310 26868 17316 26920
rect 17368 26908 17374 26920
rect 17862 26908 17868 26920
rect 17368 26880 17868 26908
rect 17368 26868 17374 26880
rect 17862 26868 17868 26880
rect 17920 26868 17926 26920
rect 21082 26868 21088 26920
rect 21140 26908 21146 26920
rect 35986 26908 35992 26920
rect 21140 26880 35992 26908
rect 21140 26868 21146 26880
rect 35986 26868 35992 26880
rect 36044 26868 36050 26920
rect 37182 26908 37188 26920
rect 36096 26880 37188 26908
rect 5350 26800 5356 26852
rect 5408 26840 5414 26852
rect 23198 26840 23204 26852
rect 5408 26812 23204 26840
rect 5408 26800 5414 26812
rect 23198 26800 23204 26812
rect 23256 26800 23262 26852
rect 27522 26800 27528 26852
rect 27580 26840 27586 26852
rect 30834 26840 30840 26852
rect 27580 26812 30840 26840
rect 27580 26800 27586 26812
rect 30834 26800 30840 26812
rect 30892 26800 30898 26852
rect 30926 26800 30932 26852
rect 30984 26840 30990 26852
rect 36096 26840 36124 26880
rect 37182 26868 37188 26880
rect 37240 26868 37246 26920
rect 37274 26868 37280 26920
rect 37332 26908 37338 26920
rect 37918 26908 37924 26920
rect 37332 26880 37924 26908
rect 37332 26868 37338 26880
rect 37918 26868 37924 26880
rect 37976 26868 37982 26920
rect 38654 26868 38660 26920
rect 38712 26908 38718 26920
rect 39301 26911 39359 26917
rect 39301 26908 39313 26911
rect 38712 26880 39313 26908
rect 38712 26868 38718 26880
rect 39301 26877 39313 26880
rect 39347 26908 39359 26911
rect 39390 26908 39396 26920
rect 39347 26880 39396 26908
rect 39347 26877 39359 26880
rect 39301 26871 39359 26877
rect 39390 26868 39396 26880
rect 39448 26868 39454 26920
rect 39853 26911 39911 26917
rect 39853 26877 39865 26911
rect 39899 26908 39911 26911
rect 41598 26908 41604 26920
rect 39899 26880 41604 26908
rect 39899 26877 39911 26880
rect 39853 26871 39911 26877
rect 41598 26868 41604 26880
rect 41656 26868 41662 26920
rect 41874 26868 41880 26920
rect 41932 26908 41938 26920
rect 48222 26908 48228 26920
rect 41932 26880 48228 26908
rect 41932 26868 41938 26880
rect 48222 26868 48228 26880
rect 48280 26868 48286 26920
rect 48406 26868 48412 26920
rect 48464 26908 48470 26920
rect 49234 26908 49240 26920
rect 48464 26880 49240 26908
rect 48464 26868 48470 26880
rect 49234 26868 49240 26880
rect 49292 26868 49298 26920
rect 49878 26868 49884 26920
rect 49936 26908 49942 26920
rect 50706 26908 50712 26920
rect 49936 26880 50712 26908
rect 49936 26868 49942 26880
rect 50706 26868 50712 26880
rect 50764 26868 50770 26920
rect 52546 26908 52552 26920
rect 51046 26880 52552 26908
rect 30984 26812 36124 26840
rect 30984 26800 30990 26812
rect 36354 26800 36360 26852
rect 36412 26840 36418 26852
rect 51046 26840 51074 26880
rect 52546 26868 52552 26880
rect 52604 26868 52610 26920
rect 52638 26868 52644 26920
rect 52696 26908 52702 26920
rect 53466 26908 53472 26920
rect 52696 26880 53472 26908
rect 52696 26868 52702 26880
rect 53466 26868 53472 26880
rect 53524 26868 53530 26920
rect 54202 26868 54208 26920
rect 54260 26908 54266 26920
rect 54938 26908 54944 26920
rect 54260 26880 54944 26908
rect 54260 26868 54266 26880
rect 54938 26868 54944 26880
rect 54996 26868 55002 26920
rect 55030 26868 55036 26920
rect 55088 26908 55094 26920
rect 59832 26908 59860 26948
rect 55088 26880 59860 26908
rect 55088 26868 55094 26880
rect 59906 26868 59912 26920
rect 59964 26908 59970 26920
rect 60108 26908 60136 26948
rect 61194 26936 61200 26948
rect 61252 26936 61258 26988
rect 85040 26976 85068 27084
rect 87506 27004 87512 27056
rect 87564 27044 87570 27056
rect 94314 27044 94320 27056
rect 87564 27016 94320 27044
rect 87564 27004 87570 27016
rect 94314 27004 94320 27016
rect 94372 27004 94378 27056
rect 94774 27044 94780 27056
rect 94735 27016 94780 27044
rect 94774 27004 94780 27016
rect 94832 27004 94838 27056
rect 86218 26976 86224 26988
rect 70366 26948 85068 26976
rect 85408 26948 86224 26976
rect 70366 26908 70394 26948
rect 59964 26880 60009 26908
rect 60108 26880 70394 26908
rect 59964 26868 59970 26880
rect 75546 26868 75552 26920
rect 75604 26908 75610 26920
rect 77386 26908 77392 26920
rect 75604 26880 77392 26908
rect 75604 26868 75610 26880
rect 77386 26868 77392 26880
rect 77444 26868 77450 26920
rect 77849 26911 77907 26917
rect 77849 26908 77861 26911
rect 77588 26880 77861 26908
rect 36412 26812 51074 26840
rect 36412 26800 36418 26812
rect 52822 26800 52828 26852
rect 52880 26840 52886 26852
rect 59262 26840 59268 26852
rect 52880 26812 59268 26840
rect 52880 26800 52886 26812
rect 59262 26800 59268 26812
rect 59320 26800 59326 26852
rect 60706 26812 61148 26840
rect 17954 26732 17960 26784
rect 18012 26772 18018 26784
rect 60706 26772 60734 26812
rect 18012 26744 60734 26772
rect 61120 26772 61148 26812
rect 63034 26800 63040 26852
rect 63092 26840 63098 26852
rect 68830 26840 68836 26852
rect 63092 26812 68836 26840
rect 63092 26800 63098 26812
rect 68830 26800 68836 26812
rect 68888 26800 68894 26852
rect 69014 26800 69020 26852
rect 69072 26840 69078 26852
rect 77018 26840 77024 26852
rect 69072 26812 77024 26840
rect 69072 26800 69078 26812
rect 77018 26800 77024 26812
rect 77076 26800 77082 26852
rect 77588 26772 77616 26880
rect 77849 26877 77861 26880
rect 77895 26908 77907 26911
rect 78079 26911 78137 26917
rect 78079 26908 78091 26911
rect 77895 26880 78091 26908
rect 77895 26877 77907 26880
rect 77849 26871 77907 26877
rect 78079 26877 78091 26880
rect 78125 26877 78137 26911
rect 78214 26908 78220 26920
rect 78175 26880 78220 26908
rect 78079 26871 78137 26877
rect 78214 26868 78220 26880
rect 78272 26868 78278 26920
rect 80882 26868 80888 26920
rect 80940 26908 80946 26920
rect 85408 26908 85436 26948
rect 86218 26936 86224 26948
rect 86276 26976 86282 26988
rect 86313 26979 86371 26985
rect 86313 26976 86325 26979
rect 86276 26948 86325 26976
rect 86276 26936 86282 26948
rect 86313 26945 86325 26948
rect 86359 26945 86371 26979
rect 86313 26939 86371 26945
rect 86494 26936 86500 26988
rect 86552 26976 86558 26988
rect 86589 26979 86647 26985
rect 86589 26976 86601 26979
rect 86552 26948 86601 26976
rect 86552 26936 86558 26948
rect 86589 26945 86601 26948
rect 86635 26945 86647 26979
rect 86589 26939 86647 26945
rect 87414 26936 87420 26988
rect 87472 26976 87478 26988
rect 97368 26985 97396 27084
rect 97353 26979 97411 26985
rect 87472 26948 97120 26976
rect 87472 26936 87478 26948
rect 86678 26908 86684 26920
rect 80940 26880 85436 26908
rect 86420 26880 86684 26908
rect 80940 26868 80946 26880
rect 78490 26800 78496 26852
rect 78548 26840 78554 26852
rect 86420 26840 86448 26880
rect 86678 26868 86684 26880
rect 86736 26868 86742 26920
rect 86862 26868 86868 26920
rect 86920 26908 86926 26920
rect 94225 26911 94283 26917
rect 94225 26908 94237 26911
rect 86920 26880 94237 26908
rect 86920 26868 86926 26880
rect 94225 26877 94237 26880
rect 94271 26877 94283 26911
rect 94498 26908 94504 26920
rect 94459 26880 94504 26908
rect 94225 26871 94283 26877
rect 94498 26868 94504 26880
rect 94556 26868 94562 26920
rect 94593 26911 94651 26917
rect 94593 26877 94605 26911
rect 94639 26877 94651 26911
rect 94593 26871 94651 26877
rect 94409 26843 94467 26849
rect 94409 26840 94421 26843
rect 78548 26812 86448 26840
rect 87248 26812 94421 26840
rect 78548 26800 78554 26812
rect 78122 26772 78128 26784
rect 61120 26744 77616 26772
rect 78083 26744 78128 26772
rect 18012 26732 18018 26744
rect 78122 26732 78128 26744
rect 78180 26732 78186 26784
rect 79410 26732 79416 26784
rect 79468 26772 79474 26784
rect 87248 26772 87276 26812
rect 94409 26809 94421 26812
rect 94455 26809 94467 26843
rect 94409 26803 94467 26809
rect 79468 26744 87276 26772
rect 79468 26732 79474 26744
rect 87506 26732 87512 26784
rect 87564 26772 87570 26784
rect 87693 26775 87751 26781
rect 87693 26772 87705 26775
rect 87564 26744 87705 26772
rect 87564 26732 87570 26744
rect 87693 26741 87705 26744
rect 87739 26741 87751 26775
rect 87693 26735 87751 26741
rect 87782 26732 87788 26784
rect 87840 26772 87846 26784
rect 94608 26772 94636 26871
rect 95142 26868 95148 26920
rect 95200 26908 95206 26920
rect 96709 26911 96767 26917
rect 96709 26908 96721 26911
rect 95200 26880 96721 26908
rect 95200 26868 95206 26880
rect 96709 26877 96721 26880
rect 96755 26877 96767 26911
rect 96890 26908 96896 26920
rect 96851 26880 96896 26908
rect 96709 26871 96767 26877
rect 96890 26868 96896 26880
rect 96948 26868 96954 26920
rect 97092 26917 97120 26948
rect 97353 26945 97365 26979
rect 97399 26945 97411 26979
rect 97353 26939 97411 26945
rect 97077 26911 97135 26917
rect 97077 26877 97089 26911
rect 97123 26877 97135 26911
rect 97442 26908 97448 26920
rect 97403 26880 97448 26908
rect 97077 26871 97135 26877
rect 97442 26868 97448 26880
rect 97500 26868 97506 26920
rect 87840 26744 94636 26772
rect 87840 26732 87846 26744
rect 97810 26732 97816 26784
rect 97868 26772 97874 26784
rect 97905 26775 97963 26781
rect 97905 26772 97917 26775
rect 97868 26744 97917 26772
rect 97868 26732 97874 26744
rect 97905 26741 97917 26744
rect 97951 26741 97963 26775
rect 97905 26735 97963 26741
rect 1104 26682 98808 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 50326 26682
rect 50378 26630 50390 26682
rect 50442 26630 50454 26682
rect 50506 26630 50518 26682
rect 50570 26630 81046 26682
rect 81098 26630 81110 26682
rect 81162 26630 81174 26682
rect 81226 26630 81238 26682
rect 81290 26630 98808 26682
rect 1104 26608 98808 26630
rect 5350 26568 5356 26580
rect 5311 26540 5356 26568
rect 5350 26528 5356 26540
rect 5408 26528 5414 26580
rect 13538 26528 13544 26580
rect 13596 26568 13602 26580
rect 16669 26571 16727 26577
rect 16669 26568 16681 26571
rect 13596 26540 16681 26568
rect 13596 26528 13602 26540
rect 16669 26537 16681 26540
rect 16715 26568 16727 26571
rect 19429 26571 19487 26577
rect 19429 26568 19441 26571
rect 16715 26540 19441 26568
rect 16715 26537 16727 26540
rect 16669 26531 16727 26537
rect 19429 26537 19441 26540
rect 19475 26537 19487 26571
rect 19429 26531 19487 26537
rect 21542 26528 21548 26580
rect 21600 26568 21606 26580
rect 30374 26568 30380 26580
rect 21600 26540 30380 26568
rect 21600 26528 21606 26540
rect 30374 26528 30380 26540
rect 30432 26528 30438 26580
rect 30558 26568 30564 26580
rect 30519 26540 30564 26568
rect 30558 26528 30564 26540
rect 30616 26528 30622 26580
rect 30834 26528 30840 26580
rect 30892 26568 30898 26580
rect 33410 26568 33416 26580
rect 30892 26540 33416 26568
rect 30892 26528 30898 26540
rect 33410 26528 33416 26540
rect 33468 26528 33474 26580
rect 35250 26528 35256 26580
rect 35308 26568 35314 26580
rect 35437 26571 35495 26577
rect 35437 26568 35449 26571
rect 35308 26540 35449 26568
rect 35308 26528 35314 26540
rect 35437 26537 35449 26540
rect 35483 26568 35495 26571
rect 35529 26571 35587 26577
rect 35529 26568 35541 26571
rect 35483 26540 35541 26568
rect 35483 26537 35495 26540
rect 35437 26531 35495 26537
rect 35529 26537 35541 26540
rect 35575 26537 35587 26571
rect 35529 26531 35587 26537
rect 36357 26571 36415 26577
rect 36357 26537 36369 26571
rect 36403 26568 36415 26571
rect 37090 26568 37096 26580
rect 36403 26540 37096 26568
rect 36403 26537 36415 26540
rect 36357 26531 36415 26537
rect 37090 26528 37096 26540
rect 37148 26528 37154 26580
rect 37182 26528 37188 26580
rect 37240 26568 37246 26580
rect 40954 26568 40960 26580
rect 37240 26540 40960 26568
rect 37240 26528 37246 26540
rect 40954 26528 40960 26540
rect 41012 26528 41018 26580
rect 41506 26528 41512 26580
rect 41564 26568 41570 26580
rect 87506 26568 87512 26580
rect 41564 26540 87512 26568
rect 41564 26528 41570 26540
rect 87506 26528 87512 26540
rect 87564 26528 87570 26580
rect 90450 26568 90456 26580
rect 90411 26540 90456 26568
rect 90450 26528 90456 26540
rect 90508 26568 90514 26580
rect 90508 26540 91324 26568
rect 90508 26528 90514 26540
rect 10318 26500 10324 26512
rect 5276 26472 10324 26500
rect 4706 26432 4712 26444
rect 4667 26404 4712 26432
rect 4706 26392 4712 26404
rect 4764 26392 4770 26444
rect 4892 26435 4950 26441
rect 4892 26401 4904 26435
rect 4938 26401 4950 26435
rect 4892 26395 4950 26401
rect 4992 26435 5050 26441
rect 4992 26401 5004 26435
rect 5038 26432 5050 26435
rect 5166 26432 5172 26444
rect 5038 26404 5172 26432
rect 5038 26401 5050 26404
rect 4992 26395 5050 26401
rect 4614 26296 4620 26308
rect 4527 26268 4620 26296
rect 4614 26256 4620 26268
rect 4672 26296 4678 26308
rect 4908 26296 4936 26395
rect 5166 26392 5172 26404
rect 5224 26392 5230 26444
rect 5276 26441 5304 26472
rect 10318 26460 10324 26472
rect 10376 26460 10382 26512
rect 20625 26503 20683 26509
rect 20625 26500 20637 26503
rect 19306 26472 20637 26500
rect 5261 26435 5319 26441
rect 5261 26401 5273 26435
rect 5307 26401 5319 26435
rect 5261 26395 5319 26401
rect 6641 26435 6699 26441
rect 6641 26401 6653 26435
rect 6687 26432 6699 26435
rect 6730 26432 6736 26444
rect 6687 26404 6736 26432
rect 6687 26401 6699 26404
rect 6641 26395 6699 26401
rect 6730 26392 6736 26404
rect 6788 26432 6794 26444
rect 6917 26435 6975 26441
rect 6917 26432 6929 26435
rect 6788 26404 6929 26432
rect 6788 26392 6794 26404
rect 6917 26401 6929 26404
rect 6963 26401 6975 26435
rect 6917 26395 6975 26401
rect 13998 26392 14004 26444
rect 14056 26432 14062 26444
rect 15381 26435 15439 26441
rect 14056 26404 15240 26432
rect 14056 26392 14062 26404
rect 5074 26324 5080 26376
rect 5132 26364 5138 26376
rect 15102 26364 15108 26376
rect 5132 26336 5177 26364
rect 15063 26336 15108 26364
rect 5132 26324 5138 26336
rect 15102 26324 15108 26336
rect 15160 26324 15166 26376
rect 15212 26364 15240 26404
rect 15381 26401 15393 26435
rect 15427 26432 15439 26435
rect 19058 26432 19064 26444
rect 15427 26404 19064 26432
rect 15427 26401 15439 26404
rect 15381 26395 15439 26401
rect 19058 26392 19064 26404
rect 19116 26392 19122 26444
rect 19306 26364 19334 26472
rect 20625 26469 20637 26472
rect 20671 26500 20683 26503
rect 20714 26500 20720 26512
rect 20671 26472 20720 26500
rect 20671 26469 20683 26472
rect 20625 26463 20683 26469
rect 20714 26460 20720 26472
rect 20772 26460 20778 26512
rect 21634 26460 21640 26512
rect 21692 26500 21698 26512
rect 33686 26500 33692 26512
rect 21692 26472 33692 26500
rect 21692 26460 21698 26472
rect 33686 26460 33692 26472
rect 33744 26460 33750 26512
rect 36722 26460 36728 26512
rect 36780 26500 36786 26512
rect 40494 26500 40500 26512
rect 36780 26472 40500 26500
rect 36780 26460 36786 26472
rect 40494 26460 40500 26472
rect 40552 26460 40558 26512
rect 46658 26460 46664 26512
rect 46716 26500 46722 26512
rect 46716 26472 49188 26500
rect 46716 26460 46722 26472
rect 20073 26435 20131 26441
rect 20073 26401 20085 26435
rect 20119 26432 20131 26435
rect 21082 26432 21088 26444
rect 20119 26404 21088 26432
rect 20119 26401 20131 26404
rect 20073 26395 20131 26401
rect 21082 26392 21088 26404
rect 21140 26392 21146 26444
rect 21266 26392 21272 26444
rect 21324 26432 21330 26444
rect 21324 26404 21680 26432
rect 21324 26392 21330 26404
rect 15212 26336 19334 26364
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26364 19487 26367
rect 21652 26364 21680 26404
rect 21910 26392 21916 26444
rect 21968 26432 21974 26444
rect 26326 26432 26332 26444
rect 21968 26404 26332 26432
rect 21968 26392 21974 26404
rect 26326 26392 26332 26404
rect 26384 26392 26390 26444
rect 26878 26392 26884 26444
rect 26936 26432 26942 26444
rect 27154 26432 27160 26444
rect 26936 26404 27160 26432
rect 26936 26392 26942 26404
rect 27154 26392 27160 26404
rect 27212 26392 27218 26444
rect 30377 26435 30435 26441
rect 30377 26401 30389 26435
rect 30423 26432 30435 26435
rect 30466 26432 30472 26444
rect 30423 26404 30472 26432
rect 30423 26401 30435 26404
rect 30377 26395 30435 26401
rect 30466 26392 30472 26404
rect 30524 26392 30530 26444
rect 30650 26392 30656 26444
rect 30708 26432 30714 26444
rect 30745 26435 30803 26441
rect 30745 26432 30757 26435
rect 30708 26404 30757 26432
rect 30708 26392 30714 26404
rect 30745 26401 30757 26404
rect 30791 26401 30803 26435
rect 30926 26432 30932 26444
rect 30887 26404 30932 26432
rect 30745 26395 30803 26401
rect 30926 26392 30932 26404
rect 30984 26392 30990 26444
rect 31018 26392 31024 26444
rect 31076 26432 31082 26444
rect 33318 26432 33324 26444
rect 31076 26404 33324 26432
rect 31076 26392 31082 26404
rect 33318 26392 33324 26404
rect 33376 26432 33382 26444
rect 34330 26432 34336 26444
rect 33376 26404 34336 26432
rect 33376 26392 33382 26404
rect 34330 26392 34336 26404
rect 34388 26392 34394 26444
rect 35437 26435 35495 26441
rect 35437 26401 35449 26435
rect 35483 26432 35495 26435
rect 35713 26435 35771 26441
rect 35713 26432 35725 26435
rect 35483 26404 35725 26432
rect 35483 26401 35495 26404
rect 35437 26395 35495 26401
rect 35713 26401 35725 26404
rect 35759 26401 35771 26435
rect 35713 26395 35771 26401
rect 35802 26392 35808 26444
rect 35860 26441 35866 26444
rect 35860 26435 35919 26441
rect 35860 26401 35873 26435
rect 35907 26401 35919 26435
rect 35986 26432 35992 26444
rect 35947 26404 35992 26432
rect 35860 26395 35919 26401
rect 35860 26392 35866 26395
rect 35986 26392 35992 26404
rect 36044 26392 36050 26444
rect 36265 26435 36323 26441
rect 36265 26401 36277 26435
rect 36311 26432 36323 26435
rect 36354 26432 36360 26444
rect 36311 26404 36360 26432
rect 36311 26401 36323 26404
rect 36265 26395 36323 26401
rect 36354 26392 36360 26404
rect 36412 26392 36418 26444
rect 36446 26392 36452 26444
rect 36504 26432 36510 26444
rect 41046 26432 41052 26444
rect 36504 26404 41052 26432
rect 36504 26392 36510 26404
rect 41046 26392 41052 26404
rect 41104 26392 41110 26444
rect 47578 26392 47584 26444
rect 47636 26432 47642 26444
rect 47857 26435 47915 26441
rect 47857 26432 47869 26435
rect 47636 26404 47869 26432
rect 47636 26392 47642 26404
rect 47857 26401 47869 26404
rect 47903 26401 47915 26435
rect 48222 26432 48228 26444
rect 48183 26404 48228 26432
rect 47857 26395 47915 26401
rect 48222 26392 48228 26404
rect 48280 26392 48286 26444
rect 48590 26432 48596 26444
rect 48551 26404 48596 26432
rect 48590 26392 48596 26404
rect 48648 26392 48654 26444
rect 33686 26364 33692 26376
rect 19475 26336 21404 26364
rect 21652 26336 33692 26364
rect 19475 26333 19487 26336
rect 19429 26327 19487 26333
rect 13446 26296 13452 26308
rect 4672 26268 13452 26296
rect 4672 26256 4678 26268
rect 13446 26256 13452 26268
rect 13504 26256 13510 26308
rect 16408 26268 16620 26296
rect 11514 26188 11520 26240
rect 11572 26228 11578 26240
rect 16408 26228 16436 26268
rect 11572 26200 16436 26228
rect 16592 26228 16620 26268
rect 17586 26256 17592 26308
rect 17644 26296 17650 26308
rect 21266 26296 21272 26308
rect 17644 26268 21272 26296
rect 17644 26256 17650 26268
rect 21266 26256 21272 26268
rect 21324 26256 21330 26308
rect 21376 26296 21404 26336
rect 33686 26324 33692 26336
rect 33744 26324 33750 26376
rect 36078 26364 36084 26376
rect 36039 26336 36084 26364
rect 36078 26324 36084 26336
rect 36136 26324 36142 26376
rect 36722 26324 36728 26376
rect 36780 26364 36786 26376
rect 42886 26364 42892 26376
rect 36780 26336 42892 26364
rect 36780 26324 36786 26336
rect 42886 26324 42892 26336
rect 42944 26324 42950 26376
rect 45370 26324 45376 26376
rect 45428 26364 45434 26376
rect 45830 26364 45836 26376
rect 45428 26336 45836 26364
rect 45428 26324 45434 26336
rect 45830 26324 45836 26336
rect 45888 26324 45894 26376
rect 48038 26364 48044 26376
rect 47999 26336 48044 26364
rect 48038 26324 48044 26336
rect 48096 26324 48102 26376
rect 48314 26324 48320 26376
rect 48372 26364 48378 26376
rect 48501 26367 48559 26373
rect 48501 26364 48513 26367
rect 48372 26336 48513 26364
rect 48372 26324 48378 26336
rect 48501 26333 48513 26336
rect 48547 26333 48559 26367
rect 49160 26364 49188 26472
rect 50062 26460 50068 26512
rect 50120 26500 50126 26512
rect 50157 26503 50215 26509
rect 50157 26500 50169 26503
rect 50120 26472 50169 26500
rect 50120 26460 50126 26472
rect 50157 26469 50169 26472
rect 50203 26469 50215 26503
rect 60550 26500 60556 26512
rect 50157 26463 50215 26469
rect 50264 26472 60556 26500
rect 50264 26444 50292 26472
rect 60550 26460 60556 26472
rect 60608 26460 60614 26512
rect 60642 26460 60648 26512
rect 60700 26500 60706 26512
rect 87782 26500 87788 26512
rect 60700 26472 87788 26500
rect 60700 26460 60706 26472
rect 87782 26460 87788 26472
rect 87840 26460 87846 26512
rect 49878 26392 49884 26444
rect 49936 26432 49942 26444
rect 49973 26435 50031 26441
rect 49973 26432 49985 26435
rect 49936 26404 49985 26432
rect 49936 26392 49942 26404
rect 49973 26401 49985 26404
rect 50019 26401 50031 26435
rect 50246 26432 50252 26444
rect 50207 26404 50252 26432
rect 49973 26395 50031 26401
rect 50246 26392 50252 26404
rect 50304 26392 50310 26444
rect 50338 26392 50344 26444
rect 50396 26432 50402 26444
rect 52546 26432 52552 26444
rect 50396 26404 52552 26432
rect 50396 26392 50402 26404
rect 52546 26392 52552 26404
rect 52604 26392 52610 26444
rect 53834 26392 53840 26444
rect 53892 26432 53898 26444
rect 57882 26432 57888 26444
rect 53892 26404 57888 26432
rect 53892 26392 53898 26404
rect 57882 26392 57888 26404
rect 57940 26432 57946 26444
rect 59262 26432 59268 26444
rect 57940 26404 59268 26432
rect 57940 26392 57946 26404
rect 59262 26392 59268 26404
rect 59320 26392 59326 26444
rect 59446 26392 59452 26444
rect 59504 26432 59510 26444
rect 60274 26432 60280 26444
rect 59504 26404 60280 26432
rect 59504 26392 59510 26404
rect 60274 26392 60280 26404
rect 60332 26392 60338 26444
rect 60366 26392 60372 26444
rect 60424 26432 60430 26444
rect 64598 26432 64604 26444
rect 60424 26404 64604 26432
rect 60424 26392 60430 26404
rect 64598 26392 64604 26404
rect 64656 26392 64662 26444
rect 64690 26392 64696 26444
rect 64748 26432 64754 26444
rect 70578 26432 70584 26444
rect 64748 26404 70584 26432
rect 64748 26392 64754 26404
rect 70578 26392 70584 26404
rect 70636 26392 70642 26444
rect 72878 26392 72884 26444
rect 72936 26432 72942 26444
rect 73798 26441 73804 26444
rect 73341 26435 73399 26441
rect 73341 26432 73353 26435
rect 72936 26404 73353 26432
rect 72936 26392 72942 26404
rect 73341 26401 73353 26404
rect 73387 26401 73399 26435
rect 73506 26435 73564 26441
rect 73506 26432 73518 26435
rect 73341 26395 73399 26401
rect 73448 26404 73518 26432
rect 72510 26364 72516 26376
rect 49160 26336 72516 26364
rect 48501 26327 48559 26333
rect 72510 26324 72516 26336
rect 72568 26324 72574 26376
rect 48682 26296 48688 26308
rect 21376 26268 48688 26296
rect 48682 26256 48688 26268
rect 48740 26256 48746 26308
rect 48866 26256 48872 26308
rect 48924 26296 48930 26308
rect 48961 26299 49019 26305
rect 48961 26296 48973 26299
rect 48924 26268 48973 26296
rect 48924 26256 48930 26268
rect 48961 26265 48973 26268
rect 49007 26265 49019 26299
rect 48961 26259 49019 26265
rect 53098 26256 53104 26308
rect 53156 26296 53162 26308
rect 60366 26296 60372 26308
rect 53156 26268 60372 26296
rect 53156 26256 53162 26268
rect 60366 26256 60372 26268
rect 60424 26256 60430 26308
rect 60458 26256 60464 26308
rect 60516 26296 60522 26308
rect 64690 26296 64696 26308
rect 60516 26268 64696 26296
rect 60516 26256 60522 26268
rect 64690 26256 64696 26268
rect 64748 26256 64754 26308
rect 73338 26256 73344 26308
rect 73396 26296 73402 26308
rect 73448 26296 73476 26404
rect 73506 26401 73518 26404
rect 73552 26401 73564 26435
rect 73506 26395 73564 26401
rect 73755 26435 73804 26441
rect 73755 26401 73767 26435
rect 73801 26401 73804 26435
rect 73755 26395 73804 26401
rect 73798 26392 73804 26395
rect 73856 26392 73862 26444
rect 73893 26435 73951 26441
rect 73893 26401 73905 26435
rect 73939 26401 73951 26435
rect 74074 26432 74080 26444
rect 74035 26404 74080 26432
rect 73893 26395 73951 26401
rect 73614 26364 73620 26376
rect 73575 26336 73620 26364
rect 73614 26324 73620 26336
rect 73672 26324 73678 26376
rect 73908 26364 73936 26395
rect 74074 26392 74080 26404
rect 74132 26392 74138 26444
rect 75086 26392 75092 26444
rect 75144 26432 75150 26444
rect 86037 26435 86095 26441
rect 86037 26432 86049 26435
rect 75144 26404 86049 26432
rect 75144 26392 75150 26404
rect 86037 26401 86049 26404
rect 86083 26432 86095 26435
rect 86310 26432 86316 26444
rect 86083 26404 86316 26432
rect 86083 26401 86095 26404
rect 86037 26395 86095 26401
rect 86310 26392 86316 26404
rect 86368 26432 86374 26444
rect 86402 26432 86408 26444
rect 86368 26404 86408 26432
rect 86368 26392 86374 26404
rect 86402 26392 86408 26404
rect 86460 26392 86466 26444
rect 86543 26435 86601 26441
rect 86543 26401 86555 26435
rect 86589 26401 86601 26435
rect 86678 26432 86684 26444
rect 86639 26404 86684 26432
rect 86543 26395 86601 26401
rect 73982 26364 73988 26376
rect 73908 26336 73988 26364
rect 73982 26324 73988 26336
rect 74040 26324 74046 26376
rect 74350 26324 74356 26376
rect 74408 26364 74414 26376
rect 86126 26364 86132 26376
rect 74408 26336 86132 26364
rect 74408 26324 74414 26336
rect 86126 26324 86132 26336
rect 86184 26324 86190 26376
rect 73396 26268 73476 26296
rect 73396 26256 73402 26268
rect 74626 26256 74632 26308
rect 74684 26296 74690 26308
rect 83550 26296 83556 26308
rect 74684 26268 83556 26296
rect 74684 26256 74690 26268
rect 83550 26256 83556 26268
rect 83608 26256 83614 26308
rect 83642 26256 83648 26308
rect 83700 26296 83706 26308
rect 86221 26299 86279 26305
rect 83700 26268 85574 26296
rect 83700 26256 83706 26268
rect 43254 26228 43260 26240
rect 16592 26200 43260 26228
rect 11572 26188 11578 26200
rect 43254 26188 43260 26200
rect 43312 26188 43318 26240
rect 43346 26188 43352 26240
rect 43404 26228 43410 26240
rect 49878 26228 49884 26240
rect 43404 26200 49884 26228
rect 43404 26188 43410 26200
rect 49878 26188 49884 26200
rect 49936 26188 49942 26240
rect 50062 26188 50068 26240
rect 50120 26228 50126 26240
rect 50525 26231 50583 26237
rect 50525 26228 50537 26231
rect 50120 26200 50537 26228
rect 50120 26188 50126 26200
rect 50525 26197 50537 26200
rect 50571 26197 50583 26231
rect 50525 26191 50583 26197
rect 52822 26188 52828 26240
rect 52880 26228 52886 26240
rect 60182 26228 60188 26240
rect 52880 26200 60188 26228
rect 52880 26188 52886 26200
rect 60182 26188 60188 26200
rect 60240 26188 60246 26240
rect 61286 26188 61292 26240
rect 61344 26228 61350 26240
rect 63494 26228 63500 26240
rect 61344 26200 63500 26228
rect 61344 26188 61350 26200
rect 63494 26188 63500 26200
rect 63552 26188 63558 26240
rect 65426 26188 65432 26240
rect 65484 26228 65490 26240
rect 73430 26228 73436 26240
rect 65484 26200 73436 26228
rect 65484 26188 65490 26200
rect 73430 26188 73436 26200
rect 73488 26188 73494 26240
rect 74258 26188 74264 26240
rect 74316 26228 74322 26240
rect 81802 26228 81808 26240
rect 74316 26200 81808 26228
rect 74316 26188 74322 26200
rect 81802 26188 81808 26200
rect 81860 26188 81866 26240
rect 85546 26228 85574 26268
rect 86221 26265 86233 26299
rect 86267 26296 86279 26299
rect 86310 26296 86316 26308
rect 86267 26268 86316 26296
rect 86267 26265 86279 26268
rect 86221 26259 86279 26265
rect 86310 26256 86316 26268
rect 86368 26256 86374 26308
rect 86558 26228 86586 26395
rect 86678 26392 86684 26404
rect 86736 26392 86742 26444
rect 86862 26441 86868 26444
rect 86809 26435 86868 26441
rect 86809 26401 86821 26435
rect 86855 26401 86868 26435
rect 86809 26395 86868 26401
rect 86862 26392 86868 26395
rect 86920 26392 86926 26444
rect 86957 26435 87015 26441
rect 86957 26401 86969 26435
rect 87003 26432 87015 26435
rect 87046 26432 87052 26444
rect 87003 26404 87052 26432
rect 87003 26401 87015 26404
rect 86957 26395 87015 26401
rect 87046 26392 87052 26404
rect 87104 26392 87110 26444
rect 91296 26441 91324 26540
rect 91281 26435 91339 26441
rect 91281 26401 91293 26435
rect 91327 26401 91339 26435
rect 91646 26432 91652 26444
rect 91607 26404 91652 26432
rect 91281 26395 91339 26401
rect 91646 26392 91652 26404
rect 91704 26392 91710 26444
rect 91830 26432 91836 26444
rect 91791 26404 91836 26432
rect 91830 26392 91836 26404
rect 91888 26392 91894 26444
rect 87966 26364 87972 26376
rect 87927 26336 87972 26364
rect 87966 26324 87972 26336
rect 88024 26364 88030 26376
rect 88153 26367 88211 26373
rect 88153 26364 88165 26367
rect 88024 26336 88165 26364
rect 88024 26324 88030 26336
rect 88153 26333 88165 26336
rect 88199 26333 88211 26367
rect 88153 26327 88211 26333
rect 88242 26324 88248 26376
rect 88300 26364 88306 26376
rect 90637 26367 90695 26373
rect 90637 26364 90649 26367
rect 88300 26336 90649 26364
rect 88300 26324 88306 26336
rect 90637 26333 90649 26336
rect 90683 26333 90695 26367
rect 90637 26327 90695 26333
rect 91373 26367 91431 26373
rect 91373 26333 91385 26367
rect 91419 26333 91431 26367
rect 91373 26327 91431 26333
rect 91388 26296 91416 26327
rect 91554 26324 91560 26376
rect 91612 26364 91618 26376
rect 91848 26364 91876 26392
rect 91612 26336 91876 26364
rect 91612 26324 91618 26336
rect 91922 26296 91928 26308
rect 91388 26268 91928 26296
rect 91922 26256 91928 26268
rect 91980 26256 91986 26308
rect 85546 26200 86586 26228
rect 1104 26138 98808 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 65686 26138
rect 65738 26086 65750 26138
rect 65802 26086 65814 26138
rect 65866 26086 65878 26138
rect 65930 26086 96406 26138
rect 96458 26086 96470 26138
rect 96522 26086 96534 26138
rect 96586 26086 96598 26138
rect 96650 26086 98808 26138
rect 1104 26064 98808 26086
rect 11698 25984 11704 26036
rect 11756 26024 11762 26036
rect 11756 25996 20208 26024
rect 11756 25984 11762 25996
rect 15102 25916 15108 25968
rect 15160 25956 15166 25968
rect 15930 25956 15936 25968
rect 15160 25928 15936 25956
rect 15160 25916 15166 25928
rect 15930 25916 15936 25928
rect 15988 25916 15994 25968
rect 20180 25956 20208 25996
rect 20346 25984 20352 26036
rect 20404 26024 20410 26036
rect 26878 26024 26884 26036
rect 20404 25996 26884 26024
rect 20404 25984 20410 25996
rect 26878 25984 26884 25996
rect 26936 25984 26942 26036
rect 41414 26024 41420 26036
rect 31726 25996 41420 26024
rect 31726 25956 31754 25996
rect 41414 25984 41420 25996
rect 41472 25984 41478 26036
rect 41506 25984 41512 26036
rect 41564 26024 41570 26036
rect 41564 25996 53419 26024
rect 41564 25984 41570 25996
rect 20180 25928 31754 25956
rect 31846 25916 31852 25968
rect 31904 25956 31910 25968
rect 36998 25956 37004 25968
rect 31904 25928 37004 25956
rect 31904 25916 31910 25928
rect 36998 25916 37004 25928
rect 37056 25916 37062 25968
rect 37458 25916 37464 25968
rect 37516 25956 37522 25968
rect 38194 25956 38200 25968
rect 37516 25928 38200 25956
rect 37516 25916 37522 25928
rect 38194 25916 38200 25928
rect 38252 25916 38258 25968
rect 38286 25916 38292 25968
rect 38344 25956 38350 25968
rect 45554 25956 45560 25968
rect 38344 25928 45560 25956
rect 38344 25916 38350 25928
rect 45554 25916 45560 25928
rect 45612 25916 45618 25968
rect 45646 25916 45652 25968
rect 45704 25956 45710 25968
rect 50430 25956 50436 25968
rect 45704 25928 50436 25956
rect 45704 25916 45710 25928
rect 50430 25916 50436 25928
rect 50488 25916 50494 25968
rect 53391 25956 53419 25996
rect 53742 25984 53748 26036
rect 53800 26024 53806 26036
rect 65426 26024 65432 26036
rect 53800 25996 65432 26024
rect 53800 25984 53806 25996
rect 65426 25984 65432 25996
rect 65484 25984 65490 26036
rect 77478 26024 77484 26036
rect 65536 25996 77484 26024
rect 65536 25956 65564 25996
rect 77478 25984 77484 25996
rect 77536 25984 77542 26036
rect 53391 25928 65564 25956
rect 68741 25959 68799 25965
rect 68741 25925 68753 25959
rect 68787 25956 68799 25959
rect 69106 25956 69112 25968
rect 68787 25928 69112 25956
rect 68787 25925 68799 25928
rect 68741 25919 68799 25925
rect 69106 25916 69112 25928
rect 69164 25916 69170 25968
rect 73430 25916 73436 25968
rect 73488 25956 73494 25968
rect 75914 25956 75920 25968
rect 73488 25928 75920 25956
rect 73488 25916 73494 25928
rect 75914 25916 75920 25928
rect 75972 25956 75978 25968
rect 91554 25956 91560 25968
rect 75972 25928 91560 25956
rect 75972 25916 75978 25928
rect 91554 25916 91560 25928
rect 91612 25916 91618 25968
rect 17218 25848 17224 25900
rect 17276 25888 17282 25900
rect 17276 25860 19196 25888
rect 17276 25848 17282 25860
rect 18874 25780 18880 25832
rect 18932 25820 18938 25832
rect 19058 25820 19064 25832
rect 18932 25792 19064 25820
rect 18932 25780 18938 25792
rect 19058 25780 19064 25792
rect 19116 25780 19122 25832
rect 19168 25820 19196 25860
rect 20456 25860 23796 25888
rect 20346 25820 20352 25832
rect 19168 25792 20352 25820
rect 20346 25780 20352 25792
rect 20404 25780 20410 25832
rect 19328 25755 19386 25761
rect 19328 25721 19340 25755
rect 19374 25752 19386 25755
rect 19886 25752 19892 25764
rect 19374 25724 19892 25752
rect 19374 25721 19386 25724
rect 19328 25715 19386 25721
rect 19886 25712 19892 25724
rect 19944 25712 19950 25764
rect 20456 25752 20484 25860
rect 22922 25820 22928 25832
rect 22883 25792 22928 25820
rect 22922 25780 22928 25792
rect 22980 25780 22986 25832
rect 23768 25820 23796 25860
rect 24486 25848 24492 25900
rect 24544 25888 24550 25900
rect 24544 25860 53144 25888
rect 24544 25848 24550 25860
rect 23768 25792 39160 25820
rect 20180 25724 20484 25752
rect 15470 25644 15476 25696
rect 15528 25684 15534 25696
rect 20180 25684 20208 25724
rect 20898 25712 20904 25764
rect 20956 25752 20962 25764
rect 39132 25752 39160 25792
rect 39206 25780 39212 25832
rect 39264 25829 39270 25832
rect 39264 25820 39274 25829
rect 39390 25820 39396 25832
rect 39264 25792 39309 25820
rect 39351 25792 39396 25820
rect 39264 25783 39274 25792
rect 39264 25780 39270 25783
rect 39390 25780 39396 25792
rect 39448 25780 39454 25832
rect 39574 25780 39580 25832
rect 39632 25820 39638 25832
rect 39850 25820 39856 25832
rect 39632 25792 39677 25820
rect 39811 25792 39856 25820
rect 39632 25780 39638 25792
rect 39850 25780 39856 25792
rect 39908 25780 39914 25832
rect 39945 25823 40003 25829
rect 39945 25789 39957 25823
rect 39991 25820 40003 25823
rect 39991 25792 43484 25820
rect 39991 25789 40003 25792
rect 39945 25783 40003 25789
rect 39960 25752 39988 25783
rect 43346 25752 43352 25764
rect 20956 25724 39068 25752
rect 39132 25724 39988 25752
rect 40052 25724 43352 25752
rect 20956 25712 20962 25724
rect 15528 25656 20208 25684
rect 15528 25644 15534 25656
rect 20254 25644 20260 25696
rect 20312 25684 20318 25696
rect 20441 25687 20499 25693
rect 20441 25684 20453 25687
rect 20312 25656 20453 25684
rect 20312 25644 20318 25656
rect 20441 25653 20453 25656
rect 20487 25653 20499 25687
rect 20441 25647 20499 25653
rect 26878 25644 26884 25696
rect 26936 25684 26942 25696
rect 34606 25684 34612 25696
rect 26936 25656 34612 25684
rect 26936 25644 26942 25656
rect 34606 25644 34612 25656
rect 34664 25684 34670 25696
rect 35802 25684 35808 25696
rect 34664 25656 35808 25684
rect 34664 25644 34670 25656
rect 35802 25644 35808 25656
rect 35860 25644 35866 25696
rect 35986 25644 35992 25696
rect 36044 25684 36050 25696
rect 38010 25684 38016 25696
rect 36044 25656 38016 25684
rect 36044 25644 36050 25656
rect 38010 25644 38016 25656
rect 38068 25644 38074 25696
rect 39040 25684 39068 25724
rect 39574 25684 39580 25696
rect 39040 25656 39580 25684
rect 39574 25644 39580 25656
rect 39632 25684 39638 25696
rect 40052 25684 40080 25724
rect 43346 25712 43352 25724
rect 43404 25712 43410 25764
rect 43456 25752 43484 25792
rect 43530 25780 43536 25832
rect 43588 25820 43594 25832
rect 52822 25820 52828 25832
rect 43588 25792 52828 25820
rect 43588 25780 43594 25792
rect 52822 25780 52828 25792
rect 52880 25780 52886 25832
rect 49786 25752 49792 25764
rect 43456 25724 49792 25752
rect 49786 25712 49792 25724
rect 49844 25712 49850 25764
rect 50430 25712 50436 25764
rect 50488 25752 50494 25764
rect 52362 25752 52368 25764
rect 50488 25724 52368 25752
rect 50488 25712 50494 25724
rect 52362 25712 52368 25724
rect 52420 25712 52426 25764
rect 53116 25752 53144 25860
rect 56226 25848 56232 25900
rect 56284 25888 56290 25900
rect 65426 25888 65432 25900
rect 56284 25860 65432 25888
rect 56284 25848 56290 25860
rect 65426 25848 65432 25860
rect 65484 25848 65490 25900
rect 86586 25888 86592 25900
rect 65536 25860 86592 25888
rect 56042 25780 56048 25832
rect 56100 25820 56106 25832
rect 61194 25820 61200 25832
rect 56100 25792 61200 25820
rect 56100 25780 56106 25792
rect 61194 25780 61200 25792
rect 61252 25780 61258 25832
rect 61654 25820 61660 25832
rect 61615 25792 61660 25820
rect 61654 25780 61660 25792
rect 61712 25780 61718 25832
rect 61746 25780 61752 25832
rect 61804 25820 61810 25832
rect 65242 25820 65248 25832
rect 61804 25792 65248 25820
rect 61804 25780 61810 25792
rect 65242 25780 65248 25792
rect 65300 25780 65306 25832
rect 65536 25752 65564 25860
rect 86586 25848 86592 25860
rect 86644 25888 86650 25900
rect 87414 25888 87420 25900
rect 86644 25860 87420 25888
rect 86644 25848 86650 25860
rect 87414 25848 87420 25860
rect 87472 25848 87478 25900
rect 66346 25820 66352 25832
rect 66307 25792 66352 25820
rect 66346 25780 66352 25792
rect 66404 25780 66410 25832
rect 67174 25820 67180 25832
rect 67135 25792 67180 25820
rect 67174 25780 67180 25792
rect 67232 25780 67238 25832
rect 67453 25823 67511 25829
rect 67453 25789 67465 25823
rect 67499 25820 67511 25823
rect 67542 25820 67548 25832
rect 67499 25792 67548 25820
rect 67499 25789 67511 25792
rect 67453 25783 67511 25789
rect 67542 25780 67548 25792
rect 67600 25780 67606 25832
rect 73246 25780 73252 25832
rect 73304 25820 73310 25832
rect 73982 25820 73988 25832
rect 73304 25792 73988 25820
rect 73304 25780 73310 25792
rect 73982 25780 73988 25792
rect 74040 25780 74046 25832
rect 80422 25820 80428 25832
rect 80383 25792 80428 25820
rect 80422 25780 80428 25792
rect 80480 25780 80486 25832
rect 53116 25724 65564 25752
rect 68112 25724 68692 25752
rect 39632 25656 40080 25684
rect 40405 25687 40463 25693
rect 39632 25644 39638 25656
rect 40405 25653 40417 25687
rect 40451 25684 40463 25687
rect 68112 25684 68140 25724
rect 40451 25656 68140 25684
rect 68664 25684 68692 25724
rect 70118 25712 70124 25764
rect 70176 25752 70182 25764
rect 82170 25752 82176 25764
rect 70176 25724 82176 25752
rect 70176 25712 70182 25724
rect 82170 25712 82176 25724
rect 82228 25752 82234 25764
rect 82722 25752 82728 25764
rect 82228 25724 82728 25752
rect 82228 25712 82234 25724
rect 82722 25712 82728 25724
rect 82780 25712 82786 25764
rect 93210 25684 93216 25696
rect 68664 25656 93216 25684
rect 40451 25653 40463 25656
rect 40405 25647 40463 25653
rect 93210 25644 93216 25656
rect 93268 25644 93274 25696
rect 1104 25594 98808 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 50326 25594
rect 50378 25542 50390 25594
rect 50442 25542 50454 25594
rect 50506 25542 50518 25594
rect 50570 25542 81046 25594
rect 81098 25542 81110 25594
rect 81162 25542 81174 25594
rect 81226 25542 81238 25594
rect 81290 25542 98808 25594
rect 1104 25520 98808 25542
rect 15194 25440 15200 25492
rect 15252 25480 15258 25492
rect 20898 25480 20904 25492
rect 15252 25452 20904 25480
rect 15252 25440 15258 25452
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 21637 25483 21695 25489
rect 21637 25449 21649 25483
rect 21683 25480 21695 25483
rect 21818 25480 21824 25492
rect 21683 25452 21824 25480
rect 21683 25449 21695 25452
rect 21637 25443 21695 25449
rect 21818 25440 21824 25452
rect 21876 25440 21882 25492
rect 21910 25440 21916 25492
rect 21968 25480 21974 25492
rect 37366 25480 37372 25492
rect 21968 25452 37372 25480
rect 21968 25440 21974 25452
rect 37366 25440 37372 25452
rect 37424 25440 37430 25492
rect 38562 25440 38568 25492
rect 38620 25480 38626 25492
rect 39390 25480 39396 25492
rect 38620 25452 39396 25480
rect 38620 25440 38626 25452
rect 39390 25440 39396 25452
rect 39448 25440 39454 25492
rect 43533 25483 43591 25489
rect 43533 25480 43545 25483
rect 39500 25452 43545 25480
rect 3050 25372 3056 25424
rect 3108 25412 3114 25424
rect 21174 25412 21180 25424
rect 3108 25384 21180 25412
rect 3108 25372 3114 25384
rect 21174 25372 21180 25384
rect 21232 25372 21238 25424
rect 21836 25412 21864 25440
rect 21836 25384 31754 25412
rect 21545 25347 21603 25353
rect 21545 25313 21557 25347
rect 21591 25344 21603 25347
rect 21726 25344 21732 25356
rect 21591 25316 21732 25344
rect 21591 25313 21603 25316
rect 21545 25307 21603 25313
rect 21726 25304 21732 25316
rect 21784 25304 21790 25356
rect 21821 25347 21879 25353
rect 21821 25313 21833 25347
rect 21867 25344 21879 25347
rect 22094 25344 22100 25356
rect 21867 25316 22100 25344
rect 21867 25313 21879 25316
rect 21821 25307 21879 25313
rect 22094 25304 22100 25316
rect 22152 25344 22158 25356
rect 22462 25344 22468 25356
rect 22152 25316 22468 25344
rect 22152 25304 22158 25316
rect 22462 25304 22468 25316
rect 22520 25304 22526 25356
rect 30926 25344 30932 25356
rect 25792 25316 30932 25344
rect 19886 25236 19892 25288
rect 19944 25276 19950 25288
rect 25792 25276 25820 25316
rect 30926 25304 30932 25316
rect 30984 25304 30990 25356
rect 31726 25344 31754 25384
rect 32122 25372 32128 25424
rect 32180 25412 32186 25424
rect 39500 25412 39528 25452
rect 43533 25449 43545 25452
rect 43579 25449 43591 25483
rect 52086 25480 52092 25492
rect 43533 25443 43591 25449
rect 43640 25452 52092 25480
rect 32180 25384 39528 25412
rect 32180 25372 32186 25384
rect 42334 25372 42340 25424
rect 42392 25412 42398 25424
rect 42610 25412 42616 25424
rect 42392 25384 42616 25412
rect 42392 25372 42398 25384
rect 42610 25372 42616 25384
rect 42668 25372 42674 25424
rect 43640 25412 43668 25452
rect 52086 25440 52092 25452
rect 52144 25440 52150 25492
rect 52365 25483 52423 25489
rect 52365 25449 52377 25483
rect 52411 25480 52423 25483
rect 53190 25480 53196 25492
rect 52411 25452 53196 25480
rect 52411 25449 52423 25452
rect 52365 25443 52423 25449
rect 53190 25440 53196 25452
rect 53248 25440 53254 25492
rect 54570 25440 54576 25492
rect 54628 25480 54634 25492
rect 56318 25480 56324 25492
rect 54628 25452 56324 25480
rect 54628 25440 54634 25452
rect 56318 25440 56324 25452
rect 56376 25440 56382 25492
rect 56502 25440 56508 25492
rect 56560 25480 56566 25492
rect 60734 25480 60740 25492
rect 56560 25452 60740 25480
rect 56560 25440 56566 25452
rect 60734 25440 60740 25452
rect 60792 25480 60798 25492
rect 61378 25480 61384 25492
rect 60792 25452 61384 25480
rect 60792 25440 60798 25452
rect 61378 25440 61384 25452
rect 61436 25440 61442 25492
rect 65242 25440 65248 25492
rect 65300 25480 65306 25492
rect 70118 25480 70124 25492
rect 65300 25452 70124 25480
rect 65300 25440 65306 25452
rect 70118 25440 70124 25452
rect 70176 25440 70182 25492
rect 70210 25440 70216 25492
rect 70268 25480 70274 25492
rect 82354 25480 82360 25492
rect 70268 25452 82360 25480
rect 70268 25440 70274 25452
rect 82354 25440 82360 25452
rect 82412 25480 82418 25492
rect 82412 25452 91416 25480
rect 82412 25440 82418 25452
rect 43272 25384 43668 25412
rect 38654 25344 38660 25356
rect 31726 25316 38660 25344
rect 38654 25304 38660 25316
rect 38712 25344 38718 25356
rect 40494 25344 40500 25356
rect 38712 25316 40500 25344
rect 38712 25304 38718 25316
rect 40494 25304 40500 25316
rect 40552 25304 40558 25356
rect 41233 25347 41291 25353
rect 40880 25316 41092 25344
rect 19944 25248 25820 25276
rect 19944 25236 19950 25248
rect 25866 25236 25872 25288
rect 25924 25276 25930 25288
rect 39022 25276 39028 25288
rect 25924 25248 39028 25276
rect 25924 25236 25930 25248
rect 39022 25236 39028 25248
rect 39080 25276 39086 25288
rect 40880 25276 40908 25316
rect 39080 25248 40908 25276
rect 40957 25279 41015 25285
rect 39080 25236 39086 25248
rect 40957 25245 40969 25279
rect 41003 25245 41015 25279
rect 41064 25276 41092 25316
rect 41233 25313 41245 25347
rect 41279 25344 41291 25347
rect 41322 25344 41328 25356
rect 41279 25316 41328 25344
rect 41279 25313 41291 25316
rect 41233 25307 41291 25313
rect 41322 25304 41328 25316
rect 41380 25304 41386 25356
rect 41506 25304 41512 25356
rect 41564 25344 41570 25356
rect 41874 25344 41880 25356
rect 41564 25316 41880 25344
rect 41564 25304 41570 25316
rect 41874 25304 41880 25316
rect 41932 25304 41938 25356
rect 43272 25276 43300 25384
rect 43714 25372 43720 25424
rect 43772 25412 43778 25424
rect 43772 25384 47532 25412
rect 43772 25372 43778 25384
rect 43622 25344 43628 25356
rect 43583 25316 43628 25344
rect 43622 25304 43628 25316
rect 43680 25304 43686 25356
rect 44082 25353 44088 25356
rect 43901 25347 43959 25353
rect 43901 25344 43913 25347
rect 43732 25316 43913 25344
rect 41064 25248 43300 25276
rect 40957 25239 41015 25245
rect 17770 25168 17776 25220
rect 17828 25208 17834 25220
rect 17828 25180 27844 25208
rect 17828 25168 17834 25180
rect 15194 25100 15200 25152
rect 15252 25140 15258 25152
rect 15378 25140 15384 25152
rect 15252 25112 15384 25140
rect 15252 25100 15258 25112
rect 15378 25100 15384 25112
rect 15436 25100 15442 25152
rect 21453 25143 21511 25149
rect 21453 25109 21465 25143
rect 21499 25140 21511 25143
rect 21818 25140 21824 25152
rect 21499 25112 21824 25140
rect 21499 25109 21511 25112
rect 21453 25103 21511 25109
rect 21818 25100 21824 25112
rect 21876 25100 21882 25152
rect 21910 25100 21916 25152
rect 21968 25140 21974 25152
rect 22005 25143 22063 25149
rect 22005 25140 22017 25143
rect 21968 25112 22017 25140
rect 21968 25100 21974 25112
rect 22005 25109 22017 25112
rect 22051 25109 22063 25143
rect 27706 25140 27712 25152
rect 27667 25112 27712 25140
rect 22005 25103 22063 25109
rect 27706 25100 27712 25112
rect 27764 25100 27770 25152
rect 27816 25140 27844 25180
rect 30466 25168 30472 25220
rect 30524 25208 30530 25220
rect 39850 25208 39856 25220
rect 30524 25180 39856 25208
rect 30524 25168 30530 25180
rect 39850 25168 39856 25180
rect 39908 25168 39914 25220
rect 40678 25168 40684 25220
rect 40736 25208 40742 25220
rect 40972 25208 41000 25239
rect 43346 25236 43352 25288
rect 43404 25276 43410 25288
rect 43732 25276 43760 25316
rect 43901 25313 43913 25316
rect 43947 25313 43959 25347
rect 43901 25307 43959 25313
rect 44029 25347 44088 25353
rect 44029 25313 44041 25347
rect 44075 25313 44088 25347
rect 44029 25307 44088 25313
rect 44082 25304 44088 25307
rect 44140 25304 44146 25356
rect 44177 25347 44235 25353
rect 44177 25313 44189 25347
rect 44223 25344 44235 25347
rect 44542 25344 44548 25356
rect 44223 25316 44548 25344
rect 44223 25313 44235 25316
rect 44177 25307 44235 25313
rect 44542 25304 44548 25316
rect 44600 25344 44606 25356
rect 47504 25344 47532 25384
rect 47578 25372 47584 25424
rect 47636 25412 47642 25424
rect 63126 25412 63132 25424
rect 47636 25384 63132 25412
rect 47636 25372 47642 25384
rect 48498 25344 48504 25356
rect 44600 25316 47440 25344
rect 47504 25316 48504 25344
rect 44600 25304 44606 25316
rect 43404 25248 43760 25276
rect 43809 25279 43867 25285
rect 43404 25236 43410 25248
rect 43809 25245 43821 25279
rect 43855 25276 43867 25279
rect 44266 25276 44272 25288
rect 43855 25248 44272 25276
rect 43855 25245 43867 25248
rect 43809 25239 43867 25245
rect 44266 25236 44272 25248
rect 44324 25276 44330 25288
rect 45646 25276 45652 25288
rect 44324 25248 45652 25276
rect 44324 25236 44330 25248
rect 45646 25236 45652 25248
rect 45704 25236 45710 25288
rect 47412 25276 47440 25316
rect 48498 25304 48504 25316
rect 48556 25344 48562 25356
rect 50982 25344 50988 25356
rect 48556 25316 50988 25344
rect 48556 25304 48562 25316
rect 50982 25304 50988 25316
rect 51040 25304 51046 25356
rect 51644 25353 51672 25384
rect 63126 25372 63132 25384
rect 63184 25372 63190 25424
rect 65426 25372 65432 25424
rect 65484 25412 65490 25424
rect 76466 25412 76472 25424
rect 65484 25384 76472 25412
rect 65484 25372 65490 25384
rect 76466 25372 76472 25384
rect 76524 25372 76530 25424
rect 82722 25372 82728 25424
rect 82780 25412 82786 25424
rect 82780 25384 91048 25412
rect 82780 25372 82786 25384
rect 51629 25347 51687 25353
rect 51629 25313 51641 25347
rect 51675 25313 51687 25347
rect 51810 25344 51816 25356
rect 51771 25316 51816 25344
rect 51629 25307 51687 25313
rect 51810 25304 51816 25316
rect 51868 25304 51874 25356
rect 52178 25344 52184 25356
rect 52139 25316 52184 25344
rect 52178 25304 52184 25316
rect 52236 25304 52242 25356
rect 53009 25347 53067 25353
rect 53009 25313 53021 25347
rect 53055 25313 53067 25347
rect 53190 25344 53196 25356
rect 53151 25316 53196 25344
rect 53009 25307 53067 25313
rect 48406 25276 48412 25288
rect 47412 25248 48412 25276
rect 48406 25236 48412 25248
rect 48464 25236 48470 25288
rect 48590 25236 48596 25288
rect 48648 25276 48654 25288
rect 49510 25276 49516 25288
rect 48648 25248 49516 25276
rect 48648 25236 48654 25248
rect 49510 25236 49516 25248
rect 49568 25276 49574 25288
rect 51902 25276 51908 25288
rect 49568 25248 51396 25276
rect 51863 25248 51908 25276
rect 49568 25236 49574 25248
rect 51258 25208 51264 25220
rect 40736 25180 41000 25208
rect 42260 25180 51264 25208
rect 40736 25168 40742 25180
rect 42260 25140 42288 25180
rect 51258 25168 51264 25180
rect 51316 25168 51322 25220
rect 51368 25208 51396 25248
rect 51902 25236 51908 25248
rect 51960 25236 51966 25288
rect 51997 25279 52055 25285
rect 51997 25245 52009 25279
rect 52043 25245 52055 25279
rect 53024 25276 53052 25307
rect 53190 25304 53196 25316
rect 53248 25304 53254 25356
rect 53285 25347 53343 25353
rect 53285 25313 53297 25347
rect 53331 25344 53343 25347
rect 53558 25344 53564 25356
rect 53331 25316 53564 25344
rect 53331 25313 53343 25316
rect 53285 25307 53343 25313
rect 53558 25304 53564 25316
rect 53616 25304 53622 25356
rect 53650 25304 53656 25356
rect 53708 25344 53714 25356
rect 53708 25316 56180 25344
rect 53708 25304 53714 25316
rect 56042 25276 56048 25288
rect 53024 25248 56048 25276
rect 51997 25239 52055 25245
rect 52012 25208 52040 25239
rect 56042 25236 56048 25248
rect 56100 25236 56106 25288
rect 56152 25276 56180 25316
rect 56226 25304 56232 25356
rect 56284 25344 56290 25356
rect 61286 25344 61292 25356
rect 56284 25316 61292 25344
rect 56284 25304 56290 25316
rect 61286 25304 61292 25316
rect 61344 25304 61350 25356
rect 61378 25304 61384 25356
rect 61436 25344 61442 25356
rect 64966 25344 64972 25356
rect 61436 25316 64972 25344
rect 61436 25304 61442 25316
rect 64966 25304 64972 25316
rect 65024 25304 65030 25356
rect 66438 25304 66444 25356
rect 66496 25344 66502 25356
rect 73617 25347 73675 25353
rect 73617 25344 73629 25347
rect 66496 25316 73629 25344
rect 66496 25304 66502 25316
rect 73617 25313 73629 25316
rect 73663 25313 73675 25347
rect 73617 25307 73675 25313
rect 81802 25304 81808 25356
rect 81860 25344 81866 25356
rect 89530 25344 89536 25356
rect 81860 25316 89536 25344
rect 81860 25304 81866 25316
rect 89530 25304 89536 25316
rect 89588 25344 89594 25356
rect 91020 25353 91048 25384
rect 91388 25353 91416 25452
rect 90637 25347 90695 25353
rect 90637 25344 90649 25347
rect 89588 25316 90649 25344
rect 89588 25304 89594 25316
rect 90637 25313 90649 25316
rect 90683 25313 90695 25347
rect 90637 25307 90695 25313
rect 91005 25347 91063 25353
rect 91005 25313 91017 25347
rect 91051 25313 91063 25347
rect 91005 25307 91063 25313
rect 91373 25347 91431 25353
rect 91373 25313 91385 25347
rect 91419 25313 91431 25347
rect 91373 25307 91431 25313
rect 74350 25276 74356 25288
rect 56152 25248 74356 25276
rect 74350 25236 74356 25248
rect 74408 25236 74414 25288
rect 90450 25236 90456 25288
rect 90508 25276 90514 25288
rect 90821 25279 90879 25285
rect 90821 25276 90833 25279
rect 90508 25248 90833 25276
rect 90508 25236 90514 25248
rect 90821 25245 90833 25248
rect 90867 25245 90879 25279
rect 91278 25276 91284 25288
rect 91239 25248 91284 25276
rect 90821 25239 90879 25245
rect 91278 25236 91284 25248
rect 91336 25236 91342 25288
rect 91388 25248 93854 25276
rect 53742 25208 53748 25220
rect 51368 25180 52040 25208
rect 52104 25180 53748 25208
rect 27816 25112 42288 25140
rect 43349 25143 43407 25149
rect 43349 25109 43361 25143
rect 43395 25140 43407 25143
rect 43622 25140 43628 25152
rect 43395 25112 43628 25140
rect 43395 25109 43407 25112
rect 43349 25103 43407 25109
rect 43622 25100 43628 25112
rect 43680 25100 43686 25152
rect 43714 25100 43720 25152
rect 43772 25140 43778 25152
rect 47486 25140 47492 25152
rect 43772 25112 47492 25140
rect 43772 25100 43778 25112
rect 47486 25100 47492 25112
rect 47544 25100 47550 25152
rect 50430 25100 50436 25152
rect 50488 25140 50494 25152
rect 52104 25140 52132 25180
rect 53742 25168 53748 25180
rect 53800 25168 53806 25220
rect 56778 25168 56784 25220
rect 56836 25208 56842 25220
rect 57514 25208 57520 25220
rect 56836 25180 57520 25208
rect 56836 25168 56842 25180
rect 57514 25168 57520 25180
rect 57572 25168 57578 25220
rect 59998 25168 60004 25220
rect 60056 25208 60062 25220
rect 60182 25208 60188 25220
rect 60056 25180 60188 25208
rect 60056 25168 60062 25180
rect 60182 25168 60188 25180
rect 60240 25168 60246 25220
rect 65610 25168 65616 25220
rect 65668 25208 65674 25220
rect 70210 25208 70216 25220
rect 65668 25180 70216 25208
rect 65668 25168 65674 25180
rect 70210 25168 70216 25180
rect 70268 25168 70274 25220
rect 73154 25168 73160 25220
rect 73212 25208 73218 25220
rect 91388 25208 91416 25248
rect 73212 25180 91416 25208
rect 93826 25208 93854 25248
rect 97442 25208 97448 25220
rect 93826 25180 97448 25208
rect 73212 25168 73218 25180
rect 97442 25168 97448 25180
rect 97500 25168 97506 25220
rect 52822 25140 52828 25152
rect 50488 25112 52132 25140
rect 52783 25112 52828 25140
rect 50488 25100 50494 25112
rect 52822 25100 52828 25112
rect 52880 25100 52886 25152
rect 53190 25100 53196 25152
rect 53248 25140 53254 25152
rect 54754 25140 54760 25152
rect 53248 25112 54760 25140
rect 53248 25100 53254 25112
rect 54754 25100 54760 25112
rect 54812 25140 54818 25152
rect 56502 25140 56508 25152
rect 54812 25112 56508 25140
rect 54812 25100 54818 25112
rect 56502 25100 56508 25112
rect 56560 25100 56566 25152
rect 56870 25100 56876 25152
rect 56928 25140 56934 25152
rect 90085 25143 90143 25149
rect 90085 25140 90097 25143
rect 56928 25112 90097 25140
rect 56928 25100 56934 25112
rect 90085 25109 90097 25112
rect 90131 25140 90143 25143
rect 90269 25143 90327 25149
rect 90269 25140 90281 25143
rect 90131 25112 90281 25140
rect 90131 25109 90143 25112
rect 90085 25103 90143 25109
rect 90269 25109 90281 25112
rect 90315 25140 90327 25143
rect 90453 25143 90511 25149
rect 90453 25140 90465 25143
rect 90315 25112 90465 25140
rect 90315 25109 90327 25112
rect 90269 25103 90327 25109
rect 90453 25109 90465 25112
rect 90499 25140 90511 25143
rect 91833 25143 91891 25149
rect 91833 25140 91845 25143
rect 90499 25112 91845 25140
rect 90499 25109 90511 25112
rect 90453 25103 90511 25109
rect 91833 25109 91845 25112
rect 91879 25140 91891 25143
rect 92109 25143 92167 25149
rect 92109 25140 92121 25143
rect 91879 25112 92121 25140
rect 91879 25109 91891 25112
rect 91833 25103 91891 25109
rect 92109 25109 92121 25112
rect 92155 25140 92167 25143
rect 92293 25143 92351 25149
rect 92293 25140 92305 25143
rect 92155 25112 92305 25140
rect 92155 25109 92167 25112
rect 92109 25103 92167 25109
rect 92293 25109 92305 25112
rect 92339 25140 92351 25143
rect 92477 25143 92535 25149
rect 92477 25140 92489 25143
rect 92339 25112 92489 25140
rect 92339 25109 92351 25112
rect 92293 25103 92351 25109
rect 92477 25109 92489 25112
rect 92523 25109 92535 25143
rect 92477 25103 92535 25109
rect 1104 25050 98808 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 65686 25050
rect 65738 24998 65750 25050
rect 65802 24998 65814 25050
rect 65866 24998 65878 25050
rect 65930 24998 96406 25050
rect 96458 24998 96470 25050
rect 96522 24998 96534 25050
rect 96586 24998 96598 25050
rect 96650 24998 98808 25050
rect 1104 24976 98808 24998
rect 9122 24896 9128 24948
rect 9180 24936 9186 24948
rect 13998 24936 14004 24948
rect 9180 24908 14004 24936
rect 9180 24896 9186 24908
rect 13998 24896 14004 24908
rect 14056 24896 14062 24948
rect 25866 24936 25872 24948
rect 17236 24908 25872 24936
rect 2225 24871 2283 24877
rect 2225 24837 2237 24871
rect 2271 24868 2283 24871
rect 2271 24840 2360 24868
rect 2271 24837 2283 24840
rect 2225 24831 2283 24837
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24800 1915 24803
rect 2332 24800 2360 24840
rect 4706 24828 4712 24880
rect 4764 24868 4770 24880
rect 17236 24868 17264 24908
rect 25866 24896 25872 24908
rect 25924 24896 25930 24948
rect 27706 24896 27712 24948
rect 27764 24936 27770 24948
rect 38286 24936 38292 24948
rect 27764 24908 38292 24936
rect 27764 24896 27770 24908
rect 38286 24896 38292 24908
rect 38344 24896 38350 24948
rect 38562 24896 38568 24948
rect 38620 24896 38626 24948
rect 39482 24896 39488 24948
rect 39540 24936 39546 24948
rect 39540 24908 52776 24936
rect 39540 24896 39546 24908
rect 36906 24868 36912 24880
rect 4764 24840 17264 24868
rect 30668 24840 36912 24868
rect 4764 24828 4770 24840
rect 3234 24800 3240 24812
rect 1903 24772 2268 24800
rect 2332 24772 3240 24800
rect 1903 24769 1915 24772
rect 1857 24763 1915 24769
rect 1486 24732 1492 24744
rect 1447 24704 1492 24732
rect 1486 24692 1492 24704
rect 1544 24692 1550 24744
rect 1672 24735 1730 24741
rect 1672 24701 1684 24735
rect 1718 24701 1730 24735
rect 1672 24695 1730 24701
rect 1688 24664 1716 24695
rect 1762 24692 1768 24744
rect 1820 24732 1826 24744
rect 2041 24735 2099 24741
rect 1820 24704 1865 24732
rect 1820 24692 1826 24704
rect 2041 24701 2053 24735
rect 2087 24732 2099 24735
rect 2130 24732 2136 24744
rect 2087 24704 2136 24732
rect 2087 24701 2099 24704
rect 2041 24695 2099 24701
rect 2130 24692 2136 24704
rect 2188 24692 2194 24744
rect 2240 24732 2268 24772
rect 3234 24760 3240 24772
rect 3292 24760 3298 24812
rect 3421 24803 3479 24809
rect 3421 24769 3433 24803
rect 3467 24769 3479 24803
rect 12710 24800 12716 24812
rect 3421 24763 3479 24769
rect 3896 24772 12716 24800
rect 2409 24735 2467 24741
rect 2409 24732 2421 24735
rect 2240 24704 2421 24732
rect 2409 24701 2421 24704
rect 2455 24732 2467 24735
rect 2866 24732 2872 24744
rect 2455 24704 2872 24732
rect 2455 24701 2467 24704
rect 2409 24695 2467 24701
rect 2866 24692 2872 24704
rect 2924 24732 2930 24744
rect 3050 24732 3056 24744
rect 2924 24704 3056 24732
rect 2924 24692 2930 24704
rect 3050 24692 3056 24704
rect 3108 24692 3114 24744
rect 3326 24732 3332 24744
rect 3287 24704 3332 24732
rect 3326 24692 3332 24704
rect 3384 24692 3390 24744
rect 1688 24636 2636 24664
rect 2608 24605 2636 24636
rect 2593 24599 2651 24605
rect 2593 24565 2605 24599
rect 2639 24596 2651 24599
rect 2682 24596 2688 24608
rect 2639 24568 2688 24596
rect 2639 24565 2651 24568
rect 2593 24559 2651 24565
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 2958 24596 2964 24608
rect 2919 24568 2964 24596
rect 2958 24556 2964 24568
rect 3016 24556 3022 24608
rect 3436 24596 3464 24763
rect 3694 24732 3700 24744
rect 3655 24704 3700 24732
rect 3694 24692 3700 24704
rect 3752 24692 3758 24744
rect 3896 24741 3924 24772
rect 12710 24760 12716 24772
rect 12768 24760 12774 24812
rect 12802 24760 12808 24812
rect 12860 24800 12866 24812
rect 16482 24800 16488 24812
rect 12860 24772 16488 24800
rect 12860 24760 12866 24772
rect 16482 24760 16488 24772
rect 16540 24760 16546 24812
rect 17126 24760 17132 24812
rect 17184 24800 17190 24812
rect 18414 24800 18420 24812
rect 17184 24772 18420 24800
rect 17184 24760 17190 24772
rect 18414 24760 18420 24772
rect 18472 24800 18478 24812
rect 24486 24800 24492 24812
rect 18472 24772 24492 24800
rect 18472 24760 18478 24772
rect 24486 24760 24492 24772
rect 24544 24760 24550 24812
rect 3881 24735 3939 24741
rect 3881 24701 3893 24735
rect 3927 24701 3939 24735
rect 3881 24695 3939 24701
rect 12161 24735 12219 24741
rect 12161 24701 12173 24735
rect 12207 24732 12219 24735
rect 12437 24735 12495 24741
rect 12437 24732 12449 24735
rect 12207 24704 12449 24732
rect 12207 24701 12219 24704
rect 12161 24695 12219 24701
rect 12437 24701 12449 24704
rect 12483 24732 12495 24735
rect 13446 24732 13452 24744
rect 12483 24704 13452 24732
rect 12483 24701 12495 24704
rect 12437 24695 12495 24701
rect 13446 24692 13452 24704
rect 13504 24692 13510 24744
rect 30668 24741 30696 24840
rect 36906 24828 36912 24840
rect 36964 24828 36970 24880
rect 37090 24828 37096 24880
rect 37148 24868 37154 24880
rect 38580 24868 38608 24896
rect 43530 24868 43536 24880
rect 37148 24840 43536 24868
rect 37148 24828 37154 24840
rect 43530 24828 43536 24840
rect 43588 24828 43594 24880
rect 44634 24828 44640 24880
rect 44692 24868 44698 24880
rect 50430 24868 50436 24880
rect 44692 24840 50436 24868
rect 44692 24828 44698 24840
rect 50430 24828 50436 24840
rect 50488 24828 50494 24880
rect 52748 24868 52776 24908
rect 52822 24896 52828 24948
rect 52880 24936 52886 24948
rect 66254 24936 66260 24948
rect 52880 24908 66260 24936
rect 52880 24896 52886 24908
rect 66254 24896 66260 24908
rect 66312 24896 66318 24948
rect 69290 24896 69296 24948
rect 69348 24936 69354 24948
rect 91278 24936 91284 24948
rect 69348 24908 91284 24936
rect 69348 24896 69354 24908
rect 91278 24896 91284 24908
rect 91336 24896 91342 24948
rect 56226 24868 56232 24880
rect 52748 24840 56232 24868
rect 56226 24828 56232 24840
rect 56284 24828 56290 24880
rect 56318 24828 56324 24880
rect 56376 24868 56382 24880
rect 69934 24868 69940 24880
rect 56376 24840 69940 24868
rect 56376 24828 56382 24840
rect 69934 24828 69940 24840
rect 69992 24828 69998 24880
rect 71406 24868 71412 24880
rect 71367 24840 71412 24868
rect 71406 24828 71412 24840
rect 71464 24828 71470 24880
rect 72694 24828 72700 24880
rect 72752 24868 72758 24880
rect 75822 24868 75828 24880
rect 72752 24840 75828 24868
rect 72752 24828 72758 24840
rect 75822 24828 75828 24840
rect 75880 24828 75886 24880
rect 35986 24760 35992 24812
rect 36044 24800 36050 24812
rect 50522 24800 50528 24812
rect 36044 24772 50528 24800
rect 36044 24760 36050 24772
rect 50522 24760 50528 24772
rect 50580 24760 50586 24812
rect 51350 24760 51356 24812
rect 51408 24800 51414 24812
rect 87966 24800 87972 24812
rect 51408 24772 87972 24800
rect 51408 24760 51414 24772
rect 87966 24760 87972 24772
rect 88024 24760 88030 24812
rect 30653 24735 30711 24741
rect 30653 24732 30665 24735
rect 22066 24704 30665 24732
rect 5074 24624 5080 24676
rect 5132 24664 5138 24676
rect 5350 24664 5356 24676
rect 5132 24636 5356 24664
rect 5132 24624 5138 24636
rect 5350 24624 5356 24636
rect 5408 24664 5414 24676
rect 22066 24664 22094 24704
rect 30653 24701 30665 24704
rect 30699 24701 30711 24735
rect 30653 24695 30711 24701
rect 36906 24692 36912 24744
rect 36964 24732 36970 24744
rect 39298 24732 39304 24744
rect 36964 24704 39304 24732
rect 36964 24692 36970 24704
rect 39298 24692 39304 24704
rect 39356 24732 39362 24744
rect 40494 24732 40500 24744
rect 39356 24704 40500 24732
rect 39356 24692 39362 24704
rect 40494 24692 40500 24704
rect 40552 24692 40558 24744
rect 40678 24692 40684 24744
rect 40736 24732 40742 24744
rect 41414 24732 41420 24744
rect 40736 24704 41420 24732
rect 40736 24692 40742 24704
rect 41414 24692 41420 24704
rect 41472 24732 41478 24744
rect 43533 24735 43591 24741
rect 43533 24732 43545 24735
rect 41472 24704 43545 24732
rect 41472 24692 41478 24704
rect 43533 24701 43545 24704
rect 43579 24701 43591 24735
rect 43806 24732 43812 24744
rect 43767 24704 43812 24732
rect 43533 24695 43591 24701
rect 43806 24692 43812 24704
rect 43864 24692 43870 24744
rect 44726 24692 44732 24744
rect 44784 24732 44790 24744
rect 44910 24732 44916 24744
rect 44784 24704 44916 24732
rect 44784 24692 44790 24704
rect 44910 24692 44916 24704
rect 44968 24732 44974 24744
rect 45189 24735 45247 24741
rect 45189 24732 45201 24735
rect 44968 24704 45201 24732
rect 44968 24692 44974 24704
rect 45189 24701 45201 24704
rect 45235 24701 45247 24735
rect 45189 24695 45247 24701
rect 45462 24692 45468 24744
rect 45520 24732 45526 24744
rect 47302 24732 47308 24744
rect 45520 24704 47308 24732
rect 45520 24692 45526 24704
rect 47302 24692 47308 24704
rect 47360 24692 47366 24744
rect 48774 24692 48780 24744
rect 48832 24732 48838 24744
rect 50893 24735 50951 24741
rect 50893 24732 50905 24735
rect 48832 24704 50905 24732
rect 48832 24692 48838 24704
rect 50893 24701 50905 24704
rect 50939 24732 50951 24735
rect 50982 24732 50988 24744
rect 50939 24704 50988 24732
rect 50939 24701 50951 24704
rect 50893 24695 50951 24701
rect 50982 24692 50988 24704
rect 51040 24692 51046 24744
rect 51166 24732 51172 24744
rect 51127 24704 51172 24732
rect 51166 24692 51172 24704
rect 51224 24692 51230 24744
rect 51534 24692 51540 24744
rect 51592 24732 51598 24744
rect 51592 24704 65472 24732
rect 51592 24692 51598 24704
rect 5408 24636 22094 24664
rect 5408 24624 5414 24636
rect 22738 24624 22744 24676
rect 22796 24664 22802 24676
rect 28074 24664 28080 24676
rect 22796 24636 28080 24664
rect 22796 24624 22802 24636
rect 28074 24624 28080 24636
rect 28132 24624 28138 24676
rect 29825 24667 29883 24673
rect 29825 24633 29837 24667
rect 29871 24664 29883 24667
rect 34238 24664 34244 24676
rect 29871 24636 34244 24664
rect 29871 24633 29883 24636
rect 29825 24627 29883 24633
rect 34238 24624 34244 24636
rect 34296 24624 34302 24676
rect 36998 24624 37004 24676
rect 37056 24664 37062 24676
rect 43622 24664 43628 24676
rect 37056 24636 43628 24664
rect 37056 24624 37062 24636
rect 43622 24624 43628 24636
rect 43680 24624 43686 24676
rect 44836 24636 45048 24664
rect 14734 24596 14740 24608
rect 3436 24568 14740 24596
rect 14734 24556 14740 24568
rect 14792 24556 14798 24608
rect 18046 24556 18052 24608
rect 18104 24596 18110 24608
rect 22554 24596 22560 24608
rect 18104 24568 22560 24596
rect 18104 24556 18110 24568
rect 22554 24556 22560 24568
rect 22612 24556 22618 24608
rect 23106 24556 23112 24608
rect 23164 24596 23170 24608
rect 30374 24596 30380 24608
rect 23164 24568 30380 24596
rect 23164 24556 23170 24568
rect 30374 24556 30380 24568
rect 30432 24556 30438 24608
rect 30834 24556 30840 24608
rect 30892 24596 30898 24608
rect 44836 24596 44864 24636
rect 30892 24568 44864 24596
rect 45020 24596 45048 24636
rect 46106 24624 46112 24676
rect 46164 24664 46170 24676
rect 50522 24664 50528 24676
rect 46164 24636 50528 24664
rect 46164 24624 46170 24636
rect 50522 24624 50528 24636
rect 50580 24624 50586 24676
rect 52196 24636 52875 24664
rect 52196 24596 52224 24636
rect 52454 24596 52460 24608
rect 45020 24568 52224 24596
rect 52415 24568 52460 24596
rect 30892 24556 30898 24568
rect 52454 24556 52460 24568
rect 52512 24556 52518 24608
rect 52847 24596 52875 24636
rect 55674 24624 55680 24676
rect 55732 24664 55738 24676
rect 63402 24664 63408 24676
rect 55732 24636 63408 24664
rect 55732 24624 55738 24636
rect 63402 24624 63408 24636
rect 63460 24624 63466 24676
rect 65444 24664 65472 24704
rect 65518 24692 65524 24744
rect 65576 24732 65582 24744
rect 72786 24732 72792 24744
rect 65576 24704 72792 24732
rect 65576 24692 65582 24704
rect 72786 24692 72792 24704
rect 72844 24692 72850 24744
rect 78033 24735 78091 24741
rect 78033 24732 78045 24735
rect 76760 24704 78045 24732
rect 66898 24664 66904 24676
rect 65444 24636 66904 24664
rect 66898 24624 66904 24636
rect 66956 24624 66962 24676
rect 67266 24624 67272 24676
rect 67324 24664 67330 24676
rect 74626 24664 74632 24676
rect 67324 24636 74632 24664
rect 67324 24624 67330 24636
rect 74626 24624 74632 24636
rect 74684 24624 74690 24676
rect 75638 24624 75644 24676
rect 75696 24664 75702 24676
rect 76653 24667 76711 24673
rect 76653 24664 76665 24667
rect 75696 24636 76665 24664
rect 75696 24624 75702 24636
rect 76653 24633 76665 24636
rect 76699 24633 76711 24667
rect 76653 24627 76711 24633
rect 76101 24599 76159 24605
rect 76101 24596 76113 24599
rect 52847 24568 76113 24596
rect 76101 24565 76113 24568
rect 76147 24596 76159 24599
rect 76285 24599 76343 24605
rect 76285 24596 76297 24599
rect 76147 24568 76297 24596
rect 76147 24565 76159 24568
rect 76101 24559 76159 24565
rect 76285 24565 76297 24568
rect 76331 24596 76343 24599
rect 76469 24599 76527 24605
rect 76469 24596 76481 24599
rect 76331 24568 76481 24596
rect 76331 24565 76343 24568
rect 76285 24559 76343 24565
rect 76469 24565 76481 24568
rect 76515 24596 76527 24599
rect 76760 24596 76788 24704
rect 78033 24701 78045 24704
rect 78079 24732 78091 24735
rect 78079 24704 78260 24732
rect 78079 24701 78091 24704
rect 78033 24695 78091 24701
rect 78232 24664 78260 24704
rect 78306 24692 78312 24744
rect 78364 24732 78370 24744
rect 78364 24704 78409 24732
rect 78364 24692 78370 24704
rect 78401 24667 78459 24673
rect 78401 24664 78413 24667
rect 78232 24636 78413 24664
rect 78401 24633 78413 24636
rect 78447 24664 78459 24667
rect 78585 24667 78643 24673
rect 78585 24664 78597 24667
rect 78447 24636 78597 24664
rect 78447 24633 78459 24636
rect 78401 24627 78459 24633
rect 78585 24633 78597 24636
rect 78631 24664 78643 24667
rect 78769 24667 78827 24673
rect 78769 24664 78781 24667
rect 78631 24636 78781 24664
rect 78631 24633 78643 24636
rect 78585 24627 78643 24633
rect 78769 24633 78781 24636
rect 78815 24633 78827 24667
rect 78769 24627 78827 24633
rect 76515 24568 76788 24596
rect 76515 24565 76527 24568
rect 76469 24559 76527 24565
rect 1104 24506 98808 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 50326 24506
rect 50378 24454 50390 24506
rect 50442 24454 50454 24506
rect 50506 24454 50518 24506
rect 50570 24454 81046 24506
rect 81098 24454 81110 24506
rect 81162 24454 81174 24506
rect 81226 24454 81238 24506
rect 81290 24454 98808 24506
rect 1104 24432 98808 24454
rect 3694 24352 3700 24404
rect 3752 24392 3758 24404
rect 12618 24392 12624 24404
rect 3752 24364 12624 24392
rect 3752 24352 3758 24364
rect 12618 24352 12624 24364
rect 12676 24392 12682 24404
rect 13354 24392 13360 24404
rect 12676 24364 13360 24392
rect 12676 24352 12682 24364
rect 13354 24352 13360 24364
rect 13412 24352 13418 24404
rect 17589 24395 17647 24401
rect 17589 24392 17601 24395
rect 17328 24364 17601 24392
rect 15102 24284 15108 24336
rect 15160 24324 15166 24336
rect 17328 24324 17356 24364
rect 17589 24361 17601 24364
rect 17635 24392 17647 24395
rect 21818 24392 21824 24404
rect 17635 24364 21680 24392
rect 21779 24364 21824 24392
rect 17635 24361 17647 24364
rect 17589 24355 17647 24361
rect 15160 24296 17356 24324
rect 15160 24284 15166 24296
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 4706 24256 4712 24268
rect 3283 24228 4712 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 4706 24216 4712 24228
rect 4764 24216 4770 24268
rect 16761 24259 16819 24265
rect 16761 24225 16773 24259
rect 16807 24225 16819 24259
rect 16761 24219 16819 24225
rect 16853 24259 16911 24265
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 16942 24256 16948 24268
rect 16899 24228 16948 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 10594 24148 10600 24200
rect 10652 24188 10658 24200
rect 10870 24188 10876 24200
rect 10652 24160 10876 24188
rect 10652 24148 10658 24160
rect 10870 24148 10876 24160
rect 10928 24188 10934 24200
rect 16025 24191 16083 24197
rect 16025 24188 16037 24191
rect 10928 24160 16037 24188
rect 10928 24148 10934 24160
rect 16025 24157 16037 24160
rect 16071 24188 16083 24191
rect 16776 24188 16804 24219
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 17126 24256 17132 24268
rect 17087 24228 17132 24256
rect 17126 24216 17132 24228
rect 17184 24216 17190 24268
rect 17328 24265 17356 24296
rect 17420 24296 17632 24324
rect 17313 24259 17371 24265
rect 17313 24225 17325 24259
rect 17359 24225 17371 24259
rect 17313 24219 17371 24225
rect 17420 24188 17448 24296
rect 17497 24259 17555 24265
rect 17497 24225 17509 24259
rect 17543 24225 17555 24259
rect 17604 24256 17632 24296
rect 19058 24284 19064 24336
rect 19116 24324 19122 24336
rect 20349 24327 20407 24333
rect 20349 24324 20361 24327
rect 19116 24296 20361 24324
rect 19116 24284 19122 24296
rect 20349 24293 20361 24296
rect 20395 24293 20407 24327
rect 21652 24324 21680 24364
rect 21818 24352 21824 24364
rect 21876 24352 21882 24404
rect 25130 24352 25136 24404
rect 25188 24392 25194 24404
rect 43530 24392 43536 24404
rect 25188 24364 43536 24392
rect 25188 24352 25194 24364
rect 43530 24352 43536 24364
rect 43588 24352 43594 24404
rect 43990 24352 43996 24404
rect 44048 24392 44054 24404
rect 44048 24364 46796 24392
rect 44048 24352 44054 24364
rect 25314 24324 25320 24336
rect 21652 24296 25320 24324
rect 20349 24287 20407 24293
rect 25314 24284 25320 24296
rect 25372 24284 25378 24336
rect 36081 24327 36139 24333
rect 36081 24293 36093 24327
rect 36127 24324 36139 24327
rect 42794 24324 42800 24336
rect 36127 24296 42800 24324
rect 36127 24293 36139 24296
rect 36081 24287 36139 24293
rect 42794 24284 42800 24296
rect 42852 24284 42858 24336
rect 43622 24284 43628 24336
rect 43680 24324 43686 24336
rect 46106 24324 46112 24336
rect 43680 24296 46112 24324
rect 43680 24284 43686 24296
rect 46106 24284 46112 24296
rect 46164 24284 46170 24336
rect 46382 24324 46388 24336
rect 46343 24296 46388 24324
rect 46382 24284 46388 24296
rect 46440 24284 46446 24336
rect 46474 24284 46480 24336
rect 46532 24324 46538 24336
rect 46532 24296 46577 24324
rect 46532 24284 46538 24296
rect 46658 24284 46664 24336
rect 46716 24284 46722 24336
rect 22554 24256 22560 24268
rect 17604 24228 21312 24256
rect 22467 24228 22560 24256
rect 17497 24219 17555 24225
rect 16071 24160 17448 24188
rect 17512 24188 17540 24219
rect 19610 24188 19616 24200
rect 17512 24160 19616 24188
rect 16071 24157 16083 24160
rect 16025 24151 16083 24157
rect 19610 24148 19616 24160
rect 19668 24148 19674 24200
rect 20349 24191 20407 24197
rect 20349 24157 20361 24191
rect 20395 24188 20407 24191
rect 20441 24191 20499 24197
rect 20441 24188 20453 24191
rect 20395 24160 20453 24188
rect 20395 24157 20407 24160
rect 20349 24151 20407 24157
rect 20441 24157 20453 24160
rect 20487 24157 20499 24191
rect 20714 24188 20720 24200
rect 20675 24160 20720 24188
rect 20441 24151 20499 24157
rect 20714 24148 20720 24160
rect 20772 24148 20778 24200
rect 21284 24188 21312 24228
rect 22554 24216 22560 24228
rect 22612 24256 22618 24268
rect 40957 24259 41015 24265
rect 40957 24256 40969 24259
rect 22612 24228 40969 24256
rect 22612 24216 22618 24228
rect 40957 24225 40969 24228
rect 41003 24256 41015 24259
rect 42242 24256 42248 24268
rect 41003 24228 42248 24256
rect 41003 24225 41015 24228
rect 40957 24219 41015 24225
rect 42242 24216 42248 24228
rect 42300 24216 42306 24268
rect 44358 24216 44364 24268
rect 44416 24256 44422 24268
rect 44726 24256 44732 24268
rect 44416 24228 44732 24256
rect 44416 24216 44422 24228
rect 44726 24216 44732 24228
rect 44784 24216 44790 24268
rect 46201 24259 46259 24265
rect 46201 24225 46213 24259
rect 46247 24256 46259 24259
rect 46290 24256 46296 24268
rect 46247 24228 46296 24256
rect 46247 24225 46259 24228
rect 46201 24219 46259 24225
rect 46290 24216 46296 24228
rect 46348 24216 46354 24268
rect 46569 24259 46627 24265
rect 46569 24225 46581 24259
rect 46615 24225 46627 24259
rect 46569 24219 46627 24225
rect 23014 24188 23020 24200
rect 21284 24160 23020 24188
rect 23014 24148 23020 24160
rect 23072 24148 23078 24200
rect 23290 24188 23296 24200
rect 23251 24160 23296 24188
rect 23290 24148 23296 24160
rect 23348 24148 23354 24200
rect 24210 24148 24216 24200
rect 24268 24188 24274 24200
rect 24762 24188 24768 24200
rect 24268 24160 24768 24188
rect 24268 24148 24274 24160
rect 24762 24148 24768 24160
rect 24820 24188 24826 24200
rect 25222 24188 25228 24200
rect 24820 24160 25228 24188
rect 24820 24148 24826 24160
rect 25222 24148 25228 24160
rect 25280 24148 25286 24200
rect 25314 24148 25320 24200
rect 25372 24188 25378 24200
rect 43990 24188 43996 24200
rect 25372 24160 43996 24188
rect 25372 24148 25378 24160
rect 43990 24148 43996 24160
rect 44048 24148 44054 24200
rect 45370 24148 45376 24200
rect 45428 24188 45434 24200
rect 45830 24188 45836 24200
rect 45428 24160 45836 24188
rect 45428 24148 45434 24160
rect 45830 24148 45836 24160
rect 45888 24148 45894 24200
rect 16393 24123 16451 24129
rect 16393 24089 16405 24123
rect 16439 24120 16451 24123
rect 40954 24120 40960 24132
rect 16439 24092 20484 24120
rect 16439 24089 16451 24092
rect 16393 24083 16451 24089
rect 3237 24055 3295 24061
rect 3237 24021 3249 24055
rect 3283 24052 3295 24055
rect 11146 24052 11152 24064
rect 3283 24024 11152 24052
rect 3283 24021 3295 24024
rect 3237 24015 3295 24021
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 19518 24012 19524 24064
rect 19576 24052 19582 24064
rect 20162 24052 20168 24064
rect 19576 24024 20168 24052
rect 19576 24012 19582 24024
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 20456 24052 20484 24092
rect 21376 24092 40960 24120
rect 21376 24052 21404 24092
rect 40954 24080 40960 24092
rect 41012 24080 41018 24132
rect 41046 24080 41052 24132
rect 41104 24120 41110 24132
rect 41141 24123 41199 24129
rect 41141 24120 41153 24123
rect 41104 24092 41153 24120
rect 41104 24080 41110 24092
rect 41141 24089 41153 24092
rect 41187 24089 41199 24123
rect 41141 24083 41199 24089
rect 46382 24080 46388 24132
rect 46440 24120 46446 24132
rect 46584 24120 46612 24219
rect 46440 24092 46612 24120
rect 46676 24120 46704 24284
rect 46768 24188 46796 24364
rect 46934 24352 46940 24404
rect 46992 24392 46998 24404
rect 65518 24392 65524 24404
rect 46992 24364 65524 24392
rect 46992 24352 46998 24364
rect 65518 24352 65524 24364
rect 65576 24352 65582 24404
rect 74994 24392 75000 24404
rect 65628 24364 75000 24392
rect 48130 24284 48136 24336
rect 48188 24324 48194 24336
rect 63494 24324 63500 24336
rect 48188 24296 63500 24324
rect 48188 24284 48194 24296
rect 63494 24284 63500 24296
rect 63552 24284 63558 24336
rect 65245 24327 65303 24333
rect 65245 24293 65257 24327
rect 65291 24324 65303 24327
rect 65628 24324 65656 24364
rect 74994 24352 75000 24364
rect 75052 24352 75058 24404
rect 86862 24392 86868 24404
rect 75104 24364 77294 24392
rect 65291 24296 65656 24324
rect 65291 24293 65303 24296
rect 65245 24287 65303 24293
rect 66254 24284 66260 24336
rect 66312 24324 66318 24336
rect 72694 24324 72700 24336
rect 66312 24296 72700 24324
rect 66312 24284 66318 24296
rect 72694 24284 72700 24296
rect 72752 24284 72758 24336
rect 72786 24284 72792 24336
rect 72844 24324 72850 24336
rect 75104 24324 75132 24364
rect 75822 24324 75828 24336
rect 72844 24296 75132 24324
rect 75783 24296 75828 24324
rect 72844 24284 72850 24296
rect 75822 24284 75828 24296
rect 75880 24284 75886 24336
rect 77266 24324 77294 24364
rect 80026 24364 86868 24392
rect 80026 24324 80054 24364
rect 86862 24352 86868 24364
rect 86920 24352 86926 24404
rect 91922 24392 91928 24404
rect 89686 24364 91928 24392
rect 89686 24324 89714 24364
rect 91922 24352 91928 24364
rect 91980 24352 91986 24404
rect 77266 24296 80054 24324
rect 83108 24296 89714 24324
rect 47302 24216 47308 24268
rect 47360 24256 47366 24268
rect 75086 24256 75092 24268
rect 47360 24228 75092 24256
rect 47360 24216 47366 24228
rect 75086 24216 75092 24228
rect 75144 24256 75150 24268
rect 75365 24259 75423 24265
rect 75365 24256 75377 24259
rect 75144 24228 75377 24256
rect 75144 24216 75150 24228
rect 75365 24225 75377 24228
rect 75411 24256 75423 24259
rect 75549 24259 75607 24265
rect 75549 24256 75561 24259
rect 75411 24228 75561 24256
rect 75411 24225 75423 24228
rect 75365 24219 75423 24225
rect 75549 24225 75561 24228
rect 75595 24225 75607 24259
rect 75730 24256 75736 24268
rect 75691 24228 75736 24256
rect 75549 24219 75607 24225
rect 75730 24216 75736 24228
rect 75788 24216 75794 24268
rect 75914 24216 75920 24268
rect 75972 24256 75978 24268
rect 78306 24256 78312 24268
rect 75972 24228 76017 24256
rect 76116 24228 78312 24256
rect 75972 24216 75978 24228
rect 72786 24188 72792 24200
rect 46768 24160 72792 24188
rect 72786 24148 72792 24160
rect 72844 24148 72850 24200
rect 46753 24123 46811 24129
rect 46753 24120 46765 24123
rect 46676 24092 46765 24120
rect 46440 24080 46446 24092
rect 46753 24089 46765 24092
rect 46799 24089 46811 24123
rect 46753 24083 46811 24089
rect 46934 24080 46940 24132
rect 46992 24120 46998 24132
rect 55674 24120 55680 24132
rect 46992 24092 55680 24120
rect 46992 24080 46998 24092
rect 55674 24080 55680 24092
rect 55732 24080 55738 24132
rect 60706 24092 70394 24120
rect 20456 24024 21404 24052
rect 23014 24012 23020 24064
rect 23072 24052 23078 24064
rect 26878 24052 26884 24064
rect 23072 24024 26884 24052
rect 23072 24012 23078 24024
rect 26878 24012 26884 24024
rect 26936 24012 26942 24064
rect 28534 24012 28540 24064
rect 28592 24052 28598 24064
rect 35986 24052 35992 24064
rect 28592 24024 35992 24052
rect 28592 24012 28598 24024
rect 35986 24012 35992 24024
rect 36044 24012 36050 24064
rect 36081 24055 36139 24061
rect 36081 24021 36093 24055
rect 36127 24052 36139 24055
rect 36357 24055 36415 24061
rect 36357 24052 36369 24055
rect 36127 24024 36369 24052
rect 36127 24021 36139 24024
rect 36081 24015 36139 24021
rect 36357 24021 36369 24024
rect 36403 24021 36415 24055
rect 36357 24015 36415 24021
rect 36446 24012 36452 24064
rect 36504 24052 36510 24064
rect 43254 24052 43260 24064
rect 36504 24024 43260 24052
rect 36504 24012 36510 24024
rect 43254 24012 43260 24024
rect 43312 24012 43318 24064
rect 44082 24012 44088 24064
rect 44140 24052 44146 24064
rect 60706 24052 60734 24092
rect 44140 24024 60734 24052
rect 44140 24012 44146 24024
rect 61194 24012 61200 24064
rect 61252 24052 61258 24064
rect 63218 24052 63224 24064
rect 61252 24024 63224 24052
rect 61252 24012 61258 24024
rect 63218 24012 63224 24024
rect 63276 24012 63282 24064
rect 63402 24012 63408 24064
rect 63460 24052 63466 24064
rect 65245 24055 65303 24061
rect 65245 24052 65257 24055
rect 63460 24024 65257 24052
rect 63460 24012 63466 24024
rect 65245 24021 65257 24024
rect 65291 24021 65303 24055
rect 65245 24015 65303 24021
rect 65426 24012 65432 24064
rect 65484 24052 65490 24064
rect 65521 24055 65579 24061
rect 65521 24052 65533 24055
rect 65484 24024 65533 24052
rect 65484 24012 65490 24024
rect 65521 24021 65533 24024
rect 65567 24021 65579 24055
rect 70366 24052 70394 24092
rect 71682 24080 71688 24132
rect 71740 24120 71746 24132
rect 74718 24120 74724 24132
rect 71740 24092 74724 24120
rect 71740 24080 71746 24092
rect 74718 24080 74724 24092
rect 74776 24080 74782 24132
rect 75086 24080 75092 24132
rect 75144 24120 75150 24132
rect 76116 24120 76144 24228
rect 78306 24216 78312 24228
rect 78364 24216 78370 24268
rect 78490 24216 78496 24268
rect 78548 24256 78554 24268
rect 83001 24259 83059 24265
rect 83001 24256 83013 24259
rect 78548 24228 83013 24256
rect 78548 24216 78554 24228
rect 83001 24225 83013 24228
rect 83047 24225 83059 24259
rect 83001 24219 83059 24225
rect 76282 24188 76288 24200
rect 76243 24160 76288 24188
rect 76282 24148 76288 24160
rect 76340 24148 76346 24200
rect 76374 24148 76380 24200
rect 76432 24188 76438 24200
rect 83108 24188 83136 24296
rect 90174 24284 90180 24336
rect 90232 24324 90238 24336
rect 90818 24324 90824 24336
rect 90232 24296 90824 24324
rect 90232 24284 90238 24296
rect 90818 24284 90824 24296
rect 90876 24284 90882 24336
rect 83182 24216 83188 24268
rect 83240 24256 83246 24268
rect 83550 24256 83556 24268
rect 83240 24228 83284 24256
rect 83463 24228 83556 24256
rect 83240 24216 83246 24228
rect 83550 24216 83556 24228
rect 83608 24256 83614 24268
rect 95326 24256 95332 24268
rect 83608 24228 95332 24256
rect 83608 24216 83614 24228
rect 95326 24216 95332 24228
rect 95384 24216 95390 24268
rect 76432 24160 83136 24188
rect 83277 24191 83335 24197
rect 76432 24148 76438 24160
rect 83277 24157 83289 24191
rect 83323 24157 83335 24191
rect 83277 24151 83335 24157
rect 83369 24191 83427 24197
rect 83369 24157 83381 24191
rect 83415 24188 83427 24191
rect 84010 24188 84016 24200
rect 83415 24160 84016 24188
rect 83415 24157 83427 24160
rect 83369 24151 83427 24157
rect 83292 24120 83320 24151
rect 84010 24148 84016 24160
rect 84068 24148 84074 24200
rect 75144 24092 76144 24120
rect 76208 24092 83320 24120
rect 75144 24080 75150 24092
rect 76006 24052 76012 24064
rect 70366 24024 76012 24052
rect 65521 24015 65579 24021
rect 76006 24012 76012 24024
rect 76064 24012 76070 24064
rect 76101 24055 76159 24061
rect 76101 24021 76113 24055
rect 76147 24052 76159 24055
rect 76208 24052 76236 24092
rect 76147 24024 76236 24052
rect 76147 24021 76159 24024
rect 76101 24015 76159 24021
rect 76282 24012 76288 24064
rect 76340 24052 76346 24064
rect 83645 24055 83703 24061
rect 83645 24052 83657 24055
rect 76340 24024 83657 24052
rect 76340 24012 76346 24024
rect 83645 24021 83657 24024
rect 83691 24021 83703 24055
rect 83645 24015 83703 24021
rect 1104 23962 98808 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 65686 23962
rect 65738 23910 65750 23962
rect 65802 23910 65814 23962
rect 65866 23910 65878 23962
rect 65930 23910 96406 23962
rect 96458 23910 96470 23962
rect 96522 23910 96534 23962
rect 96586 23910 96598 23962
rect 96650 23910 98808 23962
rect 1104 23888 98808 23910
rect 1762 23808 1768 23860
rect 1820 23848 1826 23860
rect 9490 23848 9496 23860
rect 1820 23820 9496 23848
rect 1820 23808 1826 23820
rect 9490 23808 9496 23820
rect 9548 23848 9554 23860
rect 19518 23848 19524 23860
rect 9548 23820 19524 23848
rect 9548 23808 9554 23820
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 19610 23808 19616 23860
rect 19668 23848 19674 23860
rect 20530 23848 20536 23860
rect 19668 23820 20536 23848
rect 19668 23808 19674 23820
rect 20530 23808 20536 23820
rect 20588 23848 20594 23860
rect 35526 23848 35532 23860
rect 20588 23820 35532 23848
rect 20588 23808 20594 23820
rect 35526 23808 35532 23820
rect 35584 23808 35590 23860
rect 35802 23808 35808 23860
rect 35860 23848 35866 23860
rect 35860 23820 36676 23848
rect 35860 23808 35866 23820
rect 2682 23740 2688 23792
rect 2740 23780 2746 23792
rect 20622 23780 20628 23792
rect 2740 23752 20628 23780
rect 2740 23740 2746 23752
rect 20622 23740 20628 23752
rect 20680 23780 20686 23792
rect 25130 23780 25136 23792
rect 20680 23752 25136 23780
rect 20680 23740 20686 23752
rect 25130 23740 25136 23752
rect 25188 23740 25194 23792
rect 25222 23740 25228 23792
rect 25280 23780 25286 23792
rect 25280 23752 25325 23780
rect 31726 23752 36584 23780
rect 25280 23740 25286 23752
rect 13354 23672 13360 23724
rect 13412 23712 13418 23724
rect 23934 23712 23940 23724
rect 13412 23684 23940 23712
rect 13412 23672 13418 23684
rect 23934 23672 23940 23684
rect 23992 23712 23998 23724
rect 24302 23712 24308 23724
rect 23992 23684 24308 23712
rect 23992 23672 23998 23684
rect 24302 23672 24308 23684
rect 24360 23672 24366 23724
rect 25317 23715 25375 23721
rect 24964 23684 25268 23712
rect 4801 23647 4859 23653
rect 4801 23613 4813 23647
rect 4847 23613 4859 23647
rect 4801 23607 4859 23613
rect 14461 23647 14519 23653
rect 14461 23613 14473 23647
rect 14507 23644 14519 23647
rect 24964 23644 24992 23684
rect 25130 23653 25136 23656
rect 14507 23616 24992 23644
rect 25096 23647 25136 23653
rect 14507 23613 14519 23616
rect 14461 23607 14519 23613
rect 25096 23613 25108 23647
rect 25096 23607 25136 23613
rect 4525 23579 4583 23585
rect 4525 23545 4537 23579
rect 4571 23576 4583 23579
rect 4816 23576 4844 23607
rect 25130 23604 25136 23607
rect 25188 23604 25194 23656
rect 25240 23644 25268 23684
rect 25317 23681 25329 23715
rect 25363 23712 25375 23715
rect 25682 23712 25688 23724
rect 25363 23684 25688 23712
rect 25363 23681 25375 23684
rect 25317 23675 25375 23681
rect 25682 23672 25688 23684
rect 25740 23672 25746 23724
rect 31726 23644 31754 23752
rect 34422 23672 34428 23724
rect 34480 23712 34486 23724
rect 36446 23712 36452 23724
rect 34480 23684 36452 23712
rect 34480 23672 34486 23684
rect 36446 23672 36452 23684
rect 36504 23672 36510 23724
rect 25240 23616 31754 23644
rect 36556 23644 36584 23752
rect 36648 23712 36676 23820
rect 43254 23808 43260 23860
rect 43312 23848 43318 23860
rect 45186 23848 45192 23860
rect 43312 23820 45192 23848
rect 43312 23808 43318 23820
rect 45186 23808 45192 23820
rect 45244 23808 45250 23860
rect 50338 23848 50344 23860
rect 45296 23820 50344 23848
rect 37734 23740 37740 23792
rect 37792 23780 37798 23792
rect 45002 23780 45008 23792
rect 37792 23752 45008 23780
rect 37792 23740 37798 23752
rect 45002 23740 45008 23752
rect 45060 23740 45066 23792
rect 42978 23712 42984 23724
rect 36648 23684 42984 23712
rect 42978 23672 42984 23684
rect 43036 23672 43042 23724
rect 43254 23672 43260 23724
rect 43312 23712 43318 23724
rect 43806 23712 43812 23724
rect 43312 23684 43812 23712
rect 43312 23672 43318 23684
rect 43806 23672 43812 23684
rect 43864 23672 43870 23724
rect 45296 23644 45324 23820
rect 50338 23808 50344 23820
rect 50396 23808 50402 23860
rect 51046 23820 76052 23848
rect 45370 23740 45376 23792
rect 45428 23780 45434 23792
rect 48682 23780 48688 23792
rect 45428 23752 48688 23780
rect 45428 23740 45434 23752
rect 48682 23740 48688 23752
rect 48740 23740 48746 23792
rect 50157 23783 50215 23789
rect 50157 23749 50169 23783
rect 50203 23780 50215 23783
rect 50614 23780 50620 23792
rect 50203 23752 50620 23780
rect 50203 23749 50215 23752
rect 50157 23743 50215 23749
rect 50614 23740 50620 23752
rect 50672 23780 50678 23792
rect 51046 23780 51074 23820
rect 50672 23752 51074 23780
rect 50672 23740 50678 23752
rect 53558 23740 53564 23792
rect 53616 23780 53622 23792
rect 63402 23780 63408 23792
rect 53616 23752 63408 23780
rect 53616 23740 53622 23752
rect 63402 23740 63408 23752
rect 63460 23740 63466 23792
rect 63494 23740 63500 23792
rect 63552 23780 63558 23792
rect 66349 23783 66407 23789
rect 66349 23780 66361 23783
rect 63552 23752 66361 23780
rect 63552 23740 63558 23752
rect 66349 23749 66361 23752
rect 66395 23749 66407 23783
rect 69934 23780 69940 23792
rect 69895 23752 69940 23780
rect 66349 23743 66407 23749
rect 69934 23740 69940 23752
rect 69992 23740 69998 23792
rect 72145 23783 72203 23789
rect 72145 23749 72157 23783
rect 72191 23780 72203 23783
rect 73154 23780 73160 23792
rect 72191 23752 73160 23780
rect 72191 23749 72203 23752
rect 72145 23743 72203 23749
rect 46198 23672 46204 23724
rect 46256 23712 46262 23724
rect 46658 23712 46664 23724
rect 46256 23684 46664 23712
rect 46256 23672 46262 23684
rect 46658 23672 46664 23684
rect 46716 23672 46722 23724
rect 48774 23712 48780 23724
rect 48735 23684 48780 23712
rect 48774 23672 48780 23684
rect 48832 23672 48838 23724
rect 49053 23715 49111 23721
rect 49053 23681 49065 23715
rect 49099 23712 49111 23715
rect 71866 23712 71872 23724
rect 49099 23684 71872 23712
rect 49099 23681 49111 23684
rect 49053 23675 49111 23681
rect 71866 23672 71872 23684
rect 71924 23672 71930 23724
rect 36556 23616 45324 23644
rect 47026 23604 47032 23656
rect 47084 23644 47090 23656
rect 48682 23644 48688 23656
rect 47084 23616 48688 23644
rect 47084 23604 47090 23616
rect 48682 23604 48688 23616
rect 48740 23604 48746 23656
rect 65610 23644 65616 23656
rect 48884 23616 65616 23644
rect 22094 23576 22100 23588
rect 4571 23548 22100 23576
rect 4571 23545 4583 23548
rect 4525 23539 4583 23545
rect 22094 23536 22100 23548
rect 22152 23536 22158 23588
rect 24946 23576 24952 23588
rect 24907 23548 24952 23576
rect 24946 23536 24952 23548
rect 25004 23536 25010 23588
rect 25148 23548 25728 23576
rect 18230 23468 18236 23520
rect 18288 23508 18294 23520
rect 25148 23508 25176 23548
rect 25590 23508 25596 23520
rect 18288 23480 25176 23508
rect 25551 23480 25596 23508
rect 18288 23468 18294 23480
rect 25590 23468 25596 23480
rect 25648 23468 25654 23520
rect 25700 23508 25728 23548
rect 26878 23536 26884 23588
rect 26936 23576 26942 23588
rect 34330 23576 34336 23588
rect 26936 23548 34336 23576
rect 26936 23536 26942 23548
rect 34330 23536 34336 23548
rect 34388 23576 34394 23588
rect 48884 23576 48912 23616
rect 65610 23604 65616 23616
rect 65668 23604 65674 23656
rect 65886 23604 65892 23656
rect 65944 23604 65950 23656
rect 66073 23647 66131 23653
rect 66073 23613 66085 23647
rect 66119 23644 66131 23647
rect 69014 23644 69020 23656
rect 66119 23616 69020 23644
rect 66119 23613 66131 23616
rect 66073 23607 66131 23613
rect 69014 23604 69020 23616
rect 69072 23604 69078 23656
rect 72237 23647 72295 23653
rect 72237 23613 72249 23647
rect 72283 23613 72295 23647
rect 72237 23607 72295 23613
rect 34388 23548 48912 23576
rect 49712 23548 50292 23576
rect 34388 23536 34394 23548
rect 49712 23508 49740 23548
rect 25700 23480 49740 23508
rect 50264 23508 50292 23548
rect 50338 23536 50344 23588
rect 50396 23576 50402 23588
rect 61378 23576 61384 23588
rect 50396 23548 61384 23576
rect 50396 23536 50402 23548
rect 61378 23536 61384 23548
rect 61436 23536 61442 23588
rect 61746 23536 61752 23588
rect 61804 23576 61810 23588
rect 65426 23576 65432 23588
rect 61804 23548 65432 23576
rect 61804 23536 61810 23548
rect 65426 23536 65432 23548
rect 65484 23536 65490 23588
rect 65797 23579 65855 23585
rect 65797 23576 65809 23579
rect 65720 23548 65809 23576
rect 65521 23511 65579 23517
rect 65521 23508 65533 23511
rect 50264 23480 65533 23508
rect 65521 23477 65533 23480
rect 65567 23508 65579 23511
rect 65720 23508 65748 23548
rect 65797 23545 65809 23548
rect 65843 23545 65855 23579
rect 65904 23576 65932 23604
rect 72252 23576 72280 23607
rect 72344 23576 72372 23752
rect 73154 23740 73160 23752
rect 73212 23740 73218 23792
rect 76024 23712 76052 23820
rect 76098 23808 76104 23860
rect 76156 23848 76162 23860
rect 76929 23851 76987 23857
rect 76929 23848 76941 23851
rect 76156 23820 76941 23848
rect 76156 23808 76162 23820
rect 76929 23817 76941 23820
rect 76975 23817 76987 23851
rect 76929 23811 76987 23817
rect 80054 23808 80060 23860
rect 80112 23848 80118 23860
rect 80241 23851 80299 23857
rect 80241 23848 80253 23851
rect 80112 23820 80253 23848
rect 80112 23808 80118 23820
rect 80241 23817 80253 23820
rect 80287 23817 80299 23851
rect 84010 23848 84016 23860
rect 80241 23811 80299 23817
rect 81728 23820 84016 23848
rect 76374 23740 76380 23792
rect 76432 23780 76438 23792
rect 81728 23780 81756 23820
rect 84010 23808 84016 23820
rect 84068 23808 84074 23860
rect 76432 23752 81756 23780
rect 76432 23740 76438 23752
rect 83826 23740 83832 23792
rect 83884 23780 83890 23792
rect 95329 23783 95387 23789
rect 95329 23780 95341 23783
rect 83884 23752 95341 23780
rect 83884 23740 83890 23752
rect 95329 23749 95341 23752
rect 95375 23780 95387 23783
rect 95605 23783 95663 23789
rect 95605 23780 95617 23783
rect 95375 23752 95617 23780
rect 95375 23749 95387 23752
rect 95329 23743 95387 23749
rect 95605 23749 95617 23752
rect 95651 23780 95663 23783
rect 95789 23783 95847 23789
rect 95789 23780 95801 23783
rect 95651 23752 95801 23780
rect 95651 23749 95663 23752
rect 95605 23743 95663 23749
rect 95789 23749 95801 23752
rect 95835 23780 95847 23783
rect 95835 23752 96016 23780
rect 95835 23749 95847 23752
rect 95789 23743 95847 23749
rect 83550 23712 83556 23724
rect 76024 23684 83556 23712
rect 83550 23672 83556 23684
rect 83608 23672 83614 23724
rect 95988 23712 96016 23752
rect 96249 23715 96307 23721
rect 96249 23712 96261 23715
rect 95988 23684 96261 23712
rect 96249 23681 96261 23684
rect 96295 23712 96307 23715
rect 97721 23715 97779 23721
rect 97721 23712 97733 23715
rect 96295 23684 97733 23712
rect 96295 23681 96307 23684
rect 96249 23675 96307 23681
rect 97721 23681 97733 23684
rect 97767 23712 97779 23715
rect 97905 23715 97963 23721
rect 97905 23712 97917 23715
rect 97767 23684 97917 23712
rect 97767 23681 97779 23684
rect 97721 23675 97779 23681
rect 97905 23681 97917 23684
rect 97951 23712 97963 23715
rect 98089 23715 98147 23721
rect 98089 23712 98101 23715
rect 97951 23684 98101 23712
rect 97951 23681 97963 23684
rect 97905 23675 97963 23681
rect 98089 23681 98101 23684
rect 98135 23681 98147 23715
rect 98089 23675 98147 23681
rect 72513 23647 72571 23653
rect 72513 23613 72525 23647
rect 72559 23644 72571 23647
rect 73062 23644 73068 23656
rect 72559 23616 73068 23644
rect 72559 23613 72571 23616
rect 72513 23607 72571 23613
rect 73062 23604 73068 23616
rect 73120 23604 73126 23656
rect 74997 23647 75055 23653
rect 74997 23613 75009 23647
rect 75043 23644 75055 23647
rect 75086 23644 75092 23656
rect 75043 23616 75092 23644
rect 75043 23613 75055 23616
rect 74997 23607 75055 23613
rect 75086 23604 75092 23616
rect 75144 23604 75150 23656
rect 76745 23647 76803 23653
rect 76745 23644 76757 23647
rect 75380 23616 76757 23644
rect 65904 23548 72372 23576
rect 65797 23539 65855 23545
rect 74442 23536 74448 23588
rect 74500 23576 74506 23588
rect 75242 23579 75300 23585
rect 75242 23576 75254 23579
rect 74500 23548 75254 23576
rect 74500 23536 74506 23548
rect 75242 23545 75254 23548
rect 75288 23545 75300 23579
rect 75242 23539 75300 23545
rect 65886 23508 65892 23520
rect 65567 23480 65748 23508
rect 65847 23480 65892 23508
rect 65567 23477 65579 23480
rect 65521 23471 65579 23477
rect 65886 23468 65892 23480
rect 65944 23468 65950 23520
rect 74994 23468 75000 23520
rect 75052 23508 75058 23520
rect 75380 23508 75408 23616
rect 75052 23480 75408 23508
rect 75052 23468 75058 23480
rect 75454 23468 75460 23520
rect 75512 23508 75518 23520
rect 76006 23508 76012 23520
rect 75512 23480 76012 23508
rect 75512 23468 75518 23480
rect 76006 23468 76012 23480
rect 76064 23508 76070 23520
rect 76377 23511 76435 23517
rect 76377 23508 76389 23511
rect 76064 23480 76389 23508
rect 76064 23468 76070 23480
rect 76377 23477 76389 23480
rect 76423 23477 76435 23511
rect 76484 23508 76512 23616
rect 76745 23613 76757 23616
rect 76791 23613 76803 23647
rect 77110 23644 77116 23656
rect 77071 23616 77116 23644
rect 76745 23607 76803 23613
rect 77110 23604 77116 23616
rect 77168 23604 77174 23656
rect 77202 23604 77208 23656
rect 77260 23644 77266 23656
rect 77297 23647 77355 23653
rect 77297 23644 77309 23647
rect 77260 23616 77309 23644
rect 77260 23604 77266 23616
rect 77297 23613 77309 23616
rect 77343 23613 77355 23647
rect 77297 23607 77355 23613
rect 77389 23647 77447 23653
rect 77389 23613 77401 23647
rect 77435 23613 77447 23647
rect 77389 23607 77447 23613
rect 76558 23536 76564 23588
rect 76616 23576 76622 23588
rect 77220 23576 77248 23604
rect 76616 23548 77248 23576
rect 77404 23576 77432 23607
rect 78766 23604 78772 23656
rect 78824 23644 78830 23656
rect 79137 23647 79195 23653
rect 79137 23644 79149 23647
rect 78824 23616 79149 23644
rect 78824 23604 78830 23616
rect 79137 23613 79149 23616
rect 79183 23613 79195 23647
rect 79137 23607 79195 23613
rect 84930 23604 84936 23656
rect 84988 23644 84994 23656
rect 84988 23616 93854 23644
rect 84988 23604 84994 23616
rect 90174 23576 90180 23588
rect 77404 23548 90180 23576
rect 76616 23536 76622 23548
rect 77404 23508 77432 23548
rect 90174 23536 90180 23548
rect 90232 23536 90238 23588
rect 93826 23576 93854 23616
rect 94682 23604 94688 23656
rect 94740 23644 94746 23656
rect 95973 23647 96031 23653
rect 95973 23644 95985 23647
rect 94740 23616 95985 23644
rect 94740 23604 94746 23616
rect 95973 23613 95985 23616
rect 96019 23613 96031 23647
rect 95973 23607 96031 23613
rect 93826 23548 95924 23576
rect 76484 23480 77432 23508
rect 95896 23508 95924 23548
rect 97353 23511 97411 23517
rect 97353 23508 97365 23511
rect 95896 23480 97365 23508
rect 76377 23471 76435 23477
rect 97353 23477 97365 23480
rect 97399 23477 97411 23511
rect 97353 23471 97411 23477
rect 1104 23418 98808 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 50326 23418
rect 50378 23366 50390 23418
rect 50442 23366 50454 23418
rect 50506 23366 50518 23418
rect 50570 23366 81046 23418
rect 81098 23366 81110 23418
rect 81162 23366 81174 23418
rect 81226 23366 81238 23418
rect 81290 23366 98808 23418
rect 1104 23344 98808 23366
rect 1854 23264 1860 23316
rect 1912 23304 1918 23316
rect 6914 23304 6920 23316
rect 1912 23276 6920 23304
rect 1912 23264 1918 23276
rect 6914 23264 6920 23276
rect 6972 23264 6978 23316
rect 17218 23304 17224 23316
rect 7576 23276 17224 23304
rect 2314 23196 2320 23248
rect 2372 23236 2378 23248
rect 7576 23236 7604 23276
rect 17218 23264 17224 23276
rect 17276 23264 17282 23316
rect 25685 23307 25743 23313
rect 25685 23273 25697 23307
rect 25731 23304 25743 23307
rect 25866 23304 25872 23316
rect 25731 23276 25872 23304
rect 25731 23273 25743 23276
rect 25685 23267 25743 23273
rect 25866 23264 25872 23276
rect 25924 23264 25930 23316
rect 26142 23264 26148 23316
rect 26200 23304 26206 23316
rect 26513 23307 26571 23313
rect 26513 23304 26525 23307
rect 26200 23276 26525 23304
rect 26200 23264 26206 23276
rect 26513 23273 26525 23276
rect 26559 23273 26571 23307
rect 26513 23267 26571 23273
rect 29086 23264 29092 23316
rect 29144 23304 29150 23316
rect 29914 23304 29920 23316
rect 29144 23276 29920 23304
rect 29144 23264 29150 23276
rect 29914 23264 29920 23276
rect 29972 23264 29978 23316
rect 35986 23264 35992 23316
rect 36044 23304 36050 23316
rect 36538 23304 36544 23316
rect 36044 23276 36544 23304
rect 36044 23264 36050 23276
rect 36538 23264 36544 23276
rect 36596 23264 36602 23316
rect 37918 23264 37924 23316
rect 37976 23304 37982 23316
rect 48130 23304 48136 23316
rect 37976 23276 48136 23304
rect 37976 23264 37982 23276
rect 48130 23264 48136 23276
rect 48188 23264 48194 23316
rect 48498 23304 48504 23316
rect 48459 23276 48504 23304
rect 48498 23264 48504 23276
rect 48556 23264 48562 23316
rect 48866 23264 48872 23316
rect 48924 23304 48930 23316
rect 49510 23304 49516 23316
rect 48924 23276 49516 23304
rect 48924 23264 48930 23276
rect 49510 23264 49516 23276
rect 49568 23304 49574 23316
rect 56042 23304 56048 23316
rect 49568 23276 56048 23304
rect 49568 23264 49574 23276
rect 56042 23264 56048 23276
rect 56100 23264 56106 23316
rect 56226 23264 56232 23316
rect 56284 23304 56290 23316
rect 56284 23276 70394 23304
rect 56284 23264 56290 23276
rect 2372 23208 7604 23236
rect 11149 23239 11207 23245
rect 2372 23196 2378 23208
rect 11149 23205 11161 23239
rect 11195 23236 11207 23239
rect 11422 23236 11428 23248
rect 11195 23208 11428 23236
rect 11195 23205 11207 23208
rect 11149 23199 11207 23205
rect 11422 23196 11428 23208
rect 11480 23196 11486 23248
rect 14182 23196 14188 23248
rect 14240 23236 14246 23248
rect 39206 23236 39212 23248
rect 14240 23208 39212 23236
rect 14240 23196 14246 23208
rect 39206 23196 39212 23208
rect 39264 23236 39270 23248
rect 61841 23239 61899 23245
rect 61841 23236 61853 23239
rect 39264 23208 61853 23236
rect 39264 23196 39270 23208
rect 61841 23205 61853 23208
rect 61887 23236 61899 23239
rect 66162 23236 66168 23248
rect 61887 23208 66168 23236
rect 61887 23205 61899 23208
rect 61841 23199 61899 23205
rect 6914 23128 6920 23180
rect 6972 23168 6978 23180
rect 7558 23168 7564 23180
rect 6972 23140 7564 23168
rect 6972 23128 6978 23140
rect 7558 23128 7564 23140
rect 7616 23128 7622 23180
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 14734 23168 14740 23180
rect 9272 23140 14596 23168
rect 14695 23140 14740 23168
rect 9272 23128 9278 23140
rect 9398 23060 9404 23112
rect 9456 23100 9462 23112
rect 9493 23103 9551 23109
rect 9493 23100 9505 23103
rect 9456 23072 9505 23100
rect 9456 23060 9462 23072
rect 9493 23069 9505 23072
rect 9539 23069 9551 23103
rect 9766 23100 9772 23112
rect 9727 23072 9772 23100
rect 9493 23063 9551 23069
rect 9766 23060 9772 23072
rect 9824 23060 9830 23112
rect 14568 23032 14596 23140
rect 14734 23128 14740 23140
rect 14792 23128 14798 23180
rect 14918 23168 14924 23180
rect 14879 23140 14924 23168
rect 14918 23128 14924 23140
rect 14976 23128 14982 23180
rect 15013 23171 15071 23177
rect 15013 23137 15025 23171
rect 15059 23137 15071 23171
rect 15013 23131 15071 23137
rect 15105 23171 15163 23177
rect 15105 23137 15117 23171
rect 15151 23168 15163 23171
rect 15654 23168 15660 23180
rect 15151 23140 15660 23168
rect 15151 23137 15163 23140
rect 15105 23131 15163 23137
rect 15024 23032 15052 23131
rect 15654 23128 15660 23140
rect 15712 23168 15718 23180
rect 17034 23168 17040 23180
rect 15712 23140 17040 23168
rect 15712 23128 15718 23140
rect 17034 23128 17040 23140
rect 17092 23128 17098 23180
rect 25685 23171 25743 23177
rect 25685 23137 25697 23171
rect 25731 23168 25743 23171
rect 25777 23171 25835 23177
rect 25777 23168 25789 23171
rect 25731 23140 25789 23168
rect 25731 23137 25743 23140
rect 25685 23131 25743 23137
rect 25777 23137 25789 23140
rect 25823 23137 25835 23171
rect 25777 23131 25835 23137
rect 25961 23171 26019 23177
rect 25961 23137 25973 23171
rect 26007 23137 26019 23171
rect 25961 23131 26019 23137
rect 26191 23171 26249 23177
rect 26191 23137 26203 23171
rect 26237 23137 26249 23171
rect 26191 23131 26249 23137
rect 19886 23100 19892 23112
rect 15304 23072 19892 23100
rect 15194 23032 15200 23044
rect 10428 23004 12434 23032
rect 14568 23004 15200 23032
rect 4706 22924 4712 22976
rect 4764 22964 4770 22976
rect 10428 22964 10456 23004
rect 4764 22936 10456 22964
rect 12406 22964 12434 23004
rect 15194 22992 15200 23004
rect 15252 22992 15258 23044
rect 15304 23041 15332 23072
rect 19886 23060 19892 23072
rect 19944 23060 19950 23112
rect 25222 23060 25228 23112
rect 25280 23100 25286 23112
rect 25976 23100 26004 23131
rect 25280 23072 26004 23100
rect 25280 23060 25286 23072
rect 26050 23060 26056 23112
rect 26108 23100 26114 23112
rect 26206 23100 26234 23131
rect 26326 23128 26332 23180
rect 26384 23168 26390 23180
rect 26510 23168 26516 23180
rect 26384 23140 26516 23168
rect 26384 23128 26390 23140
rect 26510 23128 26516 23140
rect 26568 23128 26574 23180
rect 33134 23168 33140 23180
rect 26804 23140 33140 23168
rect 26804 23100 26832 23140
rect 33134 23128 33140 23140
rect 33192 23168 33198 23180
rect 35618 23168 35624 23180
rect 33192 23140 35624 23168
rect 33192 23128 33198 23140
rect 35618 23128 35624 23140
rect 35676 23128 35682 23180
rect 44174 23128 44180 23180
rect 44232 23168 44238 23180
rect 44542 23168 44548 23180
rect 44232 23140 44548 23168
rect 44232 23128 44238 23140
rect 44542 23128 44548 23140
rect 44600 23128 44606 23180
rect 47486 23168 47492 23180
rect 47447 23140 47492 23168
rect 47486 23128 47492 23140
rect 47544 23168 47550 23180
rect 48406 23168 48412 23180
rect 47544 23140 48412 23168
rect 47544 23128 47550 23140
rect 48406 23128 48412 23140
rect 48464 23128 48470 23180
rect 48682 23128 48688 23180
rect 48740 23168 48746 23180
rect 49050 23168 49056 23180
rect 48740 23140 49056 23168
rect 48740 23128 48746 23140
rect 49050 23128 49056 23140
rect 49108 23128 49114 23180
rect 49142 23128 49148 23180
rect 49200 23168 49206 23180
rect 53742 23168 53748 23180
rect 49200 23140 53748 23168
rect 49200 23128 49206 23140
rect 53742 23128 53748 23140
rect 53800 23128 53806 23180
rect 53834 23128 53840 23180
rect 53892 23168 53898 23180
rect 56134 23168 56140 23180
rect 53892 23140 56140 23168
rect 53892 23128 53898 23140
rect 56134 23128 56140 23140
rect 56192 23128 56198 23180
rect 61948 23177 61976 23208
rect 66162 23196 66168 23208
rect 66220 23196 66226 23248
rect 61933 23171 61991 23177
rect 61933 23137 61945 23171
rect 61979 23168 61991 23171
rect 62114 23168 62120 23180
rect 61979 23140 62013 23168
rect 62075 23140 62120 23168
rect 61979 23137 61991 23140
rect 61933 23131 61991 23137
rect 62114 23128 62120 23140
rect 62172 23128 62178 23180
rect 62482 23128 62488 23180
rect 62540 23168 62546 23180
rect 62540 23140 62585 23168
rect 62540 23128 62546 23140
rect 64690 23128 64696 23180
rect 64748 23168 64754 23180
rect 70121 23171 70179 23177
rect 70121 23168 70133 23171
rect 64748 23140 70133 23168
rect 64748 23128 64754 23140
rect 70121 23137 70133 23140
rect 70167 23137 70179 23171
rect 70366 23168 70394 23276
rect 72234 23264 72240 23316
rect 72292 23304 72298 23316
rect 73249 23307 73307 23313
rect 73249 23304 73261 23307
rect 72292 23276 73261 23304
rect 72292 23264 72298 23276
rect 73249 23273 73261 23276
rect 73295 23273 73307 23307
rect 73249 23267 73307 23273
rect 75454 23264 75460 23316
rect 75512 23304 75518 23316
rect 76374 23304 76380 23316
rect 75512 23276 76380 23304
rect 75512 23264 75518 23276
rect 76374 23264 76380 23276
rect 76432 23264 76438 23316
rect 76742 23264 76748 23316
rect 76800 23304 76806 23316
rect 88242 23304 88248 23316
rect 76800 23276 88248 23304
rect 76800 23264 76806 23276
rect 88242 23264 88248 23276
rect 88300 23264 88306 23316
rect 72142 23196 72148 23248
rect 72200 23236 72206 23248
rect 72421 23239 72479 23245
rect 72421 23236 72433 23239
rect 72200 23208 72433 23236
rect 72200 23196 72206 23208
rect 72421 23205 72433 23208
rect 72467 23236 72479 23239
rect 72467 23208 73016 23236
rect 72467 23205 72479 23208
rect 72421 23199 72479 23205
rect 70673 23171 70731 23177
rect 70673 23168 70685 23171
rect 70366 23140 70685 23168
rect 70121 23131 70179 23137
rect 70673 23137 70685 23140
rect 70719 23168 70731 23171
rect 72050 23168 72056 23180
rect 70719 23140 72056 23168
rect 70719 23137 70731 23140
rect 70673 23131 70731 23137
rect 72050 23128 72056 23140
rect 72108 23128 72114 23180
rect 72602 23168 72608 23180
rect 72563 23140 72608 23168
rect 72602 23128 72608 23140
rect 72660 23128 72666 23180
rect 72694 23128 72700 23180
rect 72752 23177 72758 23180
rect 72988 23177 73016 23208
rect 76650 23196 76656 23248
rect 76708 23236 76714 23248
rect 90082 23236 90088 23248
rect 76708 23208 90088 23236
rect 76708 23196 76714 23208
rect 90082 23196 90088 23208
rect 90140 23196 90146 23248
rect 72752 23171 72811 23177
rect 72752 23137 72765 23171
rect 72799 23137 72811 23171
rect 72752 23131 72811 23137
rect 72973 23171 73031 23177
rect 72973 23137 72985 23171
rect 73019 23137 73031 23171
rect 72973 23131 73031 23137
rect 73157 23171 73215 23177
rect 73157 23137 73169 23171
rect 73203 23137 73215 23171
rect 73157 23131 73215 23137
rect 72752 23128 72758 23131
rect 26108 23072 26153 23100
rect 26206 23072 26832 23100
rect 26108 23060 26114 23072
rect 26206 23044 26234 23072
rect 26878 23060 26884 23112
rect 26936 23100 26942 23112
rect 46842 23100 46848 23112
rect 26936 23072 46848 23100
rect 26936 23060 26942 23072
rect 46842 23060 46848 23072
rect 46900 23060 46906 23112
rect 47670 23100 47676 23112
rect 47631 23072 47676 23100
rect 47670 23060 47676 23072
rect 47728 23060 47734 23112
rect 48038 23100 48044 23112
rect 47999 23072 48044 23100
rect 48038 23060 48044 23072
rect 48096 23060 48102 23112
rect 48130 23060 48136 23112
rect 48188 23100 48194 23112
rect 55490 23100 55496 23112
rect 48188 23072 55496 23100
rect 48188 23060 48194 23072
rect 55490 23060 55496 23072
rect 55548 23060 55554 23112
rect 55674 23060 55680 23112
rect 55732 23100 55738 23112
rect 61010 23100 61016 23112
rect 55732 23072 61016 23100
rect 55732 23060 55738 23072
rect 61010 23060 61016 23072
rect 61068 23060 61074 23112
rect 62206 23100 62212 23112
rect 62167 23072 62212 23100
rect 62206 23060 62212 23072
rect 62264 23060 62270 23112
rect 62301 23103 62359 23109
rect 62301 23069 62313 23103
rect 62347 23100 62359 23103
rect 62574 23100 62580 23112
rect 62347 23072 62580 23100
rect 62347 23069 62359 23072
rect 62301 23063 62359 23069
rect 15289 23035 15347 23041
rect 15289 23001 15301 23035
rect 15335 23001 15347 23035
rect 15289 22995 15347 23001
rect 17310 22992 17316 23044
rect 17368 23032 17374 23044
rect 25314 23032 25320 23044
rect 17368 23004 25320 23032
rect 17368 22992 17374 23004
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 26142 22992 26148 23044
rect 26200 23004 26234 23044
rect 47302 23032 47308 23044
rect 26344 23004 47308 23032
rect 26200 22992 26206 23004
rect 26344 22964 26372 23004
rect 47302 22992 47308 23004
rect 47360 22992 47366 23044
rect 48685 23035 48743 23041
rect 48685 23032 48697 23035
rect 47688 23004 48697 23032
rect 12406 22936 26372 22964
rect 4764 22924 4770 22936
rect 26878 22924 26884 22976
rect 26936 22964 26942 22976
rect 33134 22964 33140 22976
rect 26936 22936 33140 22964
rect 26936 22924 26942 22936
rect 33134 22924 33140 22936
rect 33192 22964 33198 22976
rect 37734 22964 37740 22976
rect 33192 22936 37740 22964
rect 33192 22924 33198 22936
rect 37734 22924 37740 22936
rect 37792 22924 37798 22976
rect 46014 22924 46020 22976
rect 46072 22964 46078 22976
rect 46382 22964 46388 22976
rect 46072 22936 46388 22964
rect 46072 22924 46078 22936
rect 46382 22924 46388 22936
rect 46440 22924 46446 22976
rect 46842 22924 46848 22976
rect 46900 22964 46906 22976
rect 47688 22964 47716 23004
rect 48148 22973 48176 23004
rect 48685 23001 48697 23004
rect 48731 23032 48743 23035
rect 49326 23032 49332 23044
rect 48731 23004 49332 23032
rect 48731 23001 48743 23004
rect 48685 22995 48743 23001
rect 49326 22992 49332 23004
rect 49384 22992 49390 23044
rect 49786 22992 49792 23044
rect 49844 23032 49850 23044
rect 62316 23032 62344 23063
rect 62574 23060 62580 23072
rect 62632 23060 62638 23112
rect 67174 23060 67180 23112
rect 67232 23100 67238 23112
rect 67450 23100 67456 23112
rect 67232 23072 67456 23100
rect 67232 23060 67238 23072
rect 67450 23060 67456 23072
rect 67508 23060 67514 23112
rect 67634 23060 67640 23112
rect 67692 23100 67698 23112
rect 67729 23103 67787 23109
rect 67729 23100 67741 23103
rect 67692 23072 67741 23100
rect 67692 23060 67698 23072
rect 67729 23069 67741 23072
rect 67775 23069 67787 23103
rect 67729 23063 67787 23069
rect 71958 23060 71964 23112
rect 72016 23100 72022 23112
rect 72881 23103 72939 23109
rect 72881 23100 72893 23103
rect 72016 23072 72893 23100
rect 72016 23060 72022 23072
rect 72881 23069 72893 23072
rect 72927 23069 72939 23103
rect 72881 23063 72939 23069
rect 49844 23004 62344 23032
rect 49844 22992 49850 23004
rect 62850 22992 62856 23044
rect 62908 23032 62914 23044
rect 63678 23032 63684 23044
rect 62908 23004 63684 23032
rect 62908 22992 62914 23004
rect 63678 22992 63684 23004
rect 63736 22992 63742 23044
rect 64414 22992 64420 23044
rect 64472 23032 64478 23044
rect 66530 23032 66536 23044
rect 64472 23004 66536 23032
rect 64472 22992 64478 23004
rect 66530 22992 66536 23004
rect 66588 22992 66594 23044
rect 71038 23032 71044 23044
rect 68388 23004 71044 23032
rect 46900 22936 47716 22964
rect 48133 22967 48191 22973
rect 46900 22924 46906 22936
rect 48133 22933 48145 22967
rect 48179 22964 48191 22967
rect 48271 22967 48329 22973
rect 48179 22936 48213 22964
rect 48179 22933 48191 22936
rect 48133 22927 48191 22933
rect 48271 22933 48283 22967
rect 48317 22964 48329 22967
rect 48498 22964 48504 22976
rect 48317 22936 48504 22964
rect 48317 22933 48329 22936
rect 48271 22927 48329 22933
rect 48498 22924 48504 22936
rect 48556 22924 48562 22976
rect 48774 22924 48780 22976
rect 48832 22964 48838 22976
rect 53834 22964 53840 22976
rect 48832 22936 53840 22964
rect 48832 22924 48838 22936
rect 53834 22924 53840 22936
rect 53892 22924 53898 22976
rect 53926 22924 53932 22976
rect 53984 22964 53990 22976
rect 55122 22964 55128 22976
rect 53984 22936 55128 22964
rect 53984 22924 53990 22936
rect 55122 22924 55128 22936
rect 55180 22924 55186 22976
rect 55490 22924 55496 22976
rect 55548 22964 55554 22976
rect 56226 22964 56232 22976
rect 55548 22936 56232 22964
rect 55548 22924 55554 22936
rect 56226 22924 56232 22936
rect 56284 22924 56290 22976
rect 62669 22967 62727 22973
rect 62669 22933 62681 22967
rect 62715 22964 62727 22967
rect 62758 22964 62764 22976
rect 62715 22936 62764 22964
rect 62715 22933 62727 22936
rect 62669 22927 62727 22933
rect 62758 22924 62764 22936
rect 62816 22924 62822 22976
rect 65242 22924 65248 22976
rect 65300 22964 65306 22976
rect 68388 22964 68416 23004
rect 71038 22992 71044 23004
rect 71096 23032 71102 23044
rect 71682 23032 71688 23044
rect 71096 23004 71688 23032
rect 71096 22992 71102 23004
rect 71682 22992 71688 23004
rect 71740 22992 71746 23044
rect 72234 22992 72240 23044
rect 72292 23032 72298 23044
rect 72418 23032 72424 23044
rect 72292 23004 72424 23032
rect 72292 22992 72298 23004
rect 72418 22992 72424 23004
rect 72476 22992 72482 23044
rect 65300 22936 68416 22964
rect 69017 22967 69075 22973
rect 65300 22924 65306 22936
rect 69017 22933 69029 22967
rect 69063 22964 69075 22967
rect 69106 22964 69112 22976
rect 69063 22936 69112 22964
rect 69063 22933 69075 22936
rect 69017 22927 69075 22933
rect 69106 22924 69112 22936
rect 69164 22924 69170 22976
rect 70486 22924 70492 22976
rect 70544 22964 70550 22976
rect 73172 22964 73200 23131
rect 81894 23128 81900 23180
rect 81952 23168 81958 23180
rect 89346 23168 89352 23180
rect 81952 23140 89352 23168
rect 81952 23128 81958 23140
rect 89346 23128 89352 23140
rect 89404 23128 89410 23180
rect 73430 23060 73436 23112
rect 73488 23060 73494 23112
rect 74350 23060 74356 23112
rect 74408 23100 74414 23112
rect 91094 23100 91100 23112
rect 74408 23072 91100 23100
rect 74408 23060 74414 23072
rect 91094 23060 91100 23072
rect 91152 23060 91158 23112
rect 73448 23032 73476 23060
rect 93394 23032 93400 23044
rect 73448 23004 93400 23032
rect 93394 22992 93400 23004
rect 93452 22992 93458 23044
rect 73433 22967 73491 22973
rect 73433 22964 73445 22967
rect 70544 22936 73445 22964
rect 70544 22924 70550 22936
rect 73433 22933 73445 22936
rect 73479 22933 73491 22967
rect 73433 22927 73491 22933
rect 74442 22924 74448 22976
rect 74500 22964 74506 22976
rect 78766 22964 78772 22976
rect 74500 22936 78772 22964
rect 74500 22924 74506 22936
rect 78766 22924 78772 22936
rect 78824 22924 78830 22976
rect 1104 22874 98808 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 65686 22874
rect 65738 22822 65750 22874
rect 65802 22822 65814 22874
rect 65866 22822 65878 22874
rect 65930 22822 96406 22874
rect 96458 22822 96470 22874
rect 96522 22822 96534 22874
rect 96586 22822 96598 22874
rect 96650 22822 98808 22874
rect 1104 22800 98808 22822
rect 14645 22763 14703 22769
rect 14645 22729 14657 22763
rect 14691 22760 14703 22763
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 14691 22732 14933 22760
rect 14691 22729 14703 22732
rect 14645 22723 14703 22729
rect 14921 22729 14933 22732
rect 14967 22760 14979 22763
rect 15010 22760 15016 22772
rect 14967 22732 15016 22760
rect 14967 22729 14979 22732
rect 14921 22723 14979 22729
rect 15010 22720 15016 22732
rect 15068 22720 15074 22772
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 26326 22760 26332 22772
rect 17276 22732 26332 22760
rect 17276 22720 17282 22732
rect 26326 22720 26332 22732
rect 26384 22720 26390 22772
rect 37734 22720 37740 22772
rect 37792 22760 37798 22772
rect 47670 22760 47676 22772
rect 37792 22732 47676 22760
rect 37792 22720 37798 22732
rect 47670 22720 47676 22732
rect 47728 22720 47734 22772
rect 48314 22720 48320 22772
rect 48372 22760 48378 22772
rect 48498 22760 48504 22772
rect 48372 22732 48504 22760
rect 48372 22720 48378 22732
rect 48498 22720 48504 22732
rect 48556 22720 48562 22772
rect 49878 22720 49884 22772
rect 49936 22760 49942 22772
rect 55674 22760 55680 22772
rect 49936 22732 55680 22760
rect 49936 22720 49942 22732
rect 55674 22720 55680 22732
rect 55732 22720 55738 22772
rect 56042 22720 56048 22772
rect 56100 22760 56106 22772
rect 56100 22732 65564 22760
rect 56100 22720 56106 22732
rect 2038 22652 2044 22704
rect 2096 22692 2102 22704
rect 15102 22692 15108 22704
rect 2096 22664 15108 22692
rect 2096 22652 2102 22664
rect 15102 22652 15108 22664
rect 15160 22652 15166 22704
rect 15194 22652 15200 22704
rect 15252 22692 15258 22704
rect 27154 22692 27160 22704
rect 15252 22664 27160 22692
rect 15252 22652 15258 22664
rect 27154 22652 27160 22664
rect 27212 22652 27218 22704
rect 33410 22652 33416 22704
rect 33468 22692 33474 22704
rect 33468 22664 33732 22692
rect 33468 22652 33474 22664
rect 11238 22584 11244 22636
rect 11296 22624 11302 22636
rect 11698 22624 11704 22636
rect 11296 22596 11704 22624
rect 11296 22584 11302 22596
rect 11698 22584 11704 22596
rect 11756 22624 11762 22636
rect 17310 22624 17316 22636
rect 11756 22596 17316 22624
rect 11756 22584 11762 22596
rect 17310 22584 17316 22596
rect 17368 22584 17374 22636
rect 23750 22584 23756 22636
rect 23808 22624 23814 22636
rect 33594 22624 33600 22636
rect 23808 22596 33600 22624
rect 23808 22584 23814 22596
rect 33594 22584 33600 22596
rect 33652 22584 33658 22636
rect 33704 22633 33732 22664
rect 36446 22652 36452 22704
rect 36504 22692 36510 22704
rect 64782 22692 64788 22704
rect 36504 22664 64788 22692
rect 36504 22652 36510 22664
rect 64782 22652 64788 22664
rect 64840 22652 64846 22704
rect 65426 22692 65432 22704
rect 64984 22664 65432 22692
rect 64984 22636 65012 22664
rect 65426 22652 65432 22664
rect 65484 22652 65490 22704
rect 33689 22627 33747 22633
rect 33689 22593 33701 22627
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 33870 22584 33876 22636
rect 33928 22624 33934 22636
rect 64414 22624 64420 22636
rect 33928 22596 64420 22624
rect 33928 22584 33934 22596
rect 64414 22584 64420 22596
rect 64472 22584 64478 22636
rect 64966 22624 64972 22636
rect 64927 22596 64972 22624
rect 64966 22584 64972 22596
rect 65024 22584 65030 22636
rect 65058 22584 65064 22636
rect 65116 22624 65122 22636
rect 65536 22633 65564 22732
rect 71406 22720 71412 22772
rect 71464 22760 71470 22772
rect 95786 22760 95792 22772
rect 71464 22732 95792 22760
rect 71464 22720 71470 22732
rect 95786 22720 95792 22732
rect 95844 22720 95850 22772
rect 65889 22695 65947 22701
rect 65889 22661 65901 22695
rect 65935 22692 65947 22695
rect 73798 22692 73804 22704
rect 65935 22664 73804 22692
rect 65935 22661 65947 22664
rect 65889 22655 65947 22661
rect 73798 22652 73804 22664
rect 73856 22652 73862 22704
rect 65521 22627 65579 22633
rect 65116 22596 65380 22624
rect 65116 22584 65122 22596
rect 12986 22516 12992 22568
rect 13044 22556 13050 22568
rect 33505 22559 33563 22565
rect 33505 22556 33517 22559
rect 13044 22528 33517 22556
rect 13044 22516 13050 22528
rect 33505 22525 33517 22528
rect 33551 22556 33563 22559
rect 33965 22559 34023 22565
rect 33965 22556 33977 22559
rect 33551 22528 33977 22556
rect 33551 22525 33563 22528
rect 33505 22519 33563 22525
rect 33965 22525 33977 22528
rect 34011 22525 34023 22559
rect 33965 22519 34023 22525
rect 43990 22516 43996 22568
rect 44048 22556 44054 22568
rect 55306 22556 55312 22568
rect 44048 22528 55312 22556
rect 44048 22516 44054 22528
rect 55306 22516 55312 22528
rect 55364 22516 55370 22568
rect 58802 22516 58808 22568
rect 58860 22556 58866 22568
rect 62666 22556 62672 22568
rect 58860 22528 62672 22556
rect 58860 22516 58866 22528
rect 62666 22516 62672 22528
rect 62724 22516 62730 22568
rect 63126 22516 63132 22568
rect 63184 22556 63190 22568
rect 65153 22559 65211 22565
rect 65153 22556 65165 22559
rect 63184 22528 65165 22556
rect 63184 22516 63190 22528
rect 65153 22525 65165 22528
rect 65199 22556 65211 22559
rect 65242 22556 65248 22568
rect 65199 22528 65248 22556
rect 65199 22525 65211 22528
rect 65153 22519 65211 22525
rect 65242 22516 65248 22528
rect 65300 22516 65306 22568
rect 65352 22565 65380 22596
rect 65521 22593 65533 22627
rect 65567 22624 65579 22627
rect 65567 22596 65840 22624
rect 65567 22593 65579 22596
rect 65521 22587 65579 22593
rect 65337 22559 65395 22565
rect 65337 22525 65349 22559
rect 65383 22525 65395 22559
rect 65337 22519 65395 22525
rect 65426 22516 65432 22568
rect 65484 22556 65490 22568
rect 65702 22556 65708 22568
rect 65484 22528 65529 22556
rect 65663 22528 65708 22556
rect 65484 22516 65490 22528
rect 65702 22516 65708 22528
rect 65760 22516 65766 22568
rect 65812 22556 65840 22596
rect 66530 22584 66536 22636
rect 66588 22624 66594 22636
rect 74442 22624 74448 22636
rect 66588 22596 74448 22624
rect 66588 22584 66594 22596
rect 74442 22584 74448 22596
rect 74500 22584 74506 22636
rect 75454 22624 75460 22636
rect 74552 22596 75460 22624
rect 74552 22556 74580 22596
rect 75454 22584 75460 22596
rect 75512 22584 75518 22636
rect 65812 22528 74580 22556
rect 74626 22516 74632 22568
rect 74684 22556 74690 22568
rect 74997 22559 75055 22565
rect 74997 22556 75009 22559
rect 74684 22528 75009 22556
rect 74684 22516 74690 22528
rect 74997 22525 75009 22528
rect 75043 22556 75055 22559
rect 75546 22556 75552 22568
rect 75043 22528 75552 22556
rect 75043 22525 75055 22528
rect 74997 22519 75055 22525
rect 75546 22516 75552 22528
rect 75604 22516 75610 22568
rect 76098 22556 76104 22568
rect 76059 22528 76104 22556
rect 76098 22516 76104 22528
rect 76156 22516 76162 22568
rect 12710 22448 12716 22500
rect 12768 22488 12774 22500
rect 15102 22488 15108 22500
rect 12768 22460 15108 22488
rect 12768 22448 12774 22460
rect 15102 22448 15108 22460
rect 15160 22488 15166 22500
rect 15654 22488 15660 22500
rect 15160 22460 15660 22488
rect 15160 22448 15166 22460
rect 15654 22448 15660 22460
rect 15712 22448 15718 22500
rect 19242 22448 19248 22500
rect 19300 22488 19306 22500
rect 25222 22488 25228 22500
rect 19300 22460 25228 22488
rect 19300 22448 19306 22460
rect 25222 22448 25228 22460
rect 25280 22488 25286 22500
rect 25280 22460 33824 22488
rect 25280 22448 25286 22460
rect 16482 22380 16488 22432
rect 16540 22420 16546 22432
rect 33410 22420 33416 22432
rect 16540 22392 33416 22420
rect 16540 22380 16546 22392
rect 33410 22380 33416 22392
rect 33468 22380 33474 22432
rect 33796 22420 33824 22460
rect 34624 22460 64828 22488
rect 34624 22420 34652 22460
rect 35250 22420 35256 22432
rect 33796 22392 34652 22420
rect 35163 22392 35256 22420
rect 35250 22380 35256 22392
rect 35308 22420 35314 22432
rect 48774 22420 48780 22432
rect 35308 22392 48780 22420
rect 35308 22380 35314 22392
rect 48774 22380 48780 22392
rect 48832 22380 48838 22432
rect 50706 22380 50712 22432
rect 50764 22420 50770 22432
rect 54662 22420 54668 22432
rect 50764 22392 54668 22420
rect 50764 22380 50770 22392
rect 54662 22380 54668 22392
rect 54720 22380 54726 22432
rect 55122 22380 55128 22432
rect 55180 22420 55186 22432
rect 64690 22420 64696 22432
rect 55180 22392 64696 22420
rect 55180 22380 55186 22392
rect 64690 22380 64696 22392
rect 64748 22380 64754 22432
rect 64800 22420 64828 22460
rect 65058 22448 65064 22500
rect 65116 22488 65122 22500
rect 75273 22491 75331 22497
rect 75273 22488 75285 22491
rect 65116 22460 75285 22488
rect 65116 22448 65122 22460
rect 75273 22457 75285 22460
rect 75319 22457 75331 22491
rect 96890 22488 96896 22500
rect 75273 22451 75331 22457
rect 80026 22460 96896 22488
rect 80026 22420 80054 22460
rect 96890 22448 96896 22460
rect 96948 22448 96954 22500
rect 64800 22392 80054 22420
rect 1104 22330 98808 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 50326 22330
rect 50378 22278 50390 22330
rect 50442 22278 50454 22330
rect 50506 22278 50518 22330
rect 50570 22278 81046 22330
rect 81098 22278 81110 22330
rect 81162 22278 81174 22330
rect 81226 22278 81238 22330
rect 81290 22278 98808 22330
rect 1104 22256 98808 22278
rect 20438 22176 20444 22228
rect 20496 22216 20502 22228
rect 26878 22216 26884 22228
rect 20496 22188 26884 22216
rect 20496 22176 20502 22188
rect 26878 22176 26884 22188
rect 26936 22176 26942 22228
rect 29914 22176 29920 22228
rect 29972 22216 29978 22228
rect 29972 22188 33364 22216
rect 29972 22176 29978 22188
rect 11422 22108 11428 22160
rect 11480 22148 11486 22160
rect 13538 22148 13544 22160
rect 11480 22120 13544 22148
rect 11480 22108 11486 22120
rect 13538 22108 13544 22120
rect 13596 22108 13602 22160
rect 21082 22108 21088 22160
rect 21140 22148 21146 22160
rect 25590 22148 25596 22160
rect 21140 22120 25596 22148
rect 21140 22108 21146 22120
rect 25590 22108 25596 22120
rect 25648 22108 25654 22160
rect 26234 22148 26240 22160
rect 26206 22108 26240 22148
rect 26292 22148 26298 22160
rect 33042 22148 33048 22160
rect 26292 22120 33048 22148
rect 26292 22108 26298 22120
rect 33042 22108 33048 22120
rect 33100 22108 33106 22160
rect 33336 22148 33364 22188
rect 33410 22176 33416 22228
rect 33468 22216 33474 22228
rect 35250 22216 35256 22228
rect 33468 22188 35256 22216
rect 33468 22176 33474 22188
rect 35250 22176 35256 22188
rect 35308 22176 35314 22228
rect 38562 22176 38568 22228
rect 38620 22216 38626 22228
rect 95878 22216 95884 22228
rect 38620 22188 95884 22216
rect 38620 22176 38626 22188
rect 95878 22176 95884 22188
rect 95936 22176 95942 22228
rect 36446 22148 36452 22160
rect 33336 22120 36452 22148
rect 36446 22108 36452 22120
rect 36504 22108 36510 22160
rect 37642 22108 37648 22160
rect 37700 22148 37706 22160
rect 38377 22151 38435 22157
rect 38377 22148 38389 22151
rect 37700 22120 38389 22148
rect 37700 22108 37706 22120
rect 38377 22117 38389 22120
rect 38423 22117 38435 22151
rect 46842 22148 46848 22160
rect 38377 22111 38435 22117
rect 39960 22120 46848 22148
rect 9858 22080 9864 22092
rect 9819 22052 9864 22080
rect 9858 22040 9864 22052
rect 9916 22040 9922 22092
rect 17310 22040 17316 22092
rect 17368 22080 17374 22092
rect 26206 22080 26234 22108
rect 17368 22052 26234 22080
rect 17368 22040 17374 22052
rect 30190 22040 30196 22092
rect 30248 22080 30254 22092
rect 38105 22083 38163 22089
rect 38105 22080 38117 22083
rect 30248 22052 38117 22080
rect 30248 22040 30254 22052
rect 38105 22049 38117 22052
rect 38151 22080 38163 22083
rect 38194 22080 38200 22092
rect 38151 22052 38200 22080
rect 38151 22049 38163 22052
rect 38105 22043 38163 22049
rect 38194 22040 38200 22052
rect 38252 22040 38258 22092
rect 38289 22083 38347 22089
rect 38289 22049 38301 22083
rect 38335 22049 38347 22083
rect 38470 22080 38476 22092
rect 38383 22052 38476 22080
rect 38289 22043 38347 22049
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 22012 10471 22015
rect 17126 22012 17132 22024
rect 10459 21984 17132 22012
rect 10459 21981 10471 21984
rect 10413 21975 10471 21981
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 24118 21972 24124 22024
rect 24176 22012 24182 22024
rect 38304 22012 38332 22043
rect 38470 22040 38476 22052
rect 38528 22080 38534 22092
rect 39960 22080 39988 22120
rect 46842 22108 46848 22120
rect 46900 22108 46906 22160
rect 52362 22108 52368 22160
rect 52420 22148 52426 22160
rect 52457 22151 52515 22157
rect 52457 22148 52469 22151
rect 52420 22120 52469 22148
rect 52420 22108 52426 22120
rect 52457 22117 52469 22120
rect 52503 22117 52515 22151
rect 52457 22111 52515 22117
rect 54662 22108 54668 22160
rect 54720 22148 54726 22160
rect 64598 22148 64604 22160
rect 54720 22120 64604 22148
rect 54720 22108 54726 22120
rect 64598 22108 64604 22120
rect 64656 22108 64662 22160
rect 64782 22108 64788 22160
rect 64840 22148 64846 22160
rect 70486 22148 70492 22160
rect 64840 22120 70492 22148
rect 64840 22108 64846 22120
rect 70486 22108 70492 22120
rect 70544 22108 70550 22160
rect 38528 22052 39988 22080
rect 38528 22040 38534 22052
rect 40034 22040 40040 22092
rect 40092 22080 40098 22092
rect 40494 22080 40500 22092
rect 40092 22052 40500 22080
rect 40092 22040 40098 22052
rect 40494 22040 40500 22052
rect 40552 22080 40558 22092
rect 43533 22083 43591 22089
rect 43533 22080 43545 22083
rect 40552 22052 43545 22080
rect 40552 22040 40558 22052
rect 43533 22049 43545 22052
rect 43579 22049 43591 22083
rect 43533 22043 43591 22049
rect 43625 22083 43683 22089
rect 43625 22049 43637 22083
rect 43671 22049 43683 22083
rect 43806 22080 43812 22092
rect 43767 22052 43812 22080
rect 43625 22043 43683 22049
rect 42150 22012 42156 22024
rect 24176 21984 38332 22012
rect 38488 21984 42156 22012
rect 24176 21972 24182 21984
rect 25590 21904 25596 21956
rect 25648 21944 25654 21956
rect 28994 21944 29000 21956
rect 25648 21916 29000 21944
rect 25648 21904 25654 21916
rect 28994 21904 29000 21916
rect 29052 21904 29058 21956
rect 38378 21904 38384 21956
rect 38436 21944 38442 21956
rect 38488 21944 38516 21984
rect 42150 21972 42156 21984
rect 42208 21972 42214 22024
rect 43441 21947 43499 21953
rect 38436 21916 38516 21944
rect 38580 21916 41644 21944
rect 38436 21904 38442 21916
rect 6178 21836 6184 21888
rect 6236 21876 6242 21888
rect 37918 21876 37924 21888
rect 6236 21848 37924 21876
rect 6236 21836 6242 21848
rect 37918 21836 37924 21848
rect 37976 21836 37982 21888
rect 38013 21879 38071 21885
rect 38013 21845 38025 21879
rect 38059 21876 38071 21879
rect 38194 21876 38200 21888
rect 38059 21848 38200 21876
rect 38059 21845 38071 21848
rect 38013 21839 38071 21845
rect 38194 21836 38200 21848
rect 38252 21876 38258 21888
rect 38580 21876 38608 21916
rect 38252 21848 38608 21876
rect 38657 21879 38715 21885
rect 38252 21836 38258 21848
rect 38657 21845 38669 21879
rect 38703 21876 38715 21879
rect 41506 21876 41512 21888
rect 38703 21848 41512 21876
rect 38703 21845 38715 21848
rect 38657 21839 38715 21845
rect 41506 21836 41512 21848
rect 41564 21836 41570 21888
rect 41616 21876 41644 21916
rect 43441 21913 43453 21947
rect 43487 21944 43499 21947
rect 43640 21944 43668 22043
rect 43806 22040 43812 22052
rect 43864 22040 43870 22092
rect 46750 22040 46756 22092
rect 46808 22080 46814 22092
rect 52181 22083 52239 22089
rect 52181 22080 52193 22083
rect 46808 22052 52193 22080
rect 46808 22040 46814 22052
rect 52181 22049 52193 22052
rect 52227 22080 52239 22083
rect 52638 22080 52644 22092
rect 52227 22052 52644 22080
rect 52227 22049 52239 22052
rect 52181 22043 52239 22049
rect 52638 22040 52644 22052
rect 52696 22040 52702 22092
rect 55490 22040 55496 22092
rect 55548 22080 55554 22092
rect 55766 22080 55772 22092
rect 55548 22052 55772 22080
rect 55548 22040 55554 22052
rect 55766 22040 55772 22052
rect 55824 22040 55830 22092
rect 73430 22080 73436 22092
rect 55876 22052 73436 22080
rect 43993 22015 44051 22021
rect 43993 21981 44005 22015
rect 44039 22012 44051 22015
rect 46198 22012 46204 22024
rect 44039 21984 46204 22012
rect 44039 21981 44051 21984
rect 43993 21975 44051 21981
rect 46198 21972 46204 21984
rect 46256 21972 46262 22024
rect 46290 21972 46296 22024
rect 46348 22012 46354 22024
rect 51718 22012 51724 22024
rect 46348 21984 51724 22012
rect 46348 21972 46354 21984
rect 51718 21972 51724 21984
rect 51776 21972 51782 22024
rect 53098 21972 53104 22024
rect 53156 22012 53162 22024
rect 55876 22012 55904 22052
rect 73430 22040 73436 22052
rect 73488 22040 73494 22092
rect 75362 22080 75368 22092
rect 75323 22052 75368 22080
rect 75362 22040 75368 22052
rect 75420 22040 75426 22092
rect 75914 22040 75920 22092
rect 75972 22080 75978 22092
rect 85025 22083 85083 22089
rect 85025 22080 85037 22083
rect 75972 22052 85037 22080
rect 75972 22040 75978 22052
rect 85025 22049 85037 22052
rect 85071 22049 85083 22083
rect 85393 22083 85451 22089
rect 85393 22080 85405 22083
rect 85025 22043 85083 22049
rect 85132 22052 85405 22080
rect 76006 22012 76012 22024
rect 53156 21984 55904 22012
rect 55968 21984 76012 22012
rect 53156 21972 53162 21984
rect 55968 21944 55996 21984
rect 76006 21972 76012 21984
rect 76064 21972 76070 22024
rect 84749 22015 84807 22021
rect 84749 21981 84761 22015
rect 84795 22012 84807 22015
rect 85132 22012 85160 22052
rect 85393 22049 85405 22052
rect 85439 22049 85451 22083
rect 85393 22043 85451 22049
rect 85482 22040 85488 22092
rect 85540 22080 85546 22092
rect 85761 22083 85819 22089
rect 85761 22080 85773 22083
rect 85540 22052 85773 22080
rect 85540 22040 85546 22052
rect 85761 22049 85773 22052
rect 85807 22049 85819 22083
rect 85761 22043 85819 22049
rect 85298 22012 85304 22024
rect 84795 21984 85160 22012
rect 85259 21984 85304 22012
rect 84795 21981 84807 21984
rect 84749 21975 84807 21981
rect 85298 21972 85304 21984
rect 85356 21972 85362 22024
rect 85669 22015 85727 22021
rect 85669 21981 85681 22015
rect 85715 21981 85727 22015
rect 85669 21975 85727 21981
rect 43487 21916 55996 21944
rect 43487 21913 43499 21916
rect 43441 21907 43499 21913
rect 56134 21904 56140 21956
rect 56192 21944 56198 21956
rect 56192 21916 58848 21944
rect 56192 21904 56198 21916
rect 46290 21876 46296 21888
rect 41616 21848 46296 21876
rect 46290 21836 46296 21848
rect 46348 21836 46354 21888
rect 51718 21836 51724 21888
rect 51776 21876 51782 21888
rect 53098 21876 53104 21888
rect 51776 21848 53104 21876
rect 51776 21836 51782 21848
rect 53098 21836 53104 21848
rect 53156 21836 53162 21888
rect 53190 21836 53196 21888
rect 53248 21876 53254 21888
rect 56962 21876 56968 21888
rect 53248 21848 56968 21876
rect 53248 21836 53254 21848
rect 56962 21836 56968 21848
rect 57020 21836 57026 21888
rect 58618 21876 58624 21888
rect 58579 21848 58624 21876
rect 58618 21836 58624 21848
rect 58676 21836 58682 21888
rect 58820 21876 58848 21916
rect 58894 21904 58900 21956
rect 58952 21944 58958 21956
rect 60826 21944 60832 21956
rect 58952 21916 60832 21944
rect 58952 21904 58958 21916
rect 60826 21904 60832 21916
rect 60884 21904 60890 21956
rect 60936 21916 61424 21944
rect 60936 21876 60964 21916
rect 58820 21848 60964 21876
rect 61396 21876 61424 21916
rect 62666 21904 62672 21956
rect 62724 21944 62730 21956
rect 85684 21944 85712 21975
rect 62724 21916 85712 21944
rect 62724 21904 62730 21916
rect 88242 21904 88248 21956
rect 88300 21944 88306 21956
rect 92842 21944 92848 21956
rect 88300 21916 92848 21944
rect 88300 21904 88306 21916
rect 92842 21904 92848 21916
rect 92900 21904 92906 21956
rect 84749 21879 84807 21885
rect 84749 21876 84761 21879
rect 61396 21848 84761 21876
rect 84749 21845 84761 21848
rect 84795 21876 84807 21879
rect 84841 21879 84899 21885
rect 84841 21876 84853 21879
rect 84795 21848 84853 21876
rect 84795 21845 84807 21848
rect 84749 21839 84807 21845
rect 84841 21845 84853 21848
rect 84887 21845 84899 21879
rect 84841 21839 84899 21845
rect 85114 21836 85120 21888
rect 85172 21876 85178 21888
rect 86221 21879 86279 21885
rect 86221 21876 86233 21879
rect 85172 21848 86233 21876
rect 85172 21836 85178 21848
rect 86221 21845 86233 21848
rect 86267 21845 86279 21879
rect 86221 21839 86279 21845
rect 1104 21786 98808 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 65686 21786
rect 65738 21734 65750 21786
rect 65802 21734 65814 21786
rect 65866 21734 65878 21786
rect 65930 21734 96406 21786
rect 96458 21734 96470 21786
rect 96522 21734 96534 21786
rect 96586 21734 96598 21786
rect 96650 21734 98808 21786
rect 1104 21712 98808 21734
rect 17402 21632 17408 21684
rect 17460 21672 17466 21684
rect 17770 21672 17776 21684
rect 17460 21644 17776 21672
rect 17460 21632 17466 21644
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 43717 21675 43775 21681
rect 43717 21672 43729 21675
rect 22066 21644 43729 21672
rect 5442 21564 5448 21616
rect 5500 21604 5506 21616
rect 17310 21604 17316 21616
rect 5500 21576 17316 21604
rect 5500 21564 5506 21576
rect 17310 21564 17316 21576
rect 17368 21564 17374 21616
rect 2406 21496 2412 21548
rect 2464 21536 2470 21548
rect 12437 21539 12495 21545
rect 2464 21508 2774 21536
rect 2464 21496 2470 21508
rect 2746 21332 2774 21508
rect 12437 21505 12449 21539
rect 12483 21536 12495 21539
rect 22066 21536 22094 21644
rect 43717 21641 43729 21644
rect 43763 21641 43775 21675
rect 50890 21672 50896 21684
rect 43717 21635 43775 21641
rect 43824 21644 50896 21672
rect 25866 21564 25872 21616
rect 25924 21604 25930 21616
rect 28902 21604 28908 21616
rect 25924 21576 28908 21604
rect 25924 21564 25930 21576
rect 28902 21564 28908 21576
rect 28960 21564 28966 21616
rect 32858 21604 32864 21616
rect 32819 21576 32864 21604
rect 32858 21564 32864 21576
rect 32916 21604 32922 21616
rect 33229 21607 33287 21613
rect 33229 21604 33241 21607
rect 32916 21576 33241 21604
rect 32916 21564 32922 21576
rect 33229 21573 33241 21576
rect 33275 21573 33287 21607
rect 33229 21567 33287 21573
rect 34054 21564 34060 21616
rect 34112 21604 34118 21616
rect 37090 21604 37096 21616
rect 34112 21576 37096 21604
rect 34112 21564 34118 21576
rect 37090 21564 37096 21576
rect 37148 21564 37154 21616
rect 37366 21564 37372 21616
rect 37424 21604 37430 21616
rect 40034 21604 40040 21616
rect 37424 21576 40040 21604
rect 37424 21564 37430 21576
rect 40034 21564 40040 21576
rect 40092 21564 40098 21616
rect 42242 21564 42248 21616
rect 42300 21604 42306 21616
rect 43824 21604 43852 21644
rect 50890 21632 50896 21644
rect 50948 21632 50954 21684
rect 51350 21672 51356 21684
rect 51046 21644 51356 21672
rect 43990 21604 43996 21616
rect 42300 21576 43852 21604
rect 43951 21576 43996 21604
rect 42300 21564 42306 21576
rect 43990 21564 43996 21576
rect 44048 21564 44054 21616
rect 44542 21564 44548 21616
rect 44600 21604 44606 21616
rect 51046 21604 51074 21644
rect 51350 21632 51356 21644
rect 51408 21632 51414 21684
rect 51460 21644 54984 21672
rect 44600 21576 51074 21604
rect 44600 21564 44606 21576
rect 12483 21508 22094 21536
rect 12483 21505 12495 21508
rect 12437 21499 12495 21505
rect 25406 21496 25412 21548
rect 25464 21536 25470 21548
rect 25464 21508 26060 21536
rect 25464 21496 25470 21508
rect 12066 21468 12072 21480
rect 12027 21440 12072 21468
rect 12066 21428 12072 21440
rect 12124 21428 12130 21480
rect 12158 21428 12164 21480
rect 12216 21468 12222 21480
rect 12253 21471 12311 21477
rect 12253 21468 12265 21471
rect 12216 21440 12265 21468
rect 12216 21428 12222 21440
rect 12253 21437 12265 21440
rect 12299 21437 12311 21471
rect 12253 21431 12311 21437
rect 12345 21471 12403 21477
rect 12345 21437 12357 21471
rect 12391 21437 12403 21471
rect 12618 21468 12624 21480
rect 12579 21440 12624 21468
rect 12345 21431 12403 21437
rect 12360 21400 12388 21431
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 12802 21468 12808 21480
rect 12763 21440 12808 21468
rect 12802 21428 12808 21440
rect 12860 21428 12866 21480
rect 17126 21428 17132 21480
rect 17184 21468 17190 21480
rect 25866 21468 25872 21480
rect 17184 21440 25872 21468
rect 17184 21428 17190 21440
rect 25866 21428 25872 21440
rect 25924 21428 25930 21480
rect 26032 21477 26060 21508
rect 32214 21496 32220 21548
rect 32272 21536 32278 21548
rect 34790 21536 34796 21548
rect 32272 21508 34796 21536
rect 32272 21496 32278 21508
rect 34790 21496 34796 21508
rect 34848 21496 34854 21548
rect 35342 21496 35348 21548
rect 35400 21536 35406 21548
rect 51460 21536 51488 21644
rect 54956 21604 54984 21644
rect 55030 21632 55036 21684
rect 55088 21672 55094 21684
rect 58713 21675 58771 21681
rect 58713 21672 58725 21675
rect 55088 21644 58725 21672
rect 55088 21632 55094 21644
rect 58713 21641 58725 21644
rect 58759 21641 58771 21675
rect 58713 21635 58771 21641
rect 60553 21675 60611 21681
rect 60553 21641 60565 21675
rect 60599 21672 60611 21675
rect 62666 21672 62672 21684
rect 60599 21644 62672 21672
rect 60599 21641 60611 21644
rect 60553 21635 60611 21641
rect 62666 21632 62672 21644
rect 62724 21632 62730 21684
rect 66254 21632 66260 21684
rect 66312 21672 66318 21684
rect 85482 21672 85488 21684
rect 66312 21644 85488 21672
rect 66312 21632 66318 21644
rect 85482 21632 85488 21644
rect 85540 21632 85546 21684
rect 60826 21604 60832 21616
rect 54956 21576 60832 21604
rect 60826 21564 60832 21576
rect 60884 21564 60890 21616
rect 61010 21604 61016 21616
rect 60936 21576 61016 21604
rect 52270 21536 52276 21548
rect 35400 21508 43484 21536
rect 35400 21496 35406 21508
rect 26017 21471 26075 21477
rect 26017 21437 26029 21471
rect 26063 21437 26075 21471
rect 26142 21468 26148 21480
rect 26103 21440 26148 21468
rect 26017 21431 26075 21437
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 26237 21471 26295 21477
rect 26237 21437 26249 21471
rect 26283 21437 26295 21471
rect 26237 21431 26295 21437
rect 17218 21400 17224 21412
rect 12360 21372 17224 21400
rect 17218 21360 17224 21372
rect 17276 21360 17282 21412
rect 17494 21360 17500 21412
rect 17552 21400 17558 21412
rect 25590 21400 25596 21412
rect 17552 21372 25596 21400
rect 17552 21360 17558 21372
rect 25590 21360 25596 21372
rect 25648 21360 25654 21412
rect 26252 21400 26280 21431
rect 26326 21428 26332 21480
rect 26384 21468 26390 21480
rect 26421 21471 26479 21477
rect 26421 21468 26433 21471
rect 26384 21440 26433 21468
rect 26384 21428 26390 21440
rect 26421 21437 26433 21440
rect 26467 21437 26479 21471
rect 26421 21431 26479 21437
rect 38562 21428 38568 21480
rect 38620 21468 38626 21480
rect 38620 21440 38700 21468
rect 38620 21428 38626 21440
rect 26878 21400 26884 21412
rect 26252 21372 26884 21400
rect 26878 21360 26884 21372
rect 26936 21400 26942 21412
rect 27798 21400 27804 21412
rect 26936 21372 27804 21400
rect 26936 21360 26942 21372
rect 27798 21360 27804 21372
rect 27856 21360 27862 21412
rect 33778 21360 33784 21412
rect 33836 21400 33842 21412
rect 38672 21400 38700 21440
rect 38746 21428 38752 21480
rect 38804 21468 38810 21480
rect 39390 21468 39396 21480
rect 38804 21440 39396 21468
rect 38804 21428 38810 21440
rect 39390 21428 39396 21440
rect 39448 21428 39454 21480
rect 39669 21471 39727 21477
rect 39669 21437 39681 21471
rect 39715 21468 39727 21471
rect 41141 21471 41199 21477
rect 41141 21468 41153 21471
rect 39715 21440 41153 21468
rect 39715 21437 39727 21440
rect 39669 21431 39727 21437
rect 41141 21437 41153 21440
rect 41187 21468 41199 21471
rect 41187 21440 41368 21468
rect 41187 21437 41199 21440
rect 41141 21431 41199 21437
rect 39761 21403 39819 21409
rect 39761 21400 39773 21403
rect 33836 21372 38608 21400
rect 38672 21372 39773 21400
rect 33836 21360 33842 21372
rect 16298 21332 16304 21344
rect 2746 21304 16304 21332
rect 16298 21292 16304 21304
rect 16356 21292 16362 21344
rect 26234 21292 26240 21344
rect 26292 21332 26298 21344
rect 26513 21335 26571 21341
rect 26513 21332 26525 21335
rect 26292 21304 26525 21332
rect 26292 21292 26298 21304
rect 26513 21301 26525 21304
rect 26559 21301 26571 21335
rect 26513 21295 26571 21301
rect 35250 21292 35256 21344
rect 35308 21332 35314 21344
rect 35710 21332 35716 21344
rect 35308 21304 35716 21332
rect 35308 21292 35314 21304
rect 35710 21292 35716 21304
rect 35768 21292 35774 21344
rect 37918 21292 37924 21344
rect 37976 21332 37982 21344
rect 38470 21332 38476 21344
rect 37976 21304 38476 21332
rect 37976 21292 37982 21304
rect 38470 21292 38476 21304
rect 38528 21292 38534 21344
rect 38580 21332 38608 21372
rect 39761 21369 39773 21372
rect 39807 21369 39819 21403
rect 41340 21400 41368 21440
rect 41414 21428 41420 21480
rect 41472 21468 41478 21480
rect 43456 21468 43484 21508
rect 44192 21508 51488 21536
rect 51552 21508 52132 21536
rect 52231 21508 52276 21536
rect 44192 21468 44220 21508
rect 41472 21440 41517 21468
rect 43456 21440 44220 21468
rect 41472 21428 41478 21440
rect 46198 21428 46204 21480
rect 46256 21468 46262 21480
rect 51552 21468 51580 21508
rect 52104 21477 52132 21508
rect 52270 21496 52276 21508
rect 52328 21496 52334 21548
rect 52546 21536 52552 21548
rect 52472 21508 52552 21536
rect 46256 21440 51580 21468
rect 51905 21471 51963 21477
rect 46256 21428 46262 21440
rect 51905 21437 51917 21471
rect 51951 21437 51963 21471
rect 51905 21431 51963 21437
rect 52089 21471 52147 21477
rect 52089 21437 52101 21471
rect 52135 21437 52147 21471
rect 52089 21431 52147 21437
rect 41506 21400 41512 21412
rect 41340 21372 41512 21400
rect 39761 21363 39819 21369
rect 41506 21360 41512 21372
rect 41564 21360 41570 21412
rect 44082 21360 44088 21412
rect 44140 21400 44146 21412
rect 49234 21400 49240 21412
rect 44140 21372 49240 21400
rect 44140 21360 44146 21372
rect 49234 21360 49240 21372
rect 49292 21360 49298 21412
rect 50154 21360 50160 21412
rect 50212 21400 50218 21412
rect 51920 21400 51948 21431
rect 52178 21428 52184 21480
rect 52236 21468 52242 21480
rect 52472 21477 52500 21508
rect 52546 21496 52552 21508
rect 52604 21496 52610 21548
rect 54018 21536 54024 21548
rect 53979 21508 54024 21536
rect 54018 21496 54024 21508
rect 54076 21496 54082 21548
rect 54386 21496 54392 21548
rect 54444 21536 54450 21548
rect 58618 21536 58624 21548
rect 54444 21508 58624 21536
rect 54444 21496 54450 21508
rect 58618 21496 58624 21508
rect 58676 21496 58682 21548
rect 58713 21539 58771 21545
rect 58713 21505 58725 21539
rect 58759 21536 58771 21539
rect 58986 21536 58992 21548
rect 58759 21508 58992 21536
rect 58759 21505 58771 21508
rect 58713 21499 58771 21505
rect 58986 21496 58992 21508
rect 59044 21496 59050 21548
rect 52457 21471 52515 21477
rect 52236 21440 52281 21468
rect 52236 21428 52242 21440
rect 52457 21437 52469 21471
rect 52503 21437 52515 21471
rect 52457 21431 52515 21437
rect 53742 21428 53748 21480
rect 53800 21468 53806 21480
rect 54297 21471 54355 21477
rect 54297 21468 54309 21471
rect 53800 21440 54309 21468
rect 53800 21428 53806 21440
rect 54297 21437 54309 21440
rect 54343 21437 54355 21471
rect 55674 21468 55680 21480
rect 55587 21440 55680 21468
rect 54297 21431 54355 21437
rect 55674 21428 55680 21440
rect 55732 21468 55738 21480
rect 59354 21468 59360 21480
rect 55732 21440 59360 21468
rect 55732 21428 55738 21440
rect 59354 21428 59360 21440
rect 59412 21428 59418 21480
rect 60458 21428 60464 21480
rect 60516 21468 60522 21480
rect 60645 21471 60703 21477
rect 60645 21468 60657 21471
rect 60516 21440 60657 21468
rect 60516 21428 60522 21440
rect 60645 21437 60657 21440
rect 60691 21437 60703 21471
rect 60826 21468 60832 21480
rect 60787 21440 60832 21468
rect 60645 21431 60703 21437
rect 60826 21428 60832 21440
rect 60884 21428 60890 21480
rect 60936 21477 60964 21576
rect 61010 21564 61016 21576
rect 61068 21564 61074 21616
rect 61102 21564 61108 21616
rect 61160 21604 61166 21616
rect 77938 21604 77944 21616
rect 61160 21576 77944 21604
rect 61160 21564 61166 21576
rect 77938 21564 77944 21576
rect 77996 21564 78002 21616
rect 80698 21564 80704 21616
rect 80756 21604 80762 21616
rect 86310 21604 86316 21616
rect 80756 21576 86316 21604
rect 80756 21564 80762 21576
rect 86310 21564 86316 21576
rect 86368 21564 86374 21616
rect 61838 21536 61844 21548
rect 61212 21508 61844 21536
rect 61212 21477 61240 21508
rect 61838 21496 61844 21508
rect 61896 21536 61902 21548
rect 64414 21536 64420 21548
rect 61896 21508 64420 21536
rect 61896 21496 61902 21508
rect 64414 21496 64420 21508
rect 64472 21496 64478 21548
rect 65150 21536 65156 21548
rect 65111 21508 65156 21536
rect 65150 21496 65156 21508
rect 65208 21496 65214 21548
rect 65242 21496 65248 21548
rect 65300 21536 65306 21548
rect 78030 21536 78036 21548
rect 65300 21508 78036 21536
rect 65300 21496 65306 21508
rect 78030 21496 78036 21508
rect 78088 21496 78094 21548
rect 78122 21496 78128 21548
rect 78180 21536 78186 21548
rect 93854 21536 93860 21548
rect 78180 21508 93860 21536
rect 78180 21496 78186 21508
rect 93854 21496 93860 21508
rect 93912 21496 93918 21548
rect 60924 21471 60982 21477
rect 60924 21437 60936 21471
rect 60970 21437 60982 21471
rect 60924 21431 60982 21437
rect 61013 21471 61071 21477
rect 61013 21437 61025 21471
rect 61059 21437 61071 21471
rect 61013 21431 61071 21437
rect 61180 21471 61240 21477
rect 61180 21437 61192 21471
rect 61226 21440 61240 21471
rect 61226 21437 61238 21440
rect 61180 21431 61238 21437
rect 53190 21400 53196 21412
rect 50212 21372 53196 21400
rect 50212 21360 50218 21372
rect 53190 21360 53196 21372
rect 53248 21360 53254 21412
rect 55030 21360 55036 21412
rect 55088 21400 55094 21412
rect 60553 21403 60611 21409
rect 60553 21400 60565 21403
rect 55088 21372 60565 21400
rect 55088 21360 55094 21372
rect 60553 21369 60565 21372
rect 60599 21369 60611 21403
rect 61028 21400 61056 21431
rect 61562 21428 61568 21480
rect 61620 21468 61626 21480
rect 80698 21468 80704 21480
rect 61620 21440 80704 21468
rect 61620 21428 61626 21440
rect 80698 21428 80704 21440
rect 80756 21428 80762 21480
rect 82446 21428 82452 21480
rect 82504 21468 82510 21480
rect 82541 21471 82599 21477
rect 82541 21468 82553 21471
rect 82504 21440 82553 21468
rect 82504 21428 82510 21440
rect 82541 21437 82553 21440
rect 82587 21437 82599 21471
rect 82541 21431 82599 21437
rect 62574 21400 62580 21412
rect 61028 21372 62580 21400
rect 60553 21363 60611 21369
rect 62574 21360 62580 21372
rect 62632 21360 62638 21412
rect 62666 21360 62672 21412
rect 62724 21400 62730 21412
rect 90634 21400 90640 21412
rect 62724 21372 90640 21400
rect 62724 21360 62730 21372
rect 90634 21360 90640 21372
rect 90692 21360 90698 21412
rect 38746 21332 38752 21344
rect 38580 21304 38752 21332
rect 38746 21292 38752 21304
rect 38804 21292 38810 21344
rect 40402 21292 40408 21344
rect 40460 21332 40466 21344
rect 42886 21332 42892 21344
rect 40460 21304 42892 21332
rect 40460 21292 40466 21304
rect 42886 21292 42892 21304
rect 42944 21292 42950 21344
rect 43717 21335 43775 21341
rect 43717 21301 43729 21335
rect 43763 21332 43775 21335
rect 48682 21332 48688 21344
rect 43763 21304 48688 21332
rect 43763 21301 43775 21304
rect 43717 21295 43775 21301
rect 48682 21292 48688 21304
rect 48740 21292 48746 21344
rect 50614 21292 50620 21344
rect 50672 21332 50678 21344
rect 52270 21332 52276 21344
rect 50672 21304 52276 21332
rect 50672 21292 50678 21304
rect 52270 21292 52276 21304
rect 52328 21292 52334 21344
rect 52641 21335 52699 21341
rect 52641 21301 52653 21335
rect 52687 21332 52699 21335
rect 52730 21332 52736 21344
rect 52687 21304 52736 21332
rect 52687 21301 52699 21304
rect 52641 21295 52699 21301
rect 52730 21292 52736 21304
rect 52788 21292 52794 21344
rect 55858 21292 55864 21344
rect 55916 21332 55922 21344
rect 61286 21332 61292 21344
rect 55916 21304 61292 21332
rect 55916 21292 55922 21304
rect 61286 21292 61292 21304
rect 61344 21292 61350 21344
rect 61381 21335 61439 21341
rect 61381 21301 61393 21335
rect 61427 21332 61439 21335
rect 62942 21332 62948 21344
rect 61427 21304 62948 21332
rect 61427 21301 61439 21304
rect 61381 21295 61439 21301
rect 62942 21292 62948 21304
rect 63000 21292 63006 21344
rect 63586 21292 63592 21344
rect 63644 21332 63650 21344
rect 66254 21332 66260 21344
rect 63644 21304 66260 21332
rect 63644 21292 63650 21304
rect 66254 21292 66260 21304
rect 66312 21292 66318 21344
rect 1104 21242 98808 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 50326 21242
rect 50378 21190 50390 21242
rect 50442 21190 50454 21242
rect 50506 21190 50518 21242
rect 50570 21190 81046 21242
rect 81098 21190 81110 21242
rect 81162 21190 81174 21242
rect 81226 21190 81238 21242
rect 81290 21190 98808 21242
rect 1104 21168 98808 21190
rect 1854 21128 1860 21140
rect 1815 21100 1860 21128
rect 1854 21088 1860 21100
rect 1912 21088 1918 21140
rect 2685 21131 2743 21137
rect 2685 21097 2697 21131
rect 2731 21128 2743 21131
rect 17494 21128 17500 21140
rect 2731 21100 17356 21128
rect 17455 21100 17500 21128
rect 2731 21097 2743 21100
rect 2685 21091 2743 21097
rect 1673 21063 1731 21069
rect 1673 21029 1685 21063
rect 1719 21060 1731 21063
rect 2700 21060 2728 21091
rect 1719 21032 2176 21060
rect 1719 21029 1731 21032
rect 1673 21023 1731 21029
rect 1489 20995 1547 21001
rect 1489 20961 1501 20995
rect 1535 20992 1547 20995
rect 1949 20995 2007 21001
rect 1949 20992 1961 20995
rect 1535 20964 1961 20992
rect 1535 20961 1547 20964
rect 1489 20955 1547 20961
rect 1949 20961 1961 20964
rect 1995 20992 2007 20995
rect 1995 20964 2084 20992
rect 1995 20961 2007 20964
rect 1949 20955 2007 20961
rect 2056 20856 2084 20964
rect 2148 20933 2176 21032
rect 2240 21032 2728 21060
rect 4985 21063 5043 21069
rect 2240 21001 2268 21032
rect 4985 21029 4997 21063
rect 5031 21060 5043 21063
rect 6178 21060 6184 21072
rect 5031 21032 6040 21060
rect 6139 21032 6184 21060
rect 5031 21029 5043 21032
rect 4985 21023 5043 21029
rect 2406 21001 2412 21004
rect 2225 20995 2283 21001
rect 2225 20961 2237 20995
rect 2271 20961 2283 20995
rect 2225 20955 2283 20961
rect 2353 20995 2412 21001
rect 2353 20961 2365 20995
rect 2399 20961 2412 20995
rect 2353 20955 2412 20961
rect 2406 20952 2412 20955
rect 2464 20952 2470 21004
rect 2501 20995 2559 21001
rect 2501 20961 2513 20995
rect 2547 20992 2559 20995
rect 4890 20992 4896 21004
rect 2547 20964 4896 20992
rect 2547 20961 2559 20964
rect 2501 20955 2559 20961
rect 4890 20952 4896 20964
rect 4948 20952 4954 21004
rect 5442 20992 5448 21004
rect 5403 20964 5448 20992
rect 5442 20952 5448 20964
rect 5500 20952 5506 21004
rect 5902 21001 5908 21004
rect 5849 20995 5908 21001
rect 5849 20961 5861 20995
rect 5895 20961 5908 20995
rect 5849 20955 5908 20961
rect 5902 20952 5908 20955
rect 5960 20952 5966 21004
rect 6012 21001 6040 21032
rect 6178 21020 6184 21032
rect 6236 21020 6242 21072
rect 17328 21060 17356 21100
rect 17494 21088 17500 21100
rect 17552 21088 17558 21140
rect 26142 21088 26148 21140
rect 26200 21128 26206 21140
rect 42794 21128 42800 21140
rect 26200 21100 42800 21128
rect 26200 21088 26206 21100
rect 42794 21088 42800 21100
rect 42852 21088 42858 21140
rect 42886 21088 42892 21140
rect 42944 21128 42950 21140
rect 47670 21128 47676 21140
rect 42944 21100 47676 21128
rect 42944 21088 42950 21100
rect 47670 21088 47676 21100
rect 47728 21088 47734 21140
rect 51350 21088 51356 21140
rect 51408 21128 51414 21140
rect 55858 21128 55864 21140
rect 51408 21100 55864 21128
rect 51408 21088 51414 21100
rect 55858 21088 55864 21100
rect 55916 21088 55922 21140
rect 58894 21128 58900 21140
rect 55968 21100 58900 21128
rect 18782 21060 18788 21072
rect 17328 21032 18788 21060
rect 18782 21020 18788 21032
rect 18840 21060 18846 21072
rect 55968 21060 55996 21100
rect 58894 21088 58900 21100
rect 58952 21088 58958 21140
rect 58986 21088 58992 21140
rect 59044 21128 59050 21140
rect 81526 21128 81532 21140
rect 59044 21100 81532 21128
rect 59044 21088 59050 21100
rect 81526 21088 81532 21100
rect 81584 21088 81590 21140
rect 84194 21128 84200 21140
rect 81636 21100 84200 21128
rect 18840 21032 55996 21060
rect 18840 21020 18846 21032
rect 57422 21020 57428 21072
rect 57480 21060 57486 21072
rect 61838 21060 61844 21072
rect 57480 21032 61844 21060
rect 57480 21020 57486 21032
rect 61838 21020 61844 21032
rect 61896 21020 61902 21072
rect 63405 21063 63463 21069
rect 63405 21060 63417 21063
rect 62960 21032 63417 21060
rect 5997 20995 6055 21001
rect 5997 20961 6009 20995
rect 6043 20992 6055 20995
rect 14550 20992 14556 21004
rect 6043 20964 14556 20992
rect 6043 20961 6055 20964
rect 5997 20955 6055 20961
rect 14550 20952 14556 20964
rect 14608 20952 14614 21004
rect 15930 20992 15936 21004
rect 15891 20964 15936 20992
rect 15930 20952 15936 20964
rect 15988 20952 15994 21004
rect 17954 20952 17960 21004
rect 18012 20992 18018 21004
rect 18601 20995 18659 21001
rect 18601 20992 18613 20995
rect 18012 20964 18613 20992
rect 18012 20952 18018 20964
rect 18601 20961 18613 20964
rect 18647 20961 18659 20995
rect 18601 20955 18659 20961
rect 26050 20952 26056 21004
rect 26108 20992 26114 21004
rect 44269 20995 44327 21001
rect 44269 20992 44281 20995
rect 26108 20964 44281 20992
rect 26108 20952 26114 20964
rect 44269 20961 44281 20964
rect 44315 20992 44327 20995
rect 45922 20992 45928 21004
rect 44315 20964 45928 20992
rect 44315 20961 44327 20964
rect 44269 20955 44327 20961
rect 45922 20952 45928 20964
rect 45980 20952 45986 21004
rect 46106 20952 46112 21004
rect 46164 20992 46170 21004
rect 51074 20992 51080 21004
rect 46164 20964 51080 20992
rect 46164 20952 46170 20964
rect 51074 20952 51080 20964
rect 51132 20952 51138 21004
rect 51166 20952 51172 21004
rect 51224 20992 51230 21004
rect 62960 20992 62988 21032
rect 63405 21029 63417 21032
rect 63451 21060 63463 21063
rect 63451 21032 70394 21060
rect 63451 21029 63463 21032
rect 63405 21023 63463 21029
rect 63218 20992 63224 21004
rect 51224 20964 62988 20992
rect 63179 20964 63224 20992
rect 51224 20952 51230 20964
rect 63218 20952 63224 20964
rect 63276 20952 63282 21004
rect 63497 20995 63555 21001
rect 63497 20961 63509 20995
rect 63543 20992 63555 20995
rect 63678 20992 63684 21004
rect 63543 20964 63684 20992
rect 63543 20961 63555 20964
rect 63497 20955 63555 20961
rect 63678 20952 63684 20964
rect 63736 20952 63742 21004
rect 67358 20992 67364 21004
rect 67319 20964 67364 20992
rect 67358 20952 67364 20964
rect 67416 20952 67422 21004
rect 70366 20992 70394 21032
rect 72142 21020 72148 21072
rect 72200 21060 72206 21072
rect 73706 21060 73712 21072
rect 72200 21032 73712 21060
rect 72200 21020 72206 21032
rect 73706 21020 73712 21032
rect 73764 21020 73770 21072
rect 75638 20992 75644 21004
rect 70366 20964 75644 20992
rect 75638 20952 75644 20964
rect 75696 20952 75702 21004
rect 80333 20995 80391 21001
rect 80333 20961 80345 20995
rect 80379 20992 80391 20995
rect 81636 20992 81664 21100
rect 84194 21088 84200 21100
rect 84252 21088 84258 21140
rect 81713 21063 81771 21069
rect 81713 21029 81725 21063
rect 81759 21060 81771 21063
rect 85574 21060 85580 21072
rect 81759 21032 85580 21060
rect 81759 21029 81771 21032
rect 81713 21023 81771 21029
rect 80379 20964 81664 20992
rect 80379 20961 80391 20964
rect 80333 20955 80391 20961
rect 2133 20927 2191 20933
rect 2133 20893 2145 20927
rect 2179 20924 2191 20927
rect 5169 20927 5227 20933
rect 2179 20896 5120 20924
rect 2179 20893 2191 20896
rect 2133 20887 2191 20893
rect 3418 20856 3424 20868
rect 2056 20828 3424 20856
rect 3418 20816 3424 20828
rect 3476 20816 3482 20868
rect 5092 20856 5120 20896
rect 5169 20893 5181 20927
rect 5215 20924 5227 20927
rect 5626 20924 5632 20936
rect 5215 20896 5632 20924
rect 5215 20893 5227 20896
rect 5169 20887 5227 20893
rect 5626 20884 5632 20896
rect 5684 20884 5690 20936
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20924 5779 20927
rect 6178 20924 6184 20936
rect 5767 20896 6184 20924
rect 5767 20893 5779 20896
rect 5721 20887 5779 20893
rect 6178 20884 6184 20896
rect 6236 20884 6242 20936
rect 15746 20884 15752 20936
rect 15804 20924 15810 20936
rect 16209 20927 16267 20933
rect 16209 20924 16221 20927
rect 15804 20896 16221 20924
rect 15804 20884 15810 20896
rect 16209 20893 16221 20896
rect 16255 20893 16267 20927
rect 18785 20927 18843 20933
rect 18785 20924 18797 20927
rect 16209 20887 16267 20893
rect 17052 20896 18797 20924
rect 5534 20856 5540 20868
rect 5092 20828 5540 20856
rect 5534 20816 5540 20828
rect 5592 20816 5598 20868
rect 5902 20816 5908 20868
rect 5960 20856 5966 20868
rect 8110 20856 8116 20868
rect 5960 20828 8116 20856
rect 5960 20816 5966 20828
rect 8110 20816 8116 20828
rect 8168 20816 8174 20868
rect 5353 20791 5411 20797
rect 5353 20757 5365 20791
rect 5399 20788 5411 20791
rect 6638 20788 6644 20800
rect 5399 20760 6644 20788
rect 5399 20757 5411 20760
rect 5353 20751 5411 20757
rect 6638 20748 6644 20760
rect 6696 20748 6702 20800
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 12158 20788 12164 20800
rect 11112 20760 12164 20788
rect 11112 20748 11118 20760
rect 12158 20748 12164 20760
rect 12216 20748 12222 20800
rect 14734 20748 14740 20800
rect 14792 20788 14798 20800
rect 17052 20788 17080 20896
rect 18785 20893 18797 20896
rect 18831 20924 18843 20927
rect 26786 20924 26792 20936
rect 18831 20896 26792 20924
rect 18831 20893 18843 20896
rect 18785 20887 18843 20893
rect 26786 20884 26792 20896
rect 26844 20884 26850 20936
rect 28994 20884 29000 20936
rect 29052 20924 29058 20936
rect 30098 20924 30104 20936
rect 29052 20896 30104 20924
rect 29052 20884 29058 20896
rect 30098 20884 30104 20896
rect 30156 20884 30162 20936
rect 35250 20884 35256 20936
rect 35308 20924 35314 20936
rect 35308 20896 38516 20924
rect 35308 20884 35314 20896
rect 17126 20816 17132 20868
rect 17184 20856 17190 20868
rect 17494 20856 17500 20868
rect 17184 20828 17500 20856
rect 17184 20816 17190 20828
rect 17494 20816 17500 20828
rect 17552 20816 17558 20868
rect 21726 20816 21732 20868
rect 21784 20856 21790 20868
rect 38378 20856 38384 20868
rect 21784 20828 38384 20856
rect 21784 20816 21790 20828
rect 38378 20816 38384 20828
rect 38436 20816 38442 20868
rect 38488 20856 38516 20896
rect 42794 20884 42800 20936
rect 42852 20924 42858 20936
rect 44082 20924 44088 20936
rect 42852 20896 44088 20924
rect 42852 20884 42858 20896
rect 44082 20884 44088 20896
rect 44140 20884 44146 20936
rect 44542 20924 44548 20936
rect 44503 20896 44548 20924
rect 44542 20884 44548 20896
rect 44600 20884 44606 20936
rect 78030 20924 78036 20936
rect 45572 20896 78036 20924
rect 45572 20856 45600 20896
rect 78030 20884 78036 20896
rect 78088 20884 78094 20936
rect 80054 20884 80060 20936
rect 80112 20924 80118 20936
rect 80112 20896 80157 20924
rect 80112 20884 80118 20896
rect 38488 20828 45600 20856
rect 45922 20816 45928 20868
rect 45980 20856 45986 20868
rect 46934 20856 46940 20868
rect 45980 20828 46940 20856
rect 45980 20816 45986 20828
rect 46934 20816 46940 20828
rect 46992 20816 46998 20868
rect 47946 20816 47952 20868
rect 48004 20856 48010 20868
rect 50890 20856 50896 20868
rect 48004 20828 50896 20856
rect 48004 20816 48010 20828
rect 50890 20816 50896 20828
rect 50948 20816 50954 20868
rect 51074 20816 51080 20868
rect 51132 20856 51138 20868
rect 55674 20856 55680 20868
rect 51132 20828 55680 20856
rect 51132 20816 51138 20828
rect 55674 20816 55680 20828
rect 55732 20816 55738 20868
rect 55858 20816 55864 20868
rect 55916 20856 55922 20868
rect 60550 20856 60556 20868
rect 55916 20828 60556 20856
rect 55916 20816 55922 20828
rect 60550 20816 60556 20828
rect 60608 20816 60614 20868
rect 60706 20828 70394 20856
rect 14792 20760 17080 20788
rect 14792 20748 14798 20760
rect 17218 20748 17224 20800
rect 17276 20788 17282 20800
rect 29086 20788 29092 20800
rect 17276 20760 29092 20788
rect 17276 20748 17282 20760
rect 29086 20748 29092 20760
rect 29144 20748 29150 20800
rect 35894 20748 35900 20800
rect 35952 20788 35958 20800
rect 36998 20788 37004 20800
rect 35952 20760 37004 20788
rect 35952 20748 35958 20760
rect 36998 20748 37004 20760
rect 37056 20748 37062 20800
rect 37918 20748 37924 20800
rect 37976 20788 37982 20800
rect 38286 20788 38292 20800
rect 37976 20760 38292 20788
rect 37976 20748 37982 20760
rect 38286 20748 38292 20760
rect 38344 20748 38350 20800
rect 38746 20748 38752 20800
rect 38804 20788 38810 20800
rect 60706 20788 60734 20828
rect 38804 20760 60734 20788
rect 38804 20748 38810 20760
rect 62850 20748 62856 20800
rect 62908 20788 62914 20800
rect 63037 20791 63095 20797
rect 63037 20788 63049 20791
rect 62908 20760 63049 20788
rect 62908 20748 62914 20760
rect 63037 20757 63049 20760
rect 63083 20757 63095 20791
rect 64138 20788 64144 20800
rect 64099 20760 64144 20788
rect 63037 20751 63095 20757
rect 64138 20748 64144 20760
rect 64196 20748 64202 20800
rect 64414 20748 64420 20800
rect 64472 20788 64478 20800
rect 65058 20788 65064 20800
rect 64472 20760 65064 20788
rect 64472 20748 64478 20760
rect 65058 20748 65064 20760
rect 65116 20748 65122 20800
rect 65150 20748 65156 20800
rect 65208 20788 65214 20800
rect 67450 20788 67456 20800
rect 65208 20760 67456 20788
rect 65208 20748 65214 20760
rect 67450 20748 67456 20760
rect 67508 20748 67514 20800
rect 70366 20788 70394 20828
rect 72694 20816 72700 20868
rect 72752 20856 72758 20868
rect 76650 20856 76656 20868
rect 72752 20828 76656 20856
rect 72752 20816 72758 20828
rect 76650 20816 76656 20828
rect 76708 20816 76714 20868
rect 81728 20788 81756 21023
rect 85574 21020 85580 21032
rect 85632 21020 85638 21072
rect 95329 21063 95387 21069
rect 95329 21029 95341 21063
rect 95375 21060 95387 21063
rect 95878 21060 95884 21072
rect 95375 21032 95884 21060
rect 95375 21029 95387 21032
rect 95329 21023 95387 21029
rect 95878 21020 95884 21032
rect 95936 21020 95942 21072
rect 93578 20952 93584 21004
rect 93636 20992 93642 21004
rect 93949 20995 94007 21001
rect 93949 20992 93961 20995
rect 93636 20964 93961 20992
rect 93636 20952 93642 20964
rect 93949 20961 93961 20964
rect 93995 20992 94007 20995
rect 95421 20995 95479 21001
rect 95421 20992 95433 20995
rect 93995 20964 95433 20992
rect 93995 20961 94007 20964
rect 93949 20955 94007 20961
rect 95421 20961 95433 20964
rect 95467 20992 95479 20995
rect 95605 20995 95663 21001
rect 95605 20992 95617 20995
rect 95467 20964 95617 20992
rect 95467 20961 95479 20964
rect 95421 20955 95479 20961
rect 95605 20961 95617 20964
rect 95651 20992 95663 20995
rect 95789 20995 95847 21001
rect 95789 20992 95801 20995
rect 95651 20964 95801 20992
rect 95651 20961 95663 20964
rect 95605 20955 95663 20961
rect 95789 20961 95801 20964
rect 95835 20992 95847 20995
rect 95973 20995 96031 21001
rect 95973 20992 95985 20995
rect 95835 20964 95985 20992
rect 95835 20961 95847 20964
rect 95789 20955 95847 20961
rect 95973 20961 95985 20964
rect 96019 20992 96031 20995
rect 96157 20995 96215 21001
rect 96157 20992 96169 20995
rect 96019 20964 96169 20992
rect 96019 20961 96031 20964
rect 95973 20955 96031 20961
rect 96157 20961 96169 20964
rect 96203 20961 96215 20995
rect 96157 20955 96215 20961
rect 92934 20884 92940 20936
rect 92992 20924 92998 20936
rect 93673 20927 93731 20933
rect 93673 20924 93685 20927
rect 92992 20896 93685 20924
rect 92992 20884 92998 20896
rect 93673 20893 93685 20896
rect 93719 20893 93731 20927
rect 93673 20887 93731 20893
rect 92750 20788 92756 20800
rect 70366 20760 81756 20788
rect 92711 20760 92756 20788
rect 92750 20748 92756 20760
rect 92808 20788 92814 20800
rect 93121 20791 93179 20797
rect 93121 20788 93133 20791
rect 92808 20760 93133 20788
rect 92808 20748 92814 20760
rect 93121 20757 93133 20760
rect 93167 20788 93179 20791
rect 93305 20791 93363 20797
rect 93305 20788 93317 20791
rect 93167 20760 93317 20788
rect 93167 20757 93179 20760
rect 93121 20751 93179 20757
rect 93305 20757 93317 20760
rect 93351 20788 93363 20791
rect 93489 20791 93547 20797
rect 93489 20788 93501 20791
rect 93351 20760 93501 20788
rect 93351 20757 93363 20760
rect 93305 20751 93363 20757
rect 93489 20757 93501 20760
rect 93535 20788 93547 20791
rect 93578 20788 93584 20800
rect 93535 20760 93584 20788
rect 93535 20757 93547 20760
rect 93489 20751 93547 20757
rect 93578 20748 93584 20760
rect 93636 20748 93642 20800
rect 1104 20698 98808 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 65686 20698
rect 65738 20646 65750 20698
rect 65802 20646 65814 20698
rect 65866 20646 65878 20698
rect 65930 20646 96406 20698
rect 96458 20646 96470 20698
rect 96522 20646 96534 20698
rect 96586 20646 96598 20698
rect 96650 20646 98808 20698
rect 1104 20624 98808 20646
rect 2958 20544 2964 20596
rect 3016 20584 3022 20596
rect 22462 20584 22468 20596
rect 3016 20556 22468 20584
rect 3016 20544 3022 20556
rect 22462 20544 22468 20556
rect 22520 20544 22526 20596
rect 22738 20544 22744 20596
rect 22796 20584 22802 20596
rect 22796 20556 22841 20584
rect 22796 20544 22802 20556
rect 23014 20544 23020 20596
rect 23072 20584 23078 20596
rect 44082 20584 44088 20596
rect 23072 20556 44088 20584
rect 23072 20544 23078 20556
rect 44082 20544 44088 20556
rect 44140 20544 44146 20596
rect 44634 20544 44640 20596
rect 44692 20584 44698 20596
rect 46106 20584 46112 20596
rect 44692 20556 46112 20584
rect 44692 20544 44698 20556
rect 46106 20544 46112 20556
rect 46164 20544 46170 20596
rect 46223 20556 46428 20584
rect 16850 20476 16856 20528
rect 16908 20516 16914 20528
rect 46223 20516 46251 20556
rect 16908 20488 46251 20516
rect 46400 20516 46428 20556
rect 51902 20544 51908 20596
rect 51960 20584 51966 20596
rect 53926 20584 53932 20596
rect 51960 20556 53932 20584
rect 51960 20544 51966 20556
rect 53926 20544 53932 20556
rect 53984 20544 53990 20596
rect 54018 20544 54024 20596
rect 54076 20584 54082 20596
rect 81618 20584 81624 20596
rect 54076 20556 81624 20584
rect 54076 20544 54082 20556
rect 81618 20544 81624 20556
rect 81676 20544 81682 20596
rect 93302 20544 93308 20596
rect 93360 20584 93366 20596
rect 94225 20587 94283 20593
rect 94225 20584 94237 20587
rect 93360 20556 94237 20584
rect 93360 20544 93366 20556
rect 94225 20553 94237 20556
rect 94271 20553 94283 20587
rect 94225 20547 94283 20553
rect 64506 20516 64512 20528
rect 46400 20488 64512 20516
rect 16908 20476 16914 20488
rect 64506 20476 64512 20488
rect 64564 20476 64570 20528
rect 70578 20516 70584 20528
rect 65536 20488 70440 20516
rect 70539 20488 70584 20516
rect 5534 20408 5540 20460
rect 5592 20448 5598 20460
rect 6270 20448 6276 20460
rect 5592 20420 6276 20448
rect 5592 20408 5598 20420
rect 6270 20408 6276 20420
rect 6328 20448 6334 20460
rect 22462 20448 22468 20460
rect 6328 20420 22468 20448
rect 6328 20408 6334 20420
rect 22462 20408 22468 20420
rect 22520 20408 22526 20460
rect 23014 20408 23020 20460
rect 23072 20448 23078 20460
rect 33686 20448 33692 20460
rect 23072 20420 33692 20448
rect 23072 20408 23078 20420
rect 33686 20408 33692 20420
rect 33744 20408 33750 20460
rect 33796 20420 45416 20448
rect 15657 20383 15715 20389
rect 15657 20349 15669 20383
rect 15703 20380 15715 20383
rect 33796 20380 33824 20420
rect 15703 20352 33824 20380
rect 34241 20383 34299 20389
rect 15703 20349 15715 20352
rect 15657 20343 15715 20349
rect 34241 20349 34253 20383
rect 34287 20349 34299 20383
rect 34241 20343 34299 20349
rect 15838 20272 15844 20324
rect 15896 20312 15902 20324
rect 34054 20312 34060 20324
rect 15896 20284 34060 20312
rect 15896 20272 15902 20284
rect 34054 20272 34060 20284
rect 34112 20272 34118 20324
rect 12802 20204 12808 20256
rect 12860 20244 12866 20256
rect 23198 20244 23204 20256
rect 12860 20216 23204 20244
rect 12860 20204 12866 20216
rect 23198 20204 23204 20216
rect 23256 20204 23262 20256
rect 26602 20204 26608 20256
rect 26660 20244 26666 20256
rect 27154 20244 27160 20256
rect 26660 20216 27160 20244
rect 26660 20204 26666 20216
rect 27154 20204 27160 20216
rect 27212 20204 27218 20256
rect 27246 20204 27252 20256
rect 27304 20244 27310 20256
rect 34146 20244 34152 20256
rect 27304 20216 34152 20244
rect 27304 20204 27310 20216
rect 34146 20204 34152 20216
rect 34204 20204 34210 20256
rect 34256 20244 34284 20343
rect 38838 20340 38844 20392
rect 38896 20380 38902 20392
rect 39022 20380 39028 20392
rect 38896 20352 39028 20380
rect 38896 20340 38902 20352
rect 39022 20340 39028 20352
rect 39080 20340 39086 20392
rect 45278 20380 45284 20392
rect 41386 20352 45284 20380
rect 34698 20272 34704 20324
rect 34756 20312 34762 20324
rect 41386 20312 41414 20352
rect 45278 20340 45284 20352
rect 45336 20340 45342 20392
rect 34756 20284 41414 20312
rect 45388 20312 45416 20420
rect 46934 20408 46940 20460
rect 46992 20448 46998 20460
rect 52270 20448 52276 20460
rect 46992 20420 52276 20448
rect 46992 20408 46998 20420
rect 52270 20408 52276 20420
rect 52328 20408 52334 20460
rect 53098 20408 53104 20460
rect 53156 20448 53162 20460
rect 53156 20420 54248 20448
rect 53156 20408 53162 20420
rect 45462 20340 45468 20392
rect 45520 20380 45526 20392
rect 51902 20380 51908 20392
rect 45520 20352 51908 20380
rect 45520 20340 45526 20352
rect 51902 20340 51908 20352
rect 51960 20380 51966 20392
rect 51997 20383 52055 20389
rect 51997 20380 52009 20383
rect 51960 20352 52009 20380
rect 51960 20340 51966 20352
rect 51997 20349 52009 20352
rect 52043 20349 52055 20383
rect 54110 20380 54116 20392
rect 51997 20343 52055 20349
rect 52196 20352 54116 20380
rect 52196 20312 52224 20352
rect 54110 20340 54116 20352
rect 54168 20340 54174 20392
rect 54220 20380 54248 20420
rect 54478 20408 54484 20460
rect 54536 20448 54542 20460
rect 58894 20448 58900 20460
rect 54536 20420 58900 20448
rect 54536 20408 54542 20420
rect 58894 20408 58900 20420
rect 58952 20448 58958 20460
rect 59722 20448 59728 20460
rect 58952 20420 59728 20448
rect 58952 20408 58958 20420
rect 59722 20408 59728 20420
rect 59780 20408 59786 20460
rect 62758 20408 62764 20460
rect 62816 20448 62822 20460
rect 63678 20448 63684 20460
rect 62816 20420 63684 20448
rect 62816 20408 62822 20420
rect 63678 20408 63684 20420
rect 63736 20408 63742 20460
rect 63954 20380 63960 20392
rect 54220 20352 63960 20380
rect 63954 20340 63960 20352
rect 64012 20340 64018 20392
rect 64509 20383 64567 20389
rect 64509 20349 64521 20383
rect 64555 20380 64567 20383
rect 65150 20380 65156 20392
rect 64555 20352 65156 20380
rect 64555 20349 64567 20352
rect 64509 20343 64567 20349
rect 65150 20340 65156 20352
rect 65208 20340 65214 20392
rect 65242 20340 65248 20392
rect 65300 20380 65306 20392
rect 65536 20380 65564 20488
rect 70210 20448 70216 20460
rect 70171 20420 70216 20448
rect 70210 20408 70216 20420
rect 70268 20408 70274 20460
rect 70412 20448 70440 20488
rect 70578 20476 70584 20488
rect 70636 20476 70642 20528
rect 71409 20519 71467 20525
rect 71409 20485 71421 20519
rect 71455 20516 71467 20519
rect 71774 20516 71780 20528
rect 71455 20488 71780 20516
rect 71455 20485 71467 20488
rect 71409 20479 71467 20485
rect 71774 20476 71780 20488
rect 71832 20476 71838 20528
rect 73154 20516 73160 20528
rect 71884 20488 73160 20516
rect 71884 20448 71912 20488
rect 73154 20476 73160 20488
rect 73212 20476 73218 20528
rect 81710 20516 81716 20528
rect 75288 20488 81716 20516
rect 72694 20448 72700 20460
rect 70412 20420 71912 20448
rect 72655 20420 72700 20448
rect 72694 20408 72700 20420
rect 72752 20408 72758 20460
rect 73062 20408 73068 20460
rect 73120 20448 73126 20460
rect 75288 20448 75316 20488
rect 81710 20476 81716 20488
rect 81768 20476 81774 20528
rect 81894 20476 81900 20528
rect 81952 20516 81958 20528
rect 93946 20516 93952 20528
rect 81952 20488 93952 20516
rect 81952 20476 81958 20488
rect 93946 20476 93952 20488
rect 94004 20476 94010 20528
rect 94590 20476 94596 20528
rect 94648 20516 94654 20528
rect 95142 20516 95148 20528
rect 94648 20488 95148 20516
rect 94648 20476 94654 20488
rect 95142 20476 95148 20488
rect 95200 20516 95206 20528
rect 95200 20488 97488 20516
rect 95200 20476 95206 20488
rect 80974 20448 80980 20460
rect 73120 20420 75316 20448
rect 80026 20420 80980 20448
rect 73120 20408 73126 20420
rect 65300 20352 65564 20380
rect 65300 20340 65306 20352
rect 69750 20340 69756 20392
rect 69808 20380 69814 20392
rect 69845 20383 69903 20389
rect 69845 20380 69857 20383
rect 69808 20352 69857 20380
rect 69808 20340 69814 20352
rect 69845 20349 69857 20352
rect 69891 20349 69903 20383
rect 69845 20343 69903 20349
rect 69934 20340 69940 20392
rect 69992 20389 69998 20392
rect 69992 20383 70051 20389
rect 69992 20349 70005 20383
rect 70039 20349 70051 20383
rect 70118 20380 70124 20392
rect 70079 20352 70124 20380
rect 69992 20343 70051 20349
rect 69992 20340 69998 20343
rect 70118 20340 70124 20352
rect 70176 20340 70182 20392
rect 70397 20383 70455 20389
rect 70397 20349 70409 20383
rect 70443 20380 70455 20383
rect 70762 20380 70768 20392
rect 70443 20352 70768 20380
rect 70443 20349 70455 20352
rect 70397 20343 70455 20349
rect 70762 20340 70768 20352
rect 70820 20340 70826 20392
rect 71130 20340 71136 20392
rect 71188 20380 71194 20392
rect 71961 20383 72019 20389
rect 71961 20380 71973 20383
rect 71188 20352 71973 20380
rect 71188 20340 71194 20352
rect 71961 20349 71973 20352
rect 72007 20349 72019 20383
rect 72142 20380 72148 20392
rect 72103 20352 72148 20380
rect 71961 20343 72019 20349
rect 72142 20340 72148 20352
rect 72200 20340 72206 20392
rect 72513 20383 72571 20389
rect 72513 20349 72525 20383
rect 72559 20380 72571 20383
rect 72602 20380 72608 20392
rect 72559 20352 72608 20380
rect 72559 20349 72571 20352
rect 72513 20343 72571 20349
rect 72602 20340 72608 20352
rect 72660 20340 72666 20392
rect 72878 20380 72884 20392
rect 72839 20352 72884 20380
rect 72878 20340 72884 20352
rect 72936 20340 72942 20392
rect 72970 20340 72976 20392
rect 73028 20380 73034 20392
rect 80026 20380 80054 20420
rect 80974 20408 80980 20420
rect 81032 20408 81038 20460
rect 82262 20408 82268 20460
rect 82320 20448 82326 20460
rect 97460 20457 97488 20488
rect 97445 20451 97503 20457
rect 82320 20420 97120 20448
rect 82320 20408 82326 20420
rect 73028 20352 80054 20380
rect 73028 20340 73034 20352
rect 81526 20340 81532 20392
rect 81584 20380 81590 20392
rect 81621 20383 81679 20389
rect 81621 20380 81633 20383
rect 81584 20352 81633 20380
rect 81584 20340 81590 20352
rect 81621 20349 81633 20352
rect 81667 20349 81679 20383
rect 81621 20343 81679 20349
rect 81710 20340 81716 20392
rect 81768 20380 81774 20392
rect 81805 20383 81863 20389
rect 81805 20380 81817 20383
rect 81768 20352 81817 20380
rect 81768 20340 81774 20352
rect 81805 20349 81817 20352
rect 81851 20349 81863 20383
rect 81805 20343 81863 20349
rect 81894 20340 81900 20392
rect 81952 20389 81958 20392
rect 81952 20383 82001 20389
rect 81952 20349 81955 20383
rect 81989 20349 82001 20383
rect 82078 20380 82084 20392
rect 82039 20352 82084 20380
rect 81952 20343 82001 20349
rect 81952 20340 81958 20343
rect 82078 20340 82084 20352
rect 82136 20340 82142 20392
rect 82170 20340 82176 20392
rect 82228 20380 82234 20392
rect 82354 20380 82360 20392
rect 82228 20352 82273 20380
rect 82315 20352 82360 20380
rect 82228 20340 82234 20352
rect 82354 20340 82360 20352
rect 82412 20340 82418 20392
rect 89530 20340 89536 20392
rect 89588 20380 89594 20392
rect 93489 20383 93547 20389
rect 93489 20380 93501 20383
rect 89588 20352 93501 20380
rect 89588 20340 89594 20352
rect 93489 20349 93501 20352
rect 93535 20349 93547 20383
rect 93670 20380 93676 20392
rect 93631 20352 93676 20380
rect 93489 20343 93547 20349
rect 93670 20340 93676 20352
rect 93728 20340 93734 20392
rect 93946 20389 93952 20392
rect 93774 20383 93832 20389
rect 93774 20349 93786 20383
rect 93820 20380 93832 20383
rect 93903 20383 93952 20389
rect 93820 20349 93854 20380
rect 93774 20343 93854 20349
rect 93903 20349 93915 20383
rect 93949 20349 93952 20383
rect 93903 20343 93952 20349
rect 45388 20284 52224 20312
rect 34756 20272 34762 20284
rect 52270 20272 52276 20324
rect 52328 20312 52334 20324
rect 52328 20284 52373 20312
rect 52328 20272 52334 20284
rect 52454 20272 52460 20324
rect 52512 20312 52518 20324
rect 53926 20312 53932 20324
rect 52512 20284 53932 20312
rect 52512 20272 52518 20284
rect 53926 20272 53932 20284
rect 53984 20272 53990 20324
rect 64782 20321 64788 20324
rect 64776 20312 64788 20321
rect 54036 20284 64184 20312
rect 64743 20284 64788 20312
rect 44634 20244 44640 20256
rect 34256 20216 44640 20244
rect 44634 20204 44640 20216
rect 44692 20204 44698 20256
rect 45094 20204 45100 20256
rect 45152 20244 45158 20256
rect 45278 20244 45284 20256
rect 45152 20216 45284 20244
rect 45152 20204 45158 20216
rect 45278 20204 45284 20216
rect 45336 20204 45342 20256
rect 46205 20204 46211 20256
rect 46263 20244 46269 20256
rect 54036 20244 54064 20284
rect 46263 20216 54064 20244
rect 46263 20204 46269 20216
rect 54110 20204 54116 20256
rect 54168 20244 54174 20256
rect 64046 20244 64052 20256
rect 54168 20216 64052 20244
rect 54168 20204 54174 20216
rect 64046 20204 64052 20216
rect 64104 20204 64110 20256
rect 64156 20244 64184 20284
rect 64776 20275 64788 20284
rect 64782 20272 64788 20275
rect 64840 20272 64846 20324
rect 79042 20312 79048 20324
rect 64892 20284 79048 20312
rect 64892 20244 64920 20284
rect 79042 20272 79048 20284
rect 79100 20272 79106 20324
rect 81360 20284 81940 20312
rect 64156 20216 64920 20244
rect 65058 20204 65064 20256
rect 65116 20244 65122 20256
rect 65889 20247 65947 20253
rect 65889 20244 65901 20247
rect 65116 20216 65901 20244
rect 65116 20204 65122 20216
rect 65889 20213 65901 20216
rect 65935 20213 65947 20247
rect 65889 20207 65947 20213
rect 65978 20204 65984 20256
rect 66036 20244 66042 20256
rect 70854 20244 70860 20256
rect 66036 20216 70860 20244
rect 66036 20204 66042 20216
rect 70854 20204 70860 20216
rect 70912 20244 70918 20256
rect 71130 20244 71136 20256
rect 70912 20216 71136 20244
rect 70912 20204 70918 20216
rect 71130 20204 71136 20216
rect 71188 20204 71194 20256
rect 71774 20204 71780 20256
rect 71832 20244 71838 20256
rect 72973 20247 73031 20253
rect 72973 20244 72985 20247
rect 71832 20216 72985 20244
rect 71832 20204 71838 20216
rect 72973 20213 72985 20216
rect 73019 20213 73031 20247
rect 72973 20207 73031 20213
rect 73154 20204 73160 20256
rect 73212 20244 73218 20256
rect 81360 20244 81388 20284
rect 73212 20216 81388 20244
rect 81437 20247 81495 20253
rect 73212 20204 73218 20216
rect 81437 20213 81449 20247
rect 81483 20244 81495 20247
rect 81802 20244 81808 20256
rect 81483 20216 81808 20244
rect 81483 20213 81495 20216
rect 81437 20207 81495 20213
rect 81802 20204 81808 20216
rect 81860 20204 81866 20256
rect 81912 20244 81940 20284
rect 92842 20272 92848 20324
rect 92900 20312 92906 20324
rect 93826 20312 93854 20343
rect 93946 20340 93952 20343
rect 94004 20340 94010 20392
rect 97092 20389 97120 20420
rect 97445 20417 97457 20451
rect 97491 20417 97503 20451
rect 97445 20411 97503 20417
rect 94041 20383 94099 20389
rect 94041 20349 94053 20383
rect 94087 20349 94099 20383
rect 94041 20343 94099 20349
rect 97077 20383 97135 20389
rect 97077 20349 97089 20383
rect 97123 20349 97135 20383
rect 97077 20343 97135 20349
rect 92900 20284 93854 20312
rect 92900 20272 92906 20284
rect 92290 20244 92296 20256
rect 81912 20216 92296 20244
rect 92290 20204 92296 20216
rect 92348 20204 92354 20256
rect 92658 20204 92664 20256
rect 92716 20244 92722 20256
rect 94056 20244 94084 20343
rect 92716 20216 94084 20244
rect 92716 20204 92722 20216
rect 1104 20154 98808 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 50326 20154
rect 50378 20102 50390 20154
rect 50442 20102 50454 20154
rect 50506 20102 50518 20154
rect 50570 20102 81046 20154
rect 81098 20102 81110 20154
rect 81162 20102 81174 20154
rect 81226 20102 81238 20154
rect 81290 20102 98808 20154
rect 1104 20080 98808 20102
rect 3234 20000 3240 20052
rect 3292 20040 3298 20052
rect 34054 20040 34060 20052
rect 3292 20012 34060 20040
rect 3292 20000 3298 20012
rect 34054 20000 34060 20012
rect 34112 20000 34118 20052
rect 34146 20000 34152 20052
rect 34204 20040 34210 20052
rect 38289 20043 38347 20049
rect 38289 20040 38301 20043
rect 34204 20012 38301 20040
rect 34204 20000 34210 20012
rect 38289 20009 38301 20012
rect 38335 20009 38347 20043
rect 38289 20003 38347 20009
rect 38473 20043 38531 20049
rect 38473 20009 38485 20043
rect 38519 20009 38531 20043
rect 38473 20003 38531 20009
rect 3786 19932 3792 19984
rect 3844 19972 3850 19984
rect 19242 19972 19248 19984
rect 3844 19944 19248 19972
rect 3844 19932 3850 19944
rect 19242 19932 19248 19944
rect 19300 19932 19306 19984
rect 33686 19972 33692 19984
rect 22066 19944 33692 19972
rect 1394 19904 1400 19916
rect 1355 19876 1400 19904
rect 1394 19864 1400 19876
rect 1452 19864 1458 19916
rect 9398 19864 9404 19916
rect 9456 19904 9462 19916
rect 18138 19904 18144 19916
rect 9456 19876 18144 19904
rect 9456 19864 9462 19876
rect 18138 19864 18144 19876
rect 18196 19864 18202 19916
rect 20162 19796 20168 19848
rect 20220 19836 20226 19848
rect 22066 19836 22094 19944
rect 33686 19932 33692 19944
rect 33744 19932 33750 19984
rect 26418 19864 26424 19916
rect 26476 19904 26482 19916
rect 26878 19904 26884 19916
rect 26476 19876 26884 19904
rect 26476 19864 26482 19876
rect 26878 19864 26884 19876
rect 26936 19864 26942 19916
rect 27246 19864 27252 19916
rect 27304 19904 27310 19916
rect 27522 19904 27528 19916
rect 27304 19876 27528 19904
rect 27304 19864 27310 19876
rect 27522 19864 27528 19876
rect 27580 19904 27586 19916
rect 28813 19907 28871 19913
rect 28813 19904 28825 19907
rect 27580 19876 28825 19904
rect 27580 19864 27586 19876
rect 28813 19873 28825 19876
rect 28859 19873 28871 19907
rect 33413 19907 33471 19913
rect 28813 19867 28871 19873
rect 28920 19876 31754 19904
rect 20220 19808 22094 19836
rect 20220 19796 20226 19808
rect 26970 19796 26976 19848
rect 27028 19836 27034 19848
rect 28920 19836 28948 19876
rect 29086 19836 29092 19848
rect 27028 19808 28948 19836
rect 29047 19808 29092 19836
rect 27028 19796 27034 19808
rect 29086 19796 29092 19808
rect 29144 19796 29150 19848
rect 31726 19836 31754 19876
rect 33413 19873 33425 19907
rect 33459 19904 33471 19907
rect 38488 19904 38516 20003
rect 38562 20000 38568 20052
rect 38620 20040 38626 20052
rect 38620 20012 38792 20040
rect 38620 20000 38626 20012
rect 38764 19972 38792 20012
rect 44082 20000 44088 20052
rect 44140 20040 44146 20052
rect 48314 20040 48320 20052
rect 44140 20012 48320 20040
rect 44140 20000 44146 20012
rect 48314 20000 48320 20012
rect 48372 20000 48378 20052
rect 48590 20000 48596 20052
rect 48648 20040 48654 20052
rect 78674 20040 78680 20052
rect 48648 20012 78680 20040
rect 48648 20000 48654 20012
rect 78674 20000 78680 20012
rect 78732 20040 78738 20052
rect 91830 20040 91836 20052
rect 78732 20012 91836 20040
rect 78732 20000 78738 20012
rect 91830 20000 91836 20012
rect 91888 20000 91894 20052
rect 97626 20040 97632 20052
rect 97587 20012 97632 20040
rect 97626 20000 97632 20012
rect 97684 20000 97690 20052
rect 38764 19944 54156 19972
rect 33459 19876 38516 19904
rect 38657 19907 38715 19913
rect 33459 19873 33471 19876
rect 33413 19867 33471 19873
rect 38657 19873 38669 19907
rect 38703 19904 38715 19907
rect 38746 19904 38752 19916
rect 38703 19876 38752 19904
rect 38703 19873 38715 19876
rect 38657 19867 38715 19873
rect 38746 19864 38752 19876
rect 38804 19864 38810 19916
rect 45462 19904 45468 19916
rect 38856 19876 45468 19904
rect 38289 19839 38347 19845
rect 38289 19836 38301 19839
rect 31726 19808 38301 19836
rect 38289 19805 38301 19808
rect 38335 19805 38347 19839
rect 38289 19799 38347 19805
rect 38381 19839 38439 19845
rect 38381 19805 38393 19839
rect 38427 19836 38439 19839
rect 38856 19836 38884 19876
rect 45462 19864 45468 19876
rect 45520 19864 45526 19916
rect 46934 19864 46940 19916
rect 46992 19904 46998 19916
rect 48314 19904 48320 19916
rect 46992 19876 48320 19904
rect 46992 19864 46998 19876
rect 48314 19864 48320 19876
rect 48372 19864 48378 19916
rect 48774 19904 48780 19916
rect 48735 19876 48780 19904
rect 48774 19864 48780 19876
rect 48832 19864 48838 19916
rect 54128 19904 54156 19944
rect 54202 19932 54208 19984
rect 54260 19972 54266 19984
rect 54849 19975 54907 19981
rect 54849 19972 54861 19975
rect 54260 19944 54861 19972
rect 54260 19932 54266 19944
rect 54849 19941 54861 19944
rect 54895 19941 54907 19975
rect 54849 19935 54907 19941
rect 54941 19975 54999 19981
rect 54941 19941 54953 19975
rect 54987 19972 54999 19975
rect 56594 19972 56600 19984
rect 54987 19944 56600 19972
rect 54987 19941 54999 19944
rect 54941 19935 54999 19941
rect 56594 19932 56600 19944
rect 56652 19932 56658 19984
rect 56704 19944 59676 19972
rect 54478 19904 54484 19916
rect 54128 19876 54484 19904
rect 54478 19864 54484 19876
rect 54536 19864 54542 19916
rect 54662 19904 54668 19916
rect 54623 19876 54668 19904
rect 54662 19864 54668 19876
rect 54720 19864 54726 19916
rect 55033 19907 55091 19913
rect 55033 19873 55045 19907
rect 55079 19904 55091 19907
rect 55122 19904 55128 19916
rect 55079 19876 55128 19904
rect 55079 19873 55091 19876
rect 55033 19867 55091 19873
rect 55122 19864 55128 19876
rect 55180 19864 55186 19916
rect 55674 19864 55680 19916
rect 55732 19904 55738 19916
rect 56704 19904 56732 19944
rect 55732 19876 56732 19904
rect 59449 19907 59507 19913
rect 55732 19864 55738 19876
rect 59449 19873 59461 19907
rect 59495 19873 59507 19907
rect 59648 19904 59676 19944
rect 59722 19932 59728 19984
rect 59780 19972 59786 19984
rect 59780 19944 70394 19972
rect 59780 19932 59786 19944
rect 61746 19904 61752 19916
rect 59648 19876 61752 19904
rect 59449 19867 59507 19873
rect 38427 19808 38884 19836
rect 38427 19805 38439 19808
rect 38381 19799 38439 19805
rect 43438 19796 43444 19848
rect 43496 19836 43502 19848
rect 50525 19839 50583 19845
rect 43496 19808 48314 19836
rect 43496 19796 43502 19808
rect 12066 19728 12072 19780
rect 12124 19768 12130 19780
rect 36262 19768 36268 19780
rect 12124 19740 36268 19768
rect 12124 19728 12130 19740
rect 36262 19728 36268 19740
rect 36320 19728 36326 19780
rect 38654 19768 38660 19780
rect 38212 19740 38660 19768
rect 27154 19660 27160 19712
rect 27212 19700 27218 19712
rect 33229 19703 33287 19709
rect 33229 19700 33241 19703
rect 27212 19672 33241 19700
rect 27212 19660 27218 19672
rect 33229 19669 33241 19672
rect 33275 19669 33287 19703
rect 33229 19663 33287 19669
rect 34790 19660 34796 19712
rect 34848 19700 34854 19712
rect 38212 19700 38240 19740
rect 38654 19728 38660 19740
rect 38712 19728 38718 19780
rect 39022 19728 39028 19780
rect 39080 19768 39086 19780
rect 46198 19768 46204 19780
rect 39080 19740 46204 19768
rect 39080 19728 39086 19740
rect 46198 19728 46204 19740
rect 46256 19728 46262 19780
rect 46290 19728 46296 19780
rect 46348 19768 46354 19780
rect 47762 19768 47768 19780
rect 46348 19740 47768 19768
rect 46348 19728 46354 19740
rect 47762 19728 47768 19740
rect 47820 19728 47826 19780
rect 48286 19768 48314 19808
rect 50525 19805 50537 19839
rect 50571 19836 50583 19839
rect 59464 19836 59492 19867
rect 61746 19864 61752 19876
rect 61804 19864 61810 19916
rect 64601 19907 64659 19913
rect 64601 19904 64613 19907
rect 61948 19876 64613 19904
rect 50571 19808 59492 19836
rect 50571 19805 50583 19808
rect 50525 19799 50583 19805
rect 50540 19768 50568 19799
rect 48286 19740 50568 19768
rect 53466 19728 53472 19780
rect 53524 19768 53530 19780
rect 55217 19771 55275 19777
rect 55217 19768 55229 19771
rect 53524 19740 55229 19768
rect 53524 19728 53530 19740
rect 55217 19737 55229 19740
rect 55263 19737 55275 19771
rect 55217 19731 55275 19737
rect 59265 19771 59323 19777
rect 59265 19737 59277 19771
rect 59311 19768 59323 19771
rect 61948 19768 61976 19876
rect 64601 19873 64613 19876
rect 64647 19873 64659 19907
rect 64601 19867 64659 19873
rect 62942 19796 62948 19848
rect 63000 19836 63006 19848
rect 63218 19836 63224 19848
rect 63000 19808 63224 19836
rect 63000 19796 63006 19808
rect 63218 19796 63224 19808
rect 63276 19796 63282 19848
rect 70366 19836 70394 19944
rect 73062 19932 73068 19984
rect 73120 19972 73126 19984
rect 97353 19975 97411 19981
rect 73120 19944 80054 19972
rect 73120 19932 73126 19944
rect 73982 19904 73988 19916
rect 73943 19876 73988 19904
rect 73982 19864 73988 19876
rect 74040 19904 74046 19916
rect 74626 19904 74632 19916
rect 74040 19876 74632 19904
rect 74040 19864 74046 19876
rect 74626 19864 74632 19876
rect 74684 19864 74690 19916
rect 75638 19904 75644 19916
rect 75599 19876 75644 19904
rect 75638 19864 75644 19876
rect 75696 19864 75702 19916
rect 75822 19904 75828 19916
rect 75783 19876 75828 19904
rect 75822 19864 75828 19876
rect 75880 19864 75886 19916
rect 80026 19904 80054 19944
rect 97353 19941 97365 19975
rect 97399 19972 97411 19975
rect 97534 19972 97540 19984
rect 97399 19944 97540 19972
rect 97399 19941 97411 19944
rect 97353 19935 97411 19941
rect 97534 19932 97540 19944
rect 97592 19932 97598 19984
rect 86954 19904 86960 19916
rect 80026 19876 86960 19904
rect 86954 19864 86960 19876
rect 87012 19864 87018 19916
rect 74721 19839 74779 19845
rect 74721 19836 74733 19839
rect 70366 19808 74733 19836
rect 74721 19805 74733 19808
rect 74767 19805 74779 19839
rect 74721 19799 74779 19805
rect 76193 19839 76251 19845
rect 76193 19805 76205 19839
rect 76239 19836 76251 19839
rect 76282 19836 76288 19848
rect 76239 19808 76288 19836
rect 76239 19805 76251 19808
rect 76193 19799 76251 19805
rect 76282 19796 76288 19808
rect 76340 19796 76346 19848
rect 59311 19740 61976 19768
rect 59311 19737 59323 19740
rect 59265 19731 59323 19737
rect 63954 19728 63960 19780
rect 64012 19768 64018 19780
rect 87690 19768 87696 19780
rect 64012 19740 87696 19768
rect 64012 19728 64018 19740
rect 87690 19728 87696 19740
rect 87748 19728 87754 19780
rect 34848 19672 38240 19700
rect 38289 19703 38347 19709
rect 34848 19660 34854 19672
rect 38289 19669 38301 19703
rect 38335 19700 38347 19703
rect 43898 19700 43904 19712
rect 38335 19672 43904 19700
rect 38335 19669 38347 19672
rect 38289 19663 38347 19669
rect 43898 19660 43904 19672
rect 43956 19660 43962 19712
rect 43990 19660 43996 19712
rect 44048 19700 44054 19712
rect 50154 19700 50160 19712
rect 44048 19672 50160 19700
rect 44048 19660 44054 19672
rect 50154 19660 50160 19672
rect 50212 19660 50218 19712
rect 55030 19660 55036 19712
rect 55088 19700 55094 19712
rect 57514 19700 57520 19712
rect 55088 19672 57520 19700
rect 55088 19660 55094 19672
rect 57514 19660 57520 19672
rect 57572 19660 57578 19712
rect 59354 19660 59360 19712
rect 59412 19700 59418 19712
rect 60918 19700 60924 19712
rect 59412 19672 60924 19700
rect 59412 19660 59418 19672
rect 60918 19660 60924 19672
rect 60976 19660 60982 19712
rect 61102 19660 61108 19712
rect 61160 19700 61166 19712
rect 63770 19700 63776 19712
rect 61160 19672 63776 19700
rect 61160 19660 61166 19672
rect 63770 19660 63776 19672
rect 63828 19660 63834 19712
rect 64417 19703 64475 19709
rect 64417 19669 64429 19703
rect 64463 19700 64475 19703
rect 71222 19700 71228 19712
rect 64463 19672 71228 19700
rect 64463 19669 64475 19672
rect 64417 19663 64475 19669
rect 71222 19660 71228 19672
rect 71280 19700 71286 19712
rect 71682 19700 71688 19712
rect 71280 19672 71688 19700
rect 71280 19660 71286 19672
rect 71682 19660 71688 19672
rect 71740 19660 71746 19712
rect 71774 19660 71780 19712
rect 71832 19700 71838 19712
rect 75730 19700 75736 19712
rect 71832 19672 75736 19700
rect 71832 19660 71838 19672
rect 75730 19660 75736 19672
rect 75788 19660 75794 19712
rect 1104 19610 98808 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 65686 19610
rect 65738 19558 65750 19610
rect 65802 19558 65814 19610
rect 65866 19558 65878 19610
rect 65930 19558 96406 19610
rect 96458 19558 96470 19610
rect 96522 19558 96534 19610
rect 96586 19558 96598 19610
rect 96650 19558 98808 19610
rect 1104 19536 98808 19558
rect 21910 19456 21916 19508
rect 21968 19496 21974 19508
rect 50065 19499 50123 19505
rect 50065 19496 50077 19499
rect 21968 19468 50077 19496
rect 21968 19456 21974 19468
rect 50065 19465 50077 19468
rect 50111 19496 50123 19499
rect 50430 19496 50436 19508
rect 50111 19468 50436 19496
rect 50111 19465 50123 19468
rect 50065 19459 50123 19465
rect 50430 19456 50436 19468
rect 50488 19456 50494 19508
rect 52270 19456 52276 19508
rect 52328 19496 52334 19508
rect 73982 19496 73988 19508
rect 52328 19468 73988 19496
rect 52328 19456 52334 19468
rect 73982 19456 73988 19468
rect 74040 19456 74046 19508
rect 18046 19388 18052 19440
rect 18104 19428 18110 19440
rect 34790 19428 34796 19440
rect 18104 19400 34796 19428
rect 18104 19388 18110 19400
rect 34790 19388 34796 19400
rect 34848 19388 34854 19440
rect 34882 19388 34888 19440
rect 34940 19428 34946 19440
rect 34940 19400 36216 19428
rect 34940 19388 34946 19400
rect 6730 19320 6736 19372
rect 6788 19360 6794 19372
rect 33686 19360 33692 19372
rect 6788 19332 33692 19360
rect 6788 19320 6794 19332
rect 33686 19320 33692 19332
rect 33744 19320 33750 19372
rect 4982 19252 4988 19304
rect 5040 19292 5046 19304
rect 27338 19292 27344 19304
rect 5040 19264 27344 19292
rect 5040 19252 5046 19264
rect 27338 19252 27344 19264
rect 27396 19252 27402 19304
rect 35894 19292 35900 19304
rect 35855 19264 35900 19292
rect 35894 19252 35900 19264
rect 35952 19252 35958 19304
rect 36078 19292 36084 19304
rect 36039 19264 36084 19292
rect 36078 19252 36084 19264
rect 36136 19252 36142 19304
rect 36188 19301 36216 19400
rect 36262 19388 36268 19440
rect 36320 19428 36326 19440
rect 44082 19428 44088 19440
rect 36320 19400 44088 19428
rect 36320 19388 36326 19400
rect 44082 19388 44088 19400
rect 44140 19388 44146 19440
rect 45094 19428 45100 19440
rect 44284 19400 45100 19428
rect 36630 19320 36636 19372
rect 36688 19360 36694 19372
rect 44284 19360 44312 19400
rect 45094 19388 45100 19400
rect 45152 19388 45158 19440
rect 46106 19388 46112 19440
rect 46164 19428 46170 19440
rect 47854 19428 47860 19440
rect 46164 19400 47860 19428
rect 46164 19388 46170 19400
rect 47854 19388 47860 19400
rect 47912 19388 47918 19440
rect 49329 19431 49387 19437
rect 49329 19397 49341 19431
rect 49375 19428 49387 19431
rect 49375 19400 52592 19428
rect 49375 19397 49387 19400
rect 49329 19391 49387 19397
rect 36688 19332 44312 19360
rect 44361 19363 44419 19369
rect 36688 19320 36694 19332
rect 44361 19329 44373 19363
rect 44407 19360 44419 19363
rect 44407 19332 45324 19360
rect 44407 19329 44419 19332
rect 44361 19323 44419 19329
rect 36354 19301 36360 19304
rect 36173 19295 36231 19301
rect 36173 19261 36185 19295
rect 36219 19261 36231 19295
rect 36173 19255 36231 19261
rect 36311 19295 36360 19301
rect 36311 19261 36323 19295
rect 36357 19261 36360 19295
rect 36311 19255 36360 19261
rect 36354 19252 36360 19255
rect 36412 19252 36418 19304
rect 36449 19295 36507 19301
rect 36449 19261 36461 19295
rect 36495 19292 36507 19295
rect 36538 19292 36544 19304
rect 36495 19264 36544 19292
rect 36495 19261 36507 19264
rect 36449 19255 36507 19261
rect 36538 19252 36544 19264
rect 36596 19252 36602 19304
rect 36906 19252 36912 19304
rect 36964 19292 36970 19304
rect 45296 19292 45324 19332
rect 45462 19320 45468 19372
rect 45520 19360 45526 19372
rect 48590 19360 48596 19372
rect 45520 19332 48596 19360
rect 45520 19320 45526 19332
rect 48590 19320 48596 19332
rect 48648 19320 48654 19372
rect 50062 19320 50068 19372
rect 50120 19360 50126 19372
rect 50525 19363 50583 19369
rect 50525 19360 50537 19363
rect 50120 19332 50537 19360
rect 50120 19320 50126 19332
rect 50525 19329 50537 19332
rect 50571 19329 50583 19363
rect 52564 19360 52592 19400
rect 52638 19388 52644 19440
rect 52696 19428 52702 19440
rect 56502 19428 56508 19440
rect 52696 19400 56508 19428
rect 52696 19388 52702 19400
rect 56502 19388 56508 19400
rect 56560 19388 56566 19440
rect 56594 19388 56600 19440
rect 56652 19428 56658 19440
rect 57422 19428 57428 19440
rect 56652 19400 57428 19428
rect 56652 19388 56658 19400
rect 57422 19388 57428 19400
rect 57480 19388 57486 19440
rect 57514 19388 57520 19440
rect 57572 19428 57578 19440
rect 61930 19428 61936 19440
rect 57572 19400 61936 19428
rect 57572 19388 57578 19400
rect 61930 19388 61936 19400
rect 61988 19388 61994 19440
rect 64598 19388 64604 19440
rect 64656 19428 64662 19440
rect 67266 19428 67272 19440
rect 64656 19400 67272 19428
rect 64656 19388 64662 19400
rect 67266 19388 67272 19400
rect 67324 19388 67330 19440
rect 69474 19388 69480 19440
rect 69532 19428 69538 19440
rect 72970 19428 72976 19440
rect 69532 19400 72976 19428
rect 69532 19388 69538 19400
rect 72970 19388 72976 19400
rect 73028 19388 73034 19440
rect 60734 19360 60740 19372
rect 52564 19332 60740 19360
rect 50525 19323 50583 19329
rect 60734 19320 60740 19332
rect 60792 19320 60798 19372
rect 60826 19320 60832 19372
rect 60884 19360 60890 19372
rect 61013 19363 61071 19369
rect 61013 19360 61025 19363
rect 60884 19332 61025 19360
rect 60884 19320 60890 19332
rect 60936 19329 61025 19332
rect 61059 19329 61071 19363
rect 60936 19323 61071 19329
rect 70228 19332 70624 19360
rect 60936 19306 61056 19323
rect 45830 19292 45836 19304
rect 36964 19264 45232 19292
rect 45296 19264 45836 19292
rect 36964 19252 36970 19264
rect 5534 19184 5540 19236
rect 5592 19224 5598 19236
rect 21634 19224 21640 19236
rect 5592 19196 21640 19224
rect 5592 19184 5598 19196
rect 21634 19184 21640 19196
rect 21692 19184 21698 19236
rect 23014 19184 23020 19236
rect 23072 19224 23078 19236
rect 34698 19224 34704 19236
rect 23072 19196 34704 19224
rect 23072 19184 23078 19196
rect 34698 19184 34704 19196
rect 34756 19184 34762 19236
rect 35802 19184 35808 19236
rect 35860 19224 35866 19236
rect 35860 19196 36308 19224
rect 35860 19184 35866 19196
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 22462 19156 22468 19168
rect 10192 19128 22468 19156
rect 10192 19116 10198 19128
rect 22462 19116 22468 19128
rect 22520 19116 22526 19168
rect 22738 19116 22744 19168
rect 22796 19156 22802 19168
rect 30834 19156 30840 19168
rect 22796 19128 30840 19156
rect 22796 19116 22802 19128
rect 30834 19116 30840 19128
rect 30892 19116 30898 19168
rect 36280 19156 36308 19196
rect 36722 19184 36728 19236
rect 36780 19224 36786 19236
rect 43438 19224 43444 19236
rect 36780 19196 43444 19224
rect 36780 19184 36786 19196
rect 43438 19184 43444 19196
rect 43496 19184 43502 19236
rect 36541 19159 36599 19165
rect 36541 19156 36553 19159
rect 36280 19128 36553 19156
rect 36541 19125 36553 19128
rect 36587 19125 36599 19159
rect 36541 19119 36599 19125
rect 36630 19116 36636 19168
rect 36688 19156 36694 19168
rect 44082 19156 44088 19168
rect 36688 19128 44088 19156
rect 36688 19116 36694 19128
rect 44082 19116 44088 19128
rect 44140 19116 44146 19168
rect 44634 19116 44640 19168
rect 44692 19156 44698 19168
rect 44729 19159 44787 19165
rect 44729 19156 44741 19159
rect 44692 19128 44741 19156
rect 44692 19116 44698 19128
rect 44729 19125 44741 19128
rect 44775 19125 44787 19159
rect 45204 19156 45232 19264
rect 45830 19252 45836 19264
rect 45888 19252 45894 19304
rect 46109 19295 46167 19301
rect 46109 19261 46121 19295
rect 46155 19292 46167 19295
rect 46198 19292 46204 19304
rect 46155 19264 46204 19292
rect 46155 19261 46167 19264
rect 46109 19255 46167 19261
rect 46198 19252 46204 19264
rect 46256 19252 46262 19304
rect 46934 19252 46940 19304
rect 46992 19292 46998 19304
rect 47946 19292 47952 19304
rect 46992 19264 47952 19292
rect 46992 19252 46998 19264
rect 47946 19252 47952 19264
rect 48004 19252 48010 19304
rect 50246 19292 50252 19304
rect 50207 19264 50252 19292
rect 50246 19252 50252 19264
rect 50304 19252 50310 19304
rect 50430 19292 50436 19304
rect 50391 19264 50436 19292
rect 50430 19252 50436 19264
rect 50488 19252 50494 19304
rect 50614 19292 50620 19304
rect 50575 19264 50620 19292
rect 50614 19252 50620 19264
rect 50672 19252 50678 19304
rect 50798 19292 50804 19304
rect 50759 19264 50804 19292
rect 50798 19252 50804 19264
rect 50856 19252 50862 19304
rect 52365 19295 52423 19301
rect 52365 19261 52377 19295
rect 52411 19292 52423 19295
rect 58434 19292 58440 19304
rect 52411 19264 58440 19292
rect 52411 19261 52423 19264
rect 52365 19255 52423 19261
rect 58434 19252 58440 19264
rect 58492 19252 58498 19304
rect 58618 19252 58624 19304
rect 58676 19292 58682 19304
rect 60366 19292 60372 19304
rect 58676 19264 60372 19292
rect 58676 19252 58682 19264
rect 60366 19252 60372 19264
rect 60424 19292 60430 19304
rect 60461 19295 60519 19301
rect 60461 19292 60473 19295
rect 60424 19264 60473 19292
rect 60424 19252 60430 19264
rect 60461 19261 60473 19264
rect 60507 19261 60519 19295
rect 60461 19255 60519 19261
rect 51258 19224 51264 19236
rect 50908 19196 51264 19224
rect 50798 19156 50804 19168
rect 45204 19128 50804 19156
rect 44729 19119 44787 19125
rect 50798 19116 50804 19128
rect 50856 19156 50862 19168
rect 50908 19156 50936 19196
rect 51258 19184 51264 19196
rect 51316 19184 51322 19236
rect 52638 19224 52644 19236
rect 52551 19196 52644 19224
rect 52638 19184 52644 19196
rect 52696 19224 52702 19236
rect 60642 19224 60648 19236
rect 52696 19196 60648 19224
rect 52696 19184 52702 19196
rect 60642 19184 60648 19196
rect 60700 19184 60706 19236
rect 50856 19128 50936 19156
rect 50985 19159 51043 19165
rect 50856 19116 50862 19128
rect 50985 19125 50997 19159
rect 51031 19156 51043 19159
rect 51074 19156 51080 19168
rect 51031 19128 51080 19156
rect 51031 19125 51043 19128
rect 50985 19119 51043 19125
rect 51074 19116 51080 19128
rect 51132 19116 51138 19168
rect 51166 19116 51172 19168
rect 51224 19156 51230 19168
rect 54754 19156 54760 19168
rect 51224 19128 54760 19156
rect 51224 19116 51230 19128
rect 54754 19116 54760 19128
rect 54812 19116 54818 19168
rect 55858 19116 55864 19168
rect 55916 19156 55922 19168
rect 60734 19156 60740 19168
rect 55916 19128 60740 19156
rect 55916 19116 55922 19128
rect 60734 19116 60740 19128
rect 60792 19116 60798 19168
rect 60936 19156 60964 19306
rect 61102 19252 61108 19304
rect 61160 19292 61166 19304
rect 70228 19292 70256 19332
rect 61160 19264 70256 19292
rect 70596 19292 70624 19332
rect 71866 19320 71872 19372
rect 71924 19360 71930 19372
rect 72602 19360 72608 19372
rect 71924 19332 72608 19360
rect 71924 19320 71930 19332
rect 72602 19320 72608 19332
rect 72660 19320 72666 19372
rect 98089 19363 98147 19369
rect 98089 19329 98101 19363
rect 98135 19360 98147 19363
rect 98362 19360 98368 19372
rect 98135 19332 98368 19360
rect 98135 19329 98147 19332
rect 98089 19323 98147 19329
rect 98362 19320 98368 19332
rect 98420 19320 98426 19372
rect 73246 19292 73252 19304
rect 70596 19264 73252 19292
rect 61160 19252 61166 19264
rect 73246 19252 73252 19264
rect 73304 19252 73310 19304
rect 63218 19184 63224 19236
rect 63276 19224 63282 19236
rect 63276 19196 70532 19224
rect 63276 19184 63282 19196
rect 69014 19156 69020 19168
rect 60936 19128 69020 19156
rect 69014 19116 69020 19128
rect 69072 19116 69078 19168
rect 70504 19156 70532 19196
rect 75914 19156 75920 19168
rect 70504 19128 75920 19156
rect 75914 19116 75920 19128
rect 75972 19116 75978 19168
rect 1104 19066 98808 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 50326 19066
rect 50378 19014 50390 19066
rect 50442 19014 50454 19066
rect 50506 19014 50518 19066
rect 50570 19014 81046 19066
rect 81098 19014 81110 19066
rect 81162 19014 81174 19066
rect 81226 19014 81238 19066
rect 81290 19014 98808 19066
rect 1104 18992 98808 19014
rect 5626 18912 5632 18964
rect 5684 18952 5690 18964
rect 5684 18924 12434 18952
rect 5684 18912 5690 18924
rect 6822 18844 6828 18896
rect 6880 18884 6886 18896
rect 7009 18887 7067 18893
rect 7009 18884 7021 18887
rect 6880 18856 7021 18884
rect 6880 18844 6886 18856
rect 7009 18853 7021 18856
rect 7055 18884 7067 18887
rect 7193 18887 7251 18893
rect 7193 18884 7205 18887
rect 7055 18856 7205 18884
rect 7055 18853 7067 18856
rect 7009 18847 7067 18853
rect 7193 18853 7205 18856
rect 7239 18853 7251 18887
rect 12406 18884 12434 18924
rect 13538 18912 13544 18964
rect 13596 18952 13602 18964
rect 13596 18924 16528 18952
rect 13596 18912 13602 18924
rect 16500 18884 16528 18924
rect 17310 18912 17316 18964
rect 17368 18952 17374 18964
rect 35802 18952 35808 18964
rect 17368 18924 35808 18952
rect 17368 18912 17374 18924
rect 35802 18912 35808 18924
rect 35860 18912 35866 18964
rect 36722 18912 36728 18964
rect 36780 18952 36786 18964
rect 39022 18952 39028 18964
rect 36780 18924 39028 18952
rect 36780 18912 36786 18924
rect 39022 18912 39028 18924
rect 39080 18912 39086 18964
rect 41064 18924 41276 18952
rect 41064 18884 41092 18924
rect 12406 18856 15700 18884
rect 16500 18856 41092 18884
rect 41248 18884 41276 18924
rect 44542 18912 44548 18964
rect 44600 18952 44606 18964
rect 45462 18952 45468 18964
rect 44600 18924 45468 18952
rect 44600 18912 44606 18924
rect 45462 18912 45468 18924
rect 45520 18912 45526 18964
rect 46290 18912 46296 18964
rect 46348 18952 46354 18964
rect 55858 18952 55864 18964
rect 46348 18924 55864 18952
rect 46348 18912 46354 18924
rect 55858 18912 55864 18924
rect 55916 18912 55922 18964
rect 56410 18912 56416 18964
rect 56468 18952 56474 18964
rect 59354 18952 59360 18964
rect 56468 18924 59360 18952
rect 56468 18912 56474 18924
rect 59354 18912 59360 18924
rect 59412 18912 59418 18964
rect 59446 18912 59452 18964
rect 59504 18952 59510 18964
rect 59541 18955 59599 18961
rect 59541 18952 59553 18955
rect 59504 18924 59553 18952
rect 59504 18912 59510 18924
rect 59541 18921 59553 18924
rect 59587 18921 59599 18955
rect 62114 18952 62120 18964
rect 59541 18915 59599 18921
rect 60016 18924 62120 18952
rect 60016 18884 60044 18924
rect 62114 18912 62120 18924
rect 62172 18912 62178 18964
rect 62390 18912 62396 18964
rect 62448 18952 62454 18964
rect 76098 18952 76104 18964
rect 62448 18924 76104 18952
rect 62448 18912 62454 18924
rect 76098 18912 76104 18924
rect 76156 18912 76162 18964
rect 41248 18856 60044 18884
rect 7193 18847 7251 18853
rect 4985 18819 5043 18825
rect 4985 18785 4997 18819
rect 5031 18816 5043 18819
rect 5169 18819 5227 18825
rect 5169 18816 5181 18819
rect 5031 18788 5181 18816
rect 5031 18785 5043 18788
rect 4985 18779 5043 18785
rect 5169 18785 5181 18788
rect 5215 18816 5227 18819
rect 6641 18819 6699 18825
rect 6641 18816 6653 18819
rect 5215 18788 6653 18816
rect 5215 18785 5227 18788
rect 5169 18779 5227 18785
rect 6641 18785 6653 18788
rect 6687 18816 6699 18819
rect 6840 18816 6868 18844
rect 6687 18788 6868 18816
rect 6917 18819 6975 18825
rect 6687 18785 6699 18788
rect 6641 18779 6699 18785
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 8202 18816 8208 18828
rect 6963 18788 8208 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 8202 18776 8208 18788
rect 8260 18816 8266 18828
rect 15565 18819 15623 18825
rect 15565 18816 15577 18819
rect 8260 18788 15577 18816
rect 8260 18776 8266 18788
rect 15565 18785 15577 18788
rect 15611 18785 15623 18819
rect 15672 18816 15700 18856
rect 60826 18844 60832 18896
rect 60884 18884 60890 18896
rect 63402 18884 63408 18896
rect 60884 18856 63408 18884
rect 60884 18844 60890 18856
rect 63402 18844 63408 18856
rect 63460 18844 63466 18896
rect 63494 18844 63500 18896
rect 63552 18884 63558 18896
rect 69290 18884 69296 18896
rect 63552 18856 69296 18884
rect 63552 18844 63558 18856
rect 69290 18844 69296 18856
rect 69348 18844 69354 18896
rect 71041 18887 71099 18893
rect 71041 18884 71053 18887
rect 70964 18856 71053 18884
rect 70964 18828 70992 18856
rect 71041 18853 71053 18856
rect 71087 18853 71099 18887
rect 71041 18847 71099 18853
rect 72418 18844 72424 18896
rect 72476 18884 72482 18896
rect 82078 18884 82084 18896
rect 72476 18856 82084 18884
rect 72476 18844 72482 18856
rect 82078 18844 82084 18856
rect 82136 18844 82142 18896
rect 33594 18816 33600 18828
rect 15672 18788 33600 18816
rect 15565 18779 15623 18785
rect 33594 18776 33600 18788
rect 33652 18776 33658 18828
rect 33686 18776 33692 18828
rect 33744 18816 33750 18828
rect 35250 18816 35256 18828
rect 33744 18788 35256 18816
rect 33744 18776 33750 18788
rect 35250 18776 35256 18788
rect 35308 18776 35314 18828
rect 35802 18776 35808 18828
rect 35860 18816 35866 18828
rect 35860 18788 36584 18816
rect 35860 18776 35866 18788
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 13872 18720 15853 18748
rect 13872 18708 13878 18720
rect 15841 18717 15853 18720
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 16298 18708 16304 18760
rect 16356 18748 16362 18760
rect 17954 18748 17960 18760
rect 16356 18720 17960 18748
rect 16356 18708 16362 18720
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 22646 18708 22652 18760
rect 22704 18748 22710 18760
rect 25222 18748 25228 18760
rect 22704 18720 25228 18748
rect 22704 18708 22710 18720
rect 25222 18708 25228 18720
rect 25280 18708 25286 18760
rect 25314 18708 25320 18760
rect 25372 18748 25378 18760
rect 25682 18748 25688 18760
rect 25372 18720 25688 18748
rect 25372 18708 25378 18720
rect 25682 18708 25688 18720
rect 25740 18748 25746 18760
rect 26510 18748 26516 18760
rect 25740 18720 26516 18748
rect 25740 18708 25746 18720
rect 26510 18708 26516 18720
rect 26568 18708 26574 18760
rect 26878 18708 26884 18760
rect 26936 18748 26942 18760
rect 36446 18748 36452 18760
rect 26936 18720 36452 18748
rect 26936 18708 26942 18720
rect 36446 18708 36452 18720
rect 36504 18708 36510 18760
rect 36556 18748 36584 18788
rect 36722 18776 36728 18828
rect 36780 18816 36786 18828
rect 36780 18788 41092 18816
rect 36780 18776 36786 18788
rect 40034 18748 40040 18760
rect 36556 18720 40040 18748
rect 40034 18708 40040 18720
rect 40092 18708 40098 18760
rect 41064 18748 41092 18788
rect 41322 18776 41328 18828
rect 41380 18816 41386 18828
rect 47302 18816 47308 18828
rect 41380 18788 47308 18816
rect 41380 18776 41386 18788
rect 47302 18776 47308 18788
rect 47360 18776 47366 18828
rect 50798 18776 50804 18828
rect 50856 18816 50862 18828
rect 53006 18825 53012 18828
rect 52549 18819 52607 18825
rect 52549 18816 52561 18819
rect 50856 18788 52561 18816
rect 50856 18776 50862 18788
rect 52549 18785 52561 18788
rect 52595 18785 52607 18819
rect 52953 18819 53012 18825
rect 52549 18779 52607 18785
rect 52656 18788 52868 18816
rect 52656 18748 52684 18788
rect 52840 18757 52868 18788
rect 52953 18785 52965 18819
rect 52999 18785 53012 18819
rect 52953 18779 53012 18785
rect 53006 18776 53012 18779
rect 53064 18776 53070 18828
rect 53098 18776 53104 18828
rect 53156 18816 53162 18828
rect 53156 18788 53201 18816
rect 53156 18776 53162 18788
rect 56042 18776 56048 18828
rect 56100 18816 56106 18828
rect 59354 18816 59360 18828
rect 56100 18788 59360 18816
rect 56100 18776 56106 18788
rect 59354 18776 59360 18788
rect 59412 18776 59418 18828
rect 59541 18819 59599 18825
rect 59541 18785 59553 18819
rect 59587 18816 59599 18819
rect 59722 18816 59728 18828
rect 59587 18788 59728 18816
rect 59587 18785 59599 18788
rect 59541 18779 59599 18785
rect 59722 18776 59728 18788
rect 59780 18776 59786 18828
rect 59814 18776 59820 18828
rect 59872 18816 59878 18828
rect 69474 18816 69480 18828
rect 59872 18788 69480 18816
rect 59872 18776 59878 18788
rect 69474 18776 69480 18788
rect 69532 18776 69538 18828
rect 69750 18776 69756 18828
rect 69808 18816 69814 18828
rect 70670 18816 70676 18828
rect 69808 18788 70676 18816
rect 69808 18776 69814 18788
rect 70670 18776 70676 18788
rect 70728 18776 70734 18828
rect 70762 18776 70768 18828
rect 70820 18816 70826 18828
rect 70820 18788 70865 18816
rect 70820 18776 70826 18788
rect 70946 18776 70952 18828
rect 71004 18776 71010 18828
rect 71130 18776 71136 18828
rect 71188 18816 71194 18828
rect 72878 18816 72884 18828
rect 71188 18788 72884 18816
rect 71188 18776 71194 18788
rect 72878 18776 72884 18788
rect 72936 18816 72942 18828
rect 78122 18816 78128 18828
rect 72936 18788 78128 18816
rect 72936 18776 72942 18788
rect 78122 18776 78128 18788
rect 78180 18776 78186 18828
rect 78232 18788 78444 18816
rect 41064 18720 52684 18748
rect 52733 18751 52791 18757
rect 52733 18717 52745 18751
rect 52779 18717 52791 18751
rect 52733 18711 52791 18717
rect 52825 18751 52883 18757
rect 52825 18717 52837 18751
rect 52871 18748 52883 18751
rect 78232 18748 78260 18788
rect 52871 18720 78260 18748
rect 78416 18748 78444 18788
rect 92474 18748 92480 18760
rect 78416 18720 92480 18748
rect 52871 18717 52883 18720
rect 52825 18711 52883 18717
rect 1946 18640 1952 18692
rect 2004 18680 2010 18692
rect 8570 18680 8576 18692
rect 2004 18652 6040 18680
rect 2004 18640 2010 18652
rect 5258 18572 5264 18624
rect 5316 18612 5322 18624
rect 5353 18615 5411 18621
rect 5353 18612 5365 18615
rect 5316 18584 5365 18612
rect 5316 18572 5322 18584
rect 5353 18581 5365 18584
rect 5399 18581 5411 18615
rect 6012 18612 6040 18652
rect 6932 18652 8576 18680
rect 6932 18612 6960 18652
rect 8570 18640 8576 18652
rect 8628 18640 8634 18692
rect 17218 18640 17224 18692
rect 17276 18680 17282 18692
rect 40954 18680 40960 18692
rect 17276 18652 40960 18680
rect 17276 18640 17282 18652
rect 40954 18640 40960 18652
rect 41012 18640 41018 18692
rect 52365 18683 52423 18689
rect 52365 18680 52377 18683
rect 46308 18652 52377 18680
rect 16942 18612 16948 18624
rect 6012 18584 6960 18612
rect 16903 18584 16948 18612
rect 5353 18575 5411 18581
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 46308 18612 46336 18652
rect 52365 18649 52377 18652
rect 52411 18649 52423 18683
rect 52365 18643 52423 18649
rect 52748 18680 52776 18711
rect 92474 18708 92480 18720
rect 92532 18708 92538 18760
rect 60826 18680 60832 18692
rect 52748 18652 60832 18680
rect 17184 18584 46336 18612
rect 17184 18572 17190 18584
rect 47118 18572 47124 18624
rect 47176 18612 47182 18624
rect 51718 18612 51724 18624
rect 47176 18584 51724 18612
rect 47176 18572 47182 18584
rect 51718 18572 51724 18584
rect 51776 18572 51782 18624
rect 52270 18612 52276 18624
rect 52183 18584 52276 18612
rect 52270 18572 52276 18584
rect 52328 18612 52334 18624
rect 52748 18612 52776 18652
rect 60826 18640 60832 18652
rect 60884 18640 60890 18692
rect 60918 18640 60924 18692
rect 60976 18680 60982 18692
rect 64506 18680 64512 18692
rect 60976 18652 64512 18680
rect 60976 18640 60982 18652
rect 64506 18640 64512 18652
rect 64564 18640 64570 18692
rect 65518 18640 65524 18692
rect 65576 18680 65582 18692
rect 78214 18680 78220 18692
rect 65576 18652 78220 18680
rect 65576 18640 65582 18652
rect 78214 18640 78220 18652
rect 78272 18640 78278 18692
rect 78306 18640 78312 18692
rect 78364 18680 78370 18692
rect 82722 18680 82728 18692
rect 78364 18652 82728 18680
rect 78364 18640 78370 18652
rect 82722 18640 82728 18652
rect 82780 18640 82786 18692
rect 52328 18584 52776 18612
rect 52328 18572 52334 18584
rect 54846 18572 54852 18624
rect 54904 18612 54910 18624
rect 59814 18612 59820 18624
rect 54904 18584 59820 18612
rect 54904 18572 54910 18584
rect 59814 18572 59820 18584
rect 59872 18572 59878 18624
rect 61930 18572 61936 18624
rect 61988 18612 61994 18624
rect 74629 18615 74687 18621
rect 74629 18612 74641 18615
rect 61988 18584 74641 18612
rect 61988 18572 61994 18584
rect 74629 18581 74641 18584
rect 74675 18581 74687 18615
rect 74629 18575 74687 18581
rect 76282 18572 76288 18624
rect 76340 18612 76346 18624
rect 93946 18612 93952 18624
rect 76340 18584 93952 18612
rect 76340 18572 76346 18584
rect 93946 18572 93952 18584
rect 94004 18572 94010 18624
rect 1104 18522 98808 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 65686 18522
rect 65738 18470 65750 18522
rect 65802 18470 65814 18522
rect 65866 18470 65878 18522
rect 65930 18470 96406 18522
rect 96458 18470 96470 18522
rect 96522 18470 96534 18522
rect 96586 18470 96598 18522
rect 96650 18470 98808 18522
rect 1104 18448 98808 18470
rect 3145 18411 3203 18417
rect 3145 18377 3157 18411
rect 3191 18408 3203 18411
rect 3329 18411 3387 18417
rect 3329 18408 3341 18411
rect 3191 18380 3341 18408
rect 3191 18377 3203 18380
rect 3145 18371 3203 18377
rect 3329 18377 3341 18380
rect 3375 18408 3387 18411
rect 3513 18411 3571 18417
rect 3513 18408 3525 18411
rect 3375 18380 3525 18408
rect 3375 18377 3387 18380
rect 3329 18371 3387 18377
rect 3513 18377 3525 18380
rect 3559 18408 3571 18411
rect 3789 18411 3847 18417
rect 3789 18408 3801 18411
rect 3559 18380 3801 18408
rect 3559 18377 3571 18380
rect 3513 18371 3571 18377
rect 3789 18377 3801 18380
rect 3835 18408 3847 18411
rect 5169 18411 5227 18417
rect 5169 18408 5181 18411
rect 3835 18380 5181 18408
rect 3835 18377 3847 18380
rect 3789 18371 3847 18377
rect 5169 18377 5181 18380
rect 5215 18408 5227 18411
rect 5353 18411 5411 18417
rect 5353 18408 5365 18411
rect 5215 18380 5365 18408
rect 5215 18377 5227 18380
rect 5169 18371 5227 18377
rect 5353 18377 5365 18380
rect 5399 18408 5411 18411
rect 5534 18408 5540 18420
rect 5399 18380 5540 18408
rect 5399 18377 5411 18380
rect 5353 18371 5411 18377
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 12158 18368 12164 18420
rect 12216 18408 12222 18420
rect 17218 18408 17224 18420
rect 12216 18380 17224 18408
rect 12216 18368 12222 18380
rect 17218 18368 17224 18380
rect 17276 18368 17282 18420
rect 22094 18368 22100 18420
rect 22152 18408 22158 18420
rect 33594 18408 33600 18420
rect 22152 18380 33600 18408
rect 22152 18368 22158 18380
rect 33594 18368 33600 18380
rect 33652 18368 33658 18420
rect 35342 18408 35348 18420
rect 33796 18380 35348 18408
rect 6086 18340 6092 18352
rect 4264 18312 6092 18340
rect 4264 18213 4292 18312
rect 6086 18300 6092 18312
rect 6144 18300 6150 18352
rect 7926 18300 7932 18352
rect 7984 18340 7990 18352
rect 7984 18312 10180 18340
rect 7984 18300 7990 18312
rect 4341 18275 4399 18281
rect 4341 18241 4353 18275
rect 4387 18272 4399 18275
rect 4387 18244 8248 18272
rect 4387 18241 4399 18244
rect 4341 18235 4399 18241
rect 4249 18207 4307 18213
rect 4249 18173 4261 18207
rect 4295 18173 4307 18207
rect 4249 18167 4307 18173
rect 4617 18207 4675 18213
rect 4617 18173 4629 18207
rect 4663 18173 4675 18207
rect 4617 18167 4675 18173
rect 4801 18207 4859 18213
rect 4801 18173 4813 18207
rect 4847 18173 4859 18207
rect 4982 18204 4988 18216
rect 4943 18176 4988 18204
rect 4801 18167 4859 18173
rect 4632 18068 4660 18167
rect 4816 18136 4844 18167
rect 4982 18164 4988 18176
rect 5040 18164 5046 18216
rect 8220 18204 8248 18244
rect 8294 18232 8300 18284
rect 8352 18272 8358 18284
rect 9306 18272 9312 18284
rect 8352 18244 9312 18272
rect 8352 18232 8358 18244
rect 9306 18232 9312 18244
rect 9364 18232 9370 18284
rect 10152 18272 10180 18312
rect 10502 18300 10508 18352
rect 10560 18340 10566 18352
rect 26234 18340 26240 18352
rect 10560 18312 26240 18340
rect 10560 18300 10566 18312
rect 26234 18300 26240 18312
rect 26292 18300 26298 18352
rect 26510 18300 26516 18352
rect 26568 18340 26574 18352
rect 33686 18340 33692 18352
rect 26568 18312 33692 18340
rect 26568 18300 26574 18312
rect 33686 18300 33692 18312
rect 33744 18300 33750 18352
rect 17126 18272 17132 18284
rect 10152 18244 17132 18272
rect 17126 18232 17132 18244
rect 17184 18232 17190 18284
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 33502 18272 33508 18284
rect 18012 18244 33508 18272
rect 18012 18232 18018 18244
rect 33502 18232 33508 18244
rect 33560 18232 33566 18284
rect 33796 18272 33824 18380
rect 35342 18368 35348 18380
rect 35400 18368 35406 18420
rect 35894 18368 35900 18420
rect 35952 18408 35958 18420
rect 38286 18408 38292 18420
rect 35952 18380 38292 18408
rect 35952 18368 35958 18380
rect 38286 18368 38292 18380
rect 38344 18368 38350 18420
rect 39850 18368 39856 18420
rect 39908 18408 39914 18420
rect 50706 18408 50712 18420
rect 39908 18380 50712 18408
rect 39908 18368 39914 18380
rect 50706 18368 50712 18380
rect 50764 18368 50770 18420
rect 56502 18368 56508 18420
rect 56560 18408 56566 18420
rect 65518 18408 65524 18420
rect 56560 18380 65524 18408
rect 56560 18368 56566 18380
rect 65518 18368 65524 18380
rect 65576 18368 65582 18420
rect 66254 18368 66260 18420
rect 66312 18408 66318 18420
rect 66312 18380 70808 18408
rect 66312 18368 66318 18380
rect 35161 18343 35219 18349
rect 35161 18309 35173 18343
rect 35207 18340 35219 18343
rect 35250 18340 35256 18352
rect 35207 18312 35256 18340
rect 35207 18309 35219 18312
rect 35161 18303 35219 18309
rect 35250 18300 35256 18312
rect 35308 18300 35314 18352
rect 35802 18300 35808 18352
rect 35860 18340 35866 18352
rect 36078 18340 36084 18352
rect 35860 18312 36084 18340
rect 35860 18300 35866 18312
rect 36078 18300 36084 18312
rect 36136 18300 36142 18352
rect 36446 18300 36452 18352
rect 36504 18340 36510 18352
rect 41414 18340 41420 18352
rect 36504 18312 41420 18340
rect 36504 18300 36510 18312
rect 41414 18300 41420 18312
rect 41472 18300 41478 18352
rect 43438 18300 43444 18352
rect 43496 18340 43502 18352
rect 50614 18340 50620 18352
rect 43496 18312 50620 18340
rect 43496 18300 43502 18312
rect 50614 18300 50620 18312
rect 50672 18300 50678 18352
rect 51258 18300 51264 18352
rect 51316 18340 51322 18352
rect 63586 18340 63592 18352
rect 51316 18312 63592 18340
rect 51316 18300 51322 18312
rect 63586 18300 63592 18312
rect 63644 18300 63650 18352
rect 63678 18300 63684 18352
rect 63736 18340 63742 18352
rect 65610 18340 65616 18352
rect 63736 18312 65616 18340
rect 63736 18300 63742 18312
rect 65610 18300 65616 18312
rect 65668 18300 65674 18352
rect 65794 18300 65800 18352
rect 65852 18340 65858 18352
rect 67818 18340 67824 18352
rect 65852 18312 67824 18340
rect 65852 18300 65858 18312
rect 67818 18300 67824 18312
rect 67876 18340 67882 18352
rect 69750 18340 69756 18352
rect 67876 18312 69756 18340
rect 67876 18300 67882 18312
rect 69750 18300 69756 18312
rect 69808 18300 69814 18352
rect 70780 18340 70808 18380
rect 70854 18368 70860 18420
rect 70912 18408 70918 18420
rect 92658 18408 92664 18420
rect 70912 18380 92664 18408
rect 70912 18368 70918 18380
rect 92658 18368 92664 18380
rect 92716 18368 92722 18420
rect 72973 18343 73031 18349
rect 72973 18340 72985 18343
rect 70780 18312 72985 18340
rect 72973 18309 72985 18312
rect 73019 18309 73031 18343
rect 72973 18303 73031 18309
rect 73154 18300 73160 18352
rect 73212 18349 73218 18352
rect 73212 18343 73261 18349
rect 73212 18309 73215 18343
rect 73249 18309 73261 18343
rect 73338 18340 73344 18352
rect 73299 18312 73344 18340
rect 73212 18303 73261 18309
rect 73212 18300 73218 18303
rect 73338 18300 73344 18312
rect 73396 18300 73402 18352
rect 34057 18275 34115 18281
rect 34057 18272 34069 18275
rect 33796 18244 34069 18272
rect 34057 18241 34069 18244
rect 34103 18241 34115 18275
rect 34057 18235 34115 18241
rect 34146 18232 34152 18284
rect 34204 18272 34210 18284
rect 39584 18275 39642 18281
rect 34204 18244 39527 18272
rect 34204 18232 34210 18244
rect 26878 18204 26884 18216
rect 8220 18176 26884 18204
rect 26878 18164 26884 18176
rect 26936 18164 26942 18216
rect 30374 18164 30380 18216
rect 30432 18204 30438 18216
rect 33781 18207 33839 18213
rect 33781 18204 33793 18207
rect 30432 18176 33793 18204
rect 30432 18164 30438 18176
rect 33781 18173 33793 18176
rect 33827 18173 33839 18207
rect 33781 18167 33839 18173
rect 34422 18164 34428 18216
rect 34480 18204 34486 18216
rect 36906 18204 36912 18216
rect 34480 18176 36912 18204
rect 34480 18164 34486 18176
rect 36906 18164 36912 18176
rect 36964 18164 36970 18216
rect 37274 18164 37280 18216
rect 37332 18204 37338 18216
rect 38102 18204 38108 18216
rect 37332 18176 38108 18204
rect 37332 18164 37338 18176
rect 38102 18164 38108 18176
rect 38160 18204 38166 18216
rect 38562 18204 38568 18216
rect 38160 18176 38568 18204
rect 38160 18164 38166 18176
rect 38562 18164 38568 18176
rect 38620 18164 38626 18216
rect 39298 18204 39304 18216
rect 39259 18176 39304 18204
rect 39298 18164 39304 18176
rect 39356 18164 39362 18216
rect 39499 18213 39527 18244
rect 39584 18241 39596 18275
rect 39630 18272 39642 18275
rect 39758 18272 39764 18284
rect 39630 18244 39764 18272
rect 39630 18241 39642 18244
rect 39584 18235 39642 18241
rect 39758 18232 39764 18244
rect 39816 18232 39822 18284
rect 41782 18232 41788 18284
rect 41840 18272 41846 18284
rect 56042 18272 56048 18284
rect 41840 18244 56048 18272
rect 41840 18232 41846 18244
rect 56042 18232 56048 18244
rect 56100 18232 56106 18284
rect 56134 18232 56140 18284
rect 56192 18272 56198 18284
rect 62390 18272 62396 18284
rect 56192 18244 62396 18272
rect 56192 18232 56198 18244
rect 62390 18232 62396 18244
rect 62448 18232 62454 18284
rect 62574 18232 62580 18284
rect 62632 18272 62638 18284
rect 65518 18272 65524 18284
rect 62632 18244 65524 18272
rect 62632 18232 62638 18244
rect 65518 18232 65524 18244
rect 65576 18232 65582 18284
rect 65812 18244 70164 18272
rect 39484 18207 39542 18213
rect 39484 18173 39496 18207
rect 39530 18173 39542 18207
rect 39484 18167 39542 18173
rect 39669 18207 39727 18213
rect 39669 18173 39681 18207
rect 39715 18173 39727 18207
rect 39669 18167 39727 18173
rect 39853 18207 39911 18213
rect 39853 18173 39865 18207
rect 39899 18204 39911 18207
rect 43622 18204 43628 18216
rect 39899 18176 43628 18204
rect 39899 18173 39911 18176
rect 39853 18167 39911 18173
rect 4816 18108 8524 18136
rect 8294 18068 8300 18080
rect 4632 18040 8300 18068
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 8496 18068 8524 18108
rect 8570 18096 8576 18148
rect 8628 18136 8634 18148
rect 8628 18108 22094 18136
rect 8628 18096 8634 18108
rect 13354 18068 13360 18080
rect 8496 18040 13360 18068
rect 13354 18028 13360 18040
rect 13412 18068 13418 18080
rect 13538 18068 13544 18080
rect 13412 18040 13544 18068
rect 13412 18028 13418 18040
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 22066 18068 22094 18108
rect 22922 18096 22928 18148
rect 22980 18136 22986 18148
rect 31110 18136 31116 18148
rect 22980 18108 31116 18136
rect 22980 18096 22986 18108
rect 31110 18096 31116 18108
rect 31168 18096 31174 18148
rect 31478 18096 31484 18148
rect 31536 18136 31542 18148
rect 32490 18136 32496 18148
rect 31536 18108 32496 18136
rect 31536 18096 31542 18108
rect 32490 18096 32496 18108
rect 32548 18096 32554 18148
rect 33042 18096 33048 18148
rect 33100 18136 33106 18148
rect 39117 18139 39175 18145
rect 39117 18136 39129 18139
rect 33100 18108 33548 18136
rect 33100 18096 33106 18108
rect 33410 18068 33416 18080
rect 22066 18040 33416 18068
rect 33410 18028 33416 18040
rect 33468 18028 33474 18080
rect 33520 18068 33548 18108
rect 34716 18108 39129 18136
rect 34716 18068 34744 18108
rect 39117 18105 39129 18108
rect 39163 18136 39175 18139
rect 39684 18136 39712 18167
rect 43622 18164 43628 18176
rect 43680 18164 43686 18216
rect 45830 18164 45836 18216
rect 45888 18204 45894 18216
rect 46014 18204 46020 18216
rect 45888 18176 46020 18204
rect 45888 18164 45894 18176
rect 46014 18164 46020 18176
rect 46072 18164 46078 18216
rect 46106 18164 46112 18216
rect 46164 18204 46170 18216
rect 56410 18204 56416 18216
rect 46164 18176 56416 18204
rect 46164 18164 46170 18176
rect 56410 18164 56416 18176
rect 56468 18164 56474 18216
rect 59354 18164 59360 18216
rect 59412 18204 59418 18216
rect 60550 18204 60556 18216
rect 59412 18176 60556 18204
rect 59412 18164 59418 18176
rect 60550 18164 60556 18176
rect 60608 18164 60614 18216
rect 62666 18204 62672 18216
rect 62579 18176 62672 18204
rect 62666 18164 62672 18176
rect 62724 18204 62730 18216
rect 65812 18204 65840 18244
rect 69750 18204 69756 18216
rect 62724 18176 65840 18204
rect 69711 18176 69756 18204
rect 62724 18164 62730 18176
rect 69750 18164 69756 18176
rect 69808 18164 69814 18216
rect 70026 18204 70032 18216
rect 69987 18176 70032 18204
rect 70026 18164 70032 18176
rect 70084 18164 70090 18216
rect 70136 18204 70164 18244
rect 70210 18232 70216 18284
rect 70268 18272 70274 18284
rect 73433 18275 73491 18281
rect 73433 18272 73445 18275
rect 70268 18244 73445 18272
rect 70268 18232 70274 18244
rect 73433 18241 73445 18244
rect 73479 18241 73491 18275
rect 73706 18272 73712 18284
rect 73667 18244 73712 18272
rect 73433 18235 73491 18241
rect 73706 18232 73712 18244
rect 73764 18232 73770 18284
rect 89530 18272 89536 18284
rect 89491 18244 89536 18272
rect 89530 18232 89536 18244
rect 89588 18232 89594 18284
rect 92474 18232 92480 18284
rect 92532 18272 92538 18284
rect 92934 18272 92940 18284
rect 92532 18244 92940 18272
rect 92532 18232 92538 18244
rect 92934 18232 92940 18244
rect 92992 18232 92998 18284
rect 70762 18204 70768 18216
rect 70136 18176 70768 18204
rect 70762 18164 70768 18176
rect 70820 18164 70826 18216
rect 72973 18207 73031 18213
rect 72973 18173 72985 18207
rect 73019 18204 73031 18207
rect 75917 18207 75975 18213
rect 73019 18176 73660 18204
rect 73019 18173 73031 18176
rect 72973 18167 73031 18173
rect 63218 18136 63224 18148
rect 39163 18108 60688 18136
rect 63179 18108 63224 18136
rect 39163 18105 39175 18108
rect 39117 18099 39175 18105
rect 33520 18040 34744 18068
rect 35158 18028 35164 18080
rect 35216 18068 35222 18080
rect 39206 18068 39212 18080
rect 35216 18040 39212 18068
rect 35216 18028 35222 18040
rect 39206 18028 39212 18040
rect 39264 18028 39270 18080
rect 39945 18071 40003 18077
rect 39945 18037 39957 18071
rect 39991 18068 40003 18071
rect 41230 18068 41236 18080
rect 39991 18040 41236 18068
rect 39991 18037 40003 18040
rect 39945 18031 40003 18037
rect 41230 18028 41236 18040
rect 41288 18028 41294 18080
rect 41414 18028 41420 18080
rect 41472 18068 41478 18080
rect 60458 18068 60464 18080
rect 41472 18040 60464 18068
rect 41472 18028 41478 18040
rect 60458 18028 60464 18040
rect 60516 18028 60522 18080
rect 60660 18068 60688 18108
rect 63218 18096 63224 18108
rect 63276 18096 63282 18148
rect 71409 18139 71467 18145
rect 71409 18105 71421 18139
rect 71455 18136 71467 18139
rect 71774 18136 71780 18148
rect 71455 18108 71780 18136
rect 71455 18105 71467 18108
rect 71409 18099 71467 18105
rect 71774 18096 71780 18108
rect 71832 18136 71838 18148
rect 72418 18136 72424 18148
rect 71832 18108 72424 18136
rect 71832 18096 71838 18108
rect 72418 18096 72424 18108
rect 72476 18096 72482 18148
rect 73062 18136 73068 18148
rect 73023 18108 73068 18136
rect 73062 18096 73068 18108
rect 73120 18096 73126 18148
rect 73632 18136 73660 18176
rect 75917 18173 75929 18207
rect 75963 18204 75975 18207
rect 77570 18204 77576 18216
rect 75963 18176 77576 18204
rect 75963 18173 75975 18176
rect 75917 18167 75975 18173
rect 77570 18164 77576 18176
rect 77628 18164 77634 18216
rect 82722 18164 82728 18216
rect 82780 18204 82786 18216
rect 89257 18207 89315 18213
rect 89257 18204 89269 18207
rect 82780 18176 89269 18204
rect 82780 18164 82786 18176
rect 89257 18173 89269 18176
rect 89303 18173 89315 18207
rect 92661 18207 92719 18213
rect 92661 18204 92673 18207
rect 89257 18167 89315 18173
rect 91664 18176 92673 18204
rect 91281 18139 91339 18145
rect 91281 18136 91293 18139
rect 73632 18108 80054 18136
rect 78398 18068 78404 18080
rect 60660 18040 78404 18068
rect 78398 18028 78404 18040
rect 78456 18028 78462 18080
rect 80026 18068 80054 18108
rect 89686 18108 91293 18136
rect 89686 18068 89714 18108
rect 91281 18105 91293 18108
rect 91327 18105 91339 18139
rect 91281 18099 91339 18105
rect 91186 18068 91192 18080
rect 80026 18040 89714 18068
rect 91147 18040 91192 18068
rect 91186 18028 91192 18040
rect 91244 18068 91250 18080
rect 91664 18068 91692 18176
rect 92661 18173 92673 18176
rect 92707 18173 92719 18207
rect 92661 18167 92719 18173
rect 91244 18040 91692 18068
rect 91244 18028 91250 18040
rect 1104 17978 98808 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 50326 17978
rect 50378 17926 50390 17978
rect 50442 17926 50454 17978
rect 50506 17926 50518 17978
rect 50570 17926 81046 17978
rect 81098 17926 81110 17978
rect 81162 17926 81174 17978
rect 81226 17926 81238 17978
rect 81290 17926 98808 17978
rect 1104 17904 98808 17926
rect 16298 17824 16304 17876
rect 16356 17864 16362 17876
rect 19334 17864 19340 17876
rect 16356 17836 19340 17864
rect 16356 17824 16362 17836
rect 19334 17824 19340 17836
rect 19392 17864 19398 17876
rect 19392 17836 59676 17864
rect 19392 17824 19398 17836
rect 23014 17756 23020 17808
rect 23072 17796 23078 17808
rect 40126 17796 40132 17808
rect 23072 17768 40132 17796
rect 23072 17756 23078 17768
rect 40126 17756 40132 17768
rect 40184 17756 40190 17808
rect 42794 17756 42800 17808
rect 42852 17796 42858 17808
rect 43806 17796 43812 17808
rect 42852 17768 43812 17796
rect 42852 17756 42858 17768
rect 43806 17756 43812 17768
rect 43864 17796 43870 17808
rect 45462 17796 45468 17808
rect 43864 17768 45468 17796
rect 43864 17756 43870 17768
rect 45462 17756 45468 17768
rect 45520 17756 45526 17808
rect 45554 17756 45560 17808
rect 45612 17796 45618 17808
rect 46290 17796 46296 17808
rect 45612 17768 46296 17796
rect 45612 17756 45618 17768
rect 46290 17756 46296 17768
rect 46348 17756 46354 17808
rect 46382 17756 46388 17808
rect 46440 17796 46446 17808
rect 49142 17796 49148 17808
rect 46440 17768 49148 17796
rect 46440 17756 46446 17768
rect 49142 17756 49148 17768
rect 49200 17756 49206 17808
rect 2501 17731 2559 17737
rect 2501 17697 2513 17731
rect 2547 17728 2559 17731
rect 2590 17728 2596 17740
rect 2547 17700 2596 17728
rect 2547 17697 2559 17700
rect 2501 17691 2559 17697
rect 2590 17688 2596 17700
rect 2648 17688 2654 17740
rect 2869 17731 2927 17737
rect 2869 17697 2881 17731
rect 2915 17728 2927 17731
rect 2958 17728 2964 17740
rect 2915 17700 2964 17728
rect 2915 17697 2927 17700
rect 2869 17691 2927 17697
rect 2958 17688 2964 17700
rect 3016 17688 3022 17740
rect 3053 17731 3111 17737
rect 3053 17697 3065 17731
rect 3099 17697 3111 17731
rect 3053 17691 3111 17697
rect 2130 17660 2136 17672
rect 2091 17632 2136 17660
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 2406 17660 2412 17672
rect 2367 17632 2412 17660
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 3068 17660 3096 17691
rect 20346 17688 20352 17740
rect 20404 17728 20410 17740
rect 20404 17700 21956 17728
rect 20404 17688 20410 17700
rect 21818 17660 21824 17672
rect 3068 17632 21824 17660
rect 21818 17620 21824 17632
rect 21876 17620 21882 17672
rect 21928 17660 21956 17700
rect 22646 17688 22652 17740
rect 22704 17728 22710 17740
rect 26878 17728 26884 17740
rect 22704 17700 26884 17728
rect 22704 17688 22710 17700
rect 26878 17688 26884 17700
rect 26936 17688 26942 17740
rect 53650 17728 53656 17740
rect 27172 17700 53656 17728
rect 27172 17660 27200 17700
rect 53650 17688 53656 17700
rect 53708 17688 53714 17740
rect 55876 17700 59584 17728
rect 28350 17660 28356 17672
rect 21928 17632 27200 17660
rect 28311 17632 28356 17660
rect 28350 17620 28356 17632
rect 28408 17620 28414 17672
rect 28626 17620 28632 17672
rect 28684 17660 28690 17672
rect 30466 17660 30472 17672
rect 28684 17632 30472 17660
rect 28684 17620 28690 17632
rect 30466 17620 30472 17632
rect 30524 17620 30530 17672
rect 31754 17620 31760 17672
rect 31812 17660 31818 17672
rect 40770 17660 40776 17672
rect 31812 17632 40776 17660
rect 31812 17620 31818 17632
rect 40770 17620 40776 17632
rect 40828 17620 40834 17672
rect 40954 17620 40960 17672
rect 41012 17660 41018 17672
rect 46566 17660 46572 17672
rect 41012 17632 46572 17660
rect 41012 17620 41018 17632
rect 46566 17620 46572 17632
rect 46624 17620 46630 17672
rect 48406 17620 48412 17672
rect 48464 17660 48470 17672
rect 55876 17660 55904 17700
rect 59173 17663 59231 17669
rect 59173 17660 59185 17663
rect 48464 17632 55904 17660
rect 57992 17632 59185 17660
rect 48464 17620 48470 17632
rect 1118 17552 1124 17604
rect 1176 17592 1182 17604
rect 48774 17592 48780 17604
rect 1176 17564 48780 17592
rect 1176 17552 1182 17564
rect 48774 17552 48780 17564
rect 48832 17552 48838 17604
rect 49142 17552 49148 17604
rect 49200 17592 49206 17604
rect 57885 17595 57943 17601
rect 57885 17592 57897 17595
rect 49200 17564 57897 17592
rect 49200 17552 49206 17564
rect 57885 17561 57897 17564
rect 57931 17561 57943 17595
rect 57885 17555 57943 17561
rect 6638 17484 6644 17536
rect 6696 17524 6702 17536
rect 31754 17524 31760 17536
rect 6696 17496 31760 17524
rect 6696 17484 6702 17496
rect 31754 17484 31760 17496
rect 31812 17484 31818 17536
rect 31938 17484 31944 17536
rect 31996 17524 32002 17536
rect 42610 17524 42616 17536
rect 31996 17496 42616 17524
rect 31996 17484 32002 17496
rect 42610 17484 42616 17496
rect 42668 17484 42674 17536
rect 43622 17484 43628 17536
rect 43680 17524 43686 17536
rect 56410 17524 56416 17536
rect 43680 17496 56416 17524
rect 43680 17484 43686 17496
rect 56410 17484 56416 17496
rect 56468 17484 56474 17536
rect 56594 17484 56600 17536
rect 56652 17524 56658 17536
rect 57609 17527 57667 17533
rect 57609 17524 57621 17527
rect 56652 17496 57621 17524
rect 56652 17484 56658 17496
rect 57609 17493 57621 17496
rect 57655 17524 57667 17527
rect 57992 17524 58020 17632
rect 59173 17629 59185 17632
rect 59219 17629 59231 17663
rect 59173 17623 59231 17629
rect 59449 17663 59507 17669
rect 59449 17629 59461 17663
rect 59495 17629 59507 17663
rect 59449 17623 59507 17629
rect 57655 17496 58020 17524
rect 59464 17524 59492 17623
rect 59556 17592 59584 17700
rect 59648 17660 59676 17836
rect 59722 17688 59728 17740
rect 59780 17728 59786 17740
rect 61381 17731 61439 17737
rect 61381 17728 61393 17731
rect 59780 17700 61393 17728
rect 59780 17688 59786 17700
rect 61381 17697 61393 17700
rect 61427 17697 61439 17731
rect 61381 17691 61439 17697
rect 64782 17688 64788 17740
rect 64840 17728 64846 17740
rect 72142 17728 72148 17740
rect 64840 17700 72148 17728
rect 64840 17688 64846 17700
rect 72142 17688 72148 17700
rect 72200 17688 72206 17740
rect 64966 17660 64972 17672
rect 59648 17632 64972 17660
rect 64966 17620 64972 17632
rect 65024 17660 65030 17672
rect 66254 17660 66260 17672
rect 65024 17632 66260 17660
rect 65024 17620 65030 17632
rect 66254 17620 66260 17632
rect 66312 17620 66318 17672
rect 74258 17660 74264 17672
rect 70366 17632 74264 17660
rect 70366 17592 70394 17632
rect 74258 17620 74264 17632
rect 74316 17660 74322 17672
rect 78766 17660 78772 17672
rect 74316 17632 78772 17660
rect 74316 17620 74322 17632
rect 78766 17620 78772 17632
rect 78824 17620 78830 17672
rect 59556 17564 70394 17592
rect 75178 17552 75184 17604
rect 75236 17592 75242 17604
rect 83090 17592 83096 17604
rect 75236 17564 83096 17592
rect 75236 17552 75242 17564
rect 83090 17552 83096 17564
rect 83148 17592 83154 17604
rect 83642 17592 83648 17604
rect 83148 17564 83648 17592
rect 83148 17552 83154 17564
rect 83642 17552 83648 17564
rect 83700 17552 83706 17604
rect 61286 17524 61292 17536
rect 59464 17496 61292 17524
rect 57655 17493 57667 17496
rect 57609 17487 57667 17493
rect 61286 17484 61292 17496
rect 61344 17484 61350 17536
rect 61381 17527 61439 17533
rect 61381 17493 61393 17527
rect 61427 17524 61439 17527
rect 90726 17524 90732 17536
rect 61427 17496 90732 17524
rect 61427 17493 61439 17496
rect 61381 17487 61439 17493
rect 90726 17484 90732 17496
rect 90784 17524 90790 17536
rect 94314 17524 94320 17536
rect 90784 17496 94320 17524
rect 90784 17484 90790 17496
rect 94314 17484 94320 17496
rect 94372 17484 94378 17536
rect 1104 17434 98808 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 65686 17434
rect 65738 17382 65750 17434
rect 65802 17382 65814 17434
rect 65866 17382 65878 17434
rect 65930 17382 96406 17434
rect 96458 17382 96470 17434
rect 96522 17382 96534 17434
rect 96586 17382 96598 17434
rect 96650 17382 98808 17434
rect 1104 17360 98808 17382
rect 2038 17280 2044 17332
rect 2096 17320 2102 17332
rect 2314 17320 2320 17332
rect 2096 17292 2320 17320
rect 2096 17280 2102 17292
rect 2314 17280 2320 17292
rect 2372 17280 2378 17332
rect 8018 17280 8024 17332
rect 8076 17320 8082 17332
rect 28902 17320 28908 17332
rect 8076 17292 28908 17320
rect 8076 17280 8082 17292
rect 28902 17280 28908 17292
rect 28960 17280 28966 17332
rect 36354 17320 36360 17332
rect 29012 17292 36360 17320
rect 23290 17252 23296 17264
rect 2746 17224 23296 17252
rect 2406 17144 2412 17196
rect 2464 17184 2470 17196
rect 2746 17184 2774 17224
rect 23290 17212 23296 17224
rect 23348 17252 23354 17264
rect 25590 17252 25596 17264
rect 23348 17224 25596 17252
rect 23348 17212 23354 17224
rect 25590 17212 25596 17224
rect 25648 17212 25654 17264
rect 25682 17212 25688 17264
rect 25740 17252 25746 17264
rect 29012 17252 29040 17292
rect 25740 17224 29040 17252
rect 25740 17212 25746 17224
rect 29086 17212 29092 17264
rect 29144 17252 29150 17264
rect 33962 17252 33968 17264
rect 29144 17224 33968 17252
rect 29144 17212 29150 17224
rect 33962 17212 33968 17224
rect 34020 17212 34026 17264
rect 2464 17156 2774 17184
rect 2464 17144 2470 17156
rect 17034 17144 17040 17196
rect 17092 17184 17098 17196
rect 22646 17184 22652 17196
rect 17092 17156 22652 17184
rect 17092 17144 17098 17156
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 31938 17184 31944 17196
rect 22756 17156 31944 17184
rect 13541 17119 13599 17125
rect 13541 17085 13553 17119
rect 13587 17116 13599 17119
rect 13817 17119 13875 17125
rect 13817 17116 13829 17119
rect 13587 17088 13829 17116
rect 13587 17085 13599 17088
rect 13541 17079 13599 17085
rect 13817 17085 13829 17088
rect 13863 17116 13875 17119
rect 22756 17116 22784 17156
rect 31938 17144 31944 17156
rect 31996 17144 32002 17196
rect 32030 17144 32036 17196
rect 32088 17184 32094 17196
rect 34517 17187 34575 17193
rect 34517 17184 34529 17187
rect 32088 17156 34529 17184
rect 32088 17144 32094 17156
rect 34517 17153 34529 17156
rect 34563 17153 34575 17187
rect 34517 17147 34575 17153
rect 13863 17088 22784 17116
rect 13863 17085 13875 17088
rect 13817 17079 13875 17085
rect 25590 17076 25596 17128
rect 25648 17116 25654 17128
rect 34333 17119 34391 17125
rect 34333 17116 34345 17119
rect 25648 17088 34345 17116
rect 25648 17076 25654 17088
rect 34333 17085 34345 17088
rect 34379 17116 34391 17119
rect 34422 17116 34428 17128
rect 34379 17088 34428 17116
rect 34379 17085 34391 17088
rect 34333 17079 34391 17085
rect 34422 17076 34428 17088
rect 34480 17076 34486 17128
rect 34701 17119 34759 17125
rect 34701 17085 34713 17119
rect 34747 17116 34759 17119
rect 34790 17116 34796 17128
rect 34747 17088 34796 17116
rect 34747 17085 34759 17088
rect 34701 17079 34759 17085
rect 34790 17076 34796 17088
rect 34848 17076 34854 17128
rect 34992 17116 35020 17292
rect 36354 17280 36360 17292
rect 36412 17280 36418 17332
rect 40402 17280 40408 17332
rect 40460 17320 40466 17332
rect 75178 17320 75184 17332
rect 40460 17292 75184 17320
rect 40460 17280 40466 17292
rect 75178 17280 75184 17292
rect 75236 17280 75242 17332
rect 77938 17320 77944 17332
rect 77899 17292 77944 17320
rect 77938 17280 77944 17292
rect 77996 17280 78002 17332
rect 78030 17280 78036 17332
rect 78088 17320 78094 17332
rect 78677 17323 78735 17329
rect 78677 17320 78689 17323
rect 78088 17292 78689 17320
rect 78088 17280 78094 17292
rect 78677 17289 78689 17292
rect 78723 17289 78735 17323
rect 93946 17320 93952 17332
rect 93907 17292 93952 17320
rect 78677 17283 78735 17289
rect 93946 17280 93952 17292
rect 94004 17280 94010 17332
rect 94314 17280 94320 17332
rect 94372 17320 94378 17332
rect 94409 17323 94467 17329
rect 94409 17320 94421 17323
rect 94372 17292 94421 17320
rect 94372 17280 94378 17292
rect 94409 17289 94421 17292
rect 94455 17289 94467 17323
rect 94409 17283 94467 17289
rect 35158 17212 35164 17264
rect 35216 17252 35222 17264
rect 40954 17252 40960 17264
rect 35216 17224 40960 17252
rect 35216 17212 35222 17224
rect 40954 17212 40960 17224
rect 41012 17212 41018 17264
rect 41322 17212 41328 17264
rect 41380 17252 41386 17264
rect 43530 17252 43536 17264
rect 41380 17224 43536 17252
rect 41380 17212 41386 17224
rect 43530 17212 43536 17224
rect 43588 17212 43594 17264
rect 45278 17212 45284 17264
rect 45336 17252 45342 17264
rect 48130 17252 48136 17264
rect 45336 17224 48136 17252
rect 45336 17212 45342 17224
rect 48130 17212 48136 17224
rect 48188 17212 48194 17264
rect 72142 17252 72148 17264
rect 48240 17224 72148 17252
rect 35894 17144 35900 17196
rect 35952 17184 35958 17196
rect 46382 17184 46388 17196
rect 35952 17156 46388 17184
rect 35952 17144 35958 17156
rect 46382 17144 46388 17156
rect 46440 17144 46446 17196
rect 46566 17144 46572 17196
rect 46624 17184 46630 17196
rect 48240 17184 48268 17224
rect 72142 17212 72148 17224
rect 72200 17252 72206 17264
rect 72970 17252 72976 17264
rect 72200 17224 72976 17252
rect 72200 17212 72206 17224
rect 72970 17212 72976 17224
rect 73028 17212 73034 17264
rect 78766 17212 78772 17264
rect 78824 17252 78830 17264
rect 94041 17255 94099 17261
rect 94041 17252 94053 17255
rect 78824 17224 94053 17252
rect 78824 17212 78830 17224
rect 94041 17221 94053 17224
rect 94087 17252 94099 17255
rect 94593 17255 94651 17261
rect 94593 17252 94605 17255
rect 94087 17224 94605 17252
rect 94087 17221 94099 17224
rect 94041 17215 94099 17221
rect 94593 17221 94605 17224
rect 94639 17221 94651 17255
rect 94593 17215 94651 17221
rect 46624 17156 48268 17184
rect 46624 17144 46630 17156
rect 50706 17144 50712 17196
rect 50764 17184 50770 17196
rect 57146 17184 57152 17196
rect 50764 17156 57152 17184
rect 50764 17144 50770 17156
rect 57146 17144 57152 17156
rect 57204 17184 57210 17196
rect 64782 17184 64788 17196
rect 57204 17156 64788 17184
rect 57204 17144 57210 17156
rect 64782 17144 64788 17156
rect 64840 17144 64846 17196
rect 69290 17144 69296 17196
rect 69348 17184 69354 17196
rect 69842 17184 69848 17196
rect 69348 17156 69848 17184
rect 69348 17144 69354 17156
rect 69842 17144 69848 17156
rect 69900 17144 69906 17196
rect 94133 17187 94191 17193
rect 94133 17184 94145 17187
rect 77680 17156 78628 17184
rect 35069 17119 35127 17125
rect 35069 17116 35081 17119
rect 34992 17088 35081 17116
rect 35069 17085 35081 17088
rect 35115 17085 35127 17119
rect 35069 17079 35127 17085
rect 35250 17076 35256 17128
rect 35308 17116 35314 17128
rect 35621 17119 35679 17125
rect 35308 17088 35572 17116
rect 35308 17076 35314 17088
rect 7834 17008 7840 17060
rect 7892 17048 7898 17060
rect 8110 17048 8116 17060
rect 7892 17020 8116 17048
rect 7892 17008 7898 17020
rect 8110 17008 8116 17020
rect 8168 17048 8174 17060
rect 32030 17048 32036 17060
rect 8168 17020 32036 17048
rect 8168 17008 8174 17020
rect 32030 17008 32036 17020
rect 32088 17008 32094 17060
rect 35544 17048 35572 17088
rect 35621 17085 35633 17119
rect 35667 17116 35679 17119
rect 45554 17116 45560 17128
rect 35667 17088 45560 17116
rect 35667 17085 35679 17088
rect 35621 17079 35679 17085
rect 45554 17076 45560 17088
rect 45612 17076 45618 17128
rect 46290 17076 46296 17128
rect 46348 17116 46354 17128
rect 51350 17116 51356 17128
rect 46348 17088 51356 17116
rect 46348 17076 46354 17088
rect 51350 17076 51356 17088
rect 51408 17076 51414 17128
rect 56410 17076 56416 17128
rect 56468 17116 56474 17128
rect 57514 17116 57520 17128
rect 56468 17088 57520 17116
rect 56468 17076 56474 17088
rect 57514 17076 57520 17088
rect 57572 17076 57578 17128
rect 58710 17076 58716 17128
rect 58768 17116 58774 17128
rect 77680 17125 77708 17156
rect 77665 17119 77723 17125
rect 77665 17116 77677 17119
rect 58768 17088 77677 17116
rect 58768 17076 58774 17088
rect 77665 17085 77677 17088
rect 77711 17085 77723 17119
rect 78030 17116 78036 17128
rect 77991 17088 78036 17116
rect 77665 17079 77723 17085
rect 78030 17076 78036 17088
rect 78088 17076 78094 17128
rect 78214 17116 78220 17128
rect 78175 17088 78220 17116
rect 78214 17076 78220 17088
rect 78272 17076 78278 17128
rect 78306 17076 78312 17128
rect 78364 17116 78370 17128
rect 78490 17125 78496 17128
rect 78437 17119 78496 17125
rect 78364 17088 78409 17116
rect 78364 17076 78370 17088
rect 78437 17085 78449 17119
rect 78483 17085 78496 17119
rect 78437 17079 78496 17085
rect 78490 17076 78496 17079
rect 78548 17076 78554 17128
rect 78600 17125 78628 17156
rect 93826 17156 94145 17184
rect 78585 17119 78643 17125
rect 78585 17085 78597 17119
rect 78631 17116 78643 17119
rect 83274 17116 83280 17128
rect 78631 17088 83280 17116
rect 78631 17085 78643 17088
rect 78585 17079 78643 17085
rect 83274 17076 83280 17088
rect 83332 17076 83338 17128
rect 87506 17116 87512 17128
rect 87467 17088 87512 17116
rect 87506 17076 87512 17088
rect 87564 17076 87570 17128
rect 93581 17119 93639 17125
rect 93581 17085 93593 17119
rect 93627 17085 93639 17119
rect 93581 17079 93639 17085
rect 45094 17048 45100 17060
rect 34072 17020 35204 17048
rect 35544 17020 45100 17048
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 34072 16980 34100 17020
rect 34238 16980 34244 16992
rect 11204 16952 34100 16980
rect 34151 16952 34244 16980
rect 11204 16940 11210 16952
rect 34238 16940 34244 16952
rect 34296 16980 34302 16992
rect 35066 16980 35072 16992
rect 34296 16952 35072 16980
rect 34296 16940 34302 16952
rect 35066 16940 35072 16952
rect 35124 16940 35130 16992
rect 35176 16980 35204 17020
rect 45094 17008 45100 17020
rect 45152 17008 45158 17060
rect 49326 17008 49332 17060
rect 49384 17048 49390 17060
rect 93213 17051 93271 17057
rect 93213 17048 93225 17051
rect 49384 17020 93225 17048
rect 49384 17008 49390 17020
rect 93213 17017 93225 17020
rect 93259 17048 93271 17051
rect 93596 17048 93624 17079
rect 93259 17020 93624 17048
rect 93259 17017 93271 17020
rect 93213 17011 93271 17017
rect 93397 16983 93455 16989
rect 93397 16980 93409 16983
rect 35176 16952 93409 16980
rect 93397 16949 93409 16952
rect 93443 16980 93455 16983
rect 93826 16980 93854 17156
rect 94133 17153 94145 17156
rect 94179 17153 94191 17187
rect 94133 17147 94191 17153
rect 93443 16952 93854 16980
rect 93443 16949 93455 16952
rect 93397 16943 93455 16949
rect 1104 16890 98808 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 50326 16890
rect 50378 16838 50390 16890
rect 50442 16838 50454 16890
rect 50506 16838 50518 16890
rect 50570 16838 81046 16890
rect 81098 16838 81110 16890
rect 81162 16838 81174 16890
rect 81226 16838 81238 16890
rect 81290 16838 98808 16890
rect 1104 16816 98808 16838
rect 11606 16736 11612 16788
rect 11664 16776 11670 16788
rect 17126 16776 17132 16788
rect 11664 16748 17132 16776
rect 11664 16736 11670 16748
rect 17126 16736 17132 16748
rect 17184 16736 17190 16788
rect 40218 16776 40224 16788
rect 17236 16748 40224 16776
rect 10318 16668 10324 16720
rect 10376 16708 10382 16720
rect 17236 16708 17264 16748
rect 40218 16736 40224 16748
rect 40276 16736 40282 16788
rect 57974 16776 57980 16788
rect 46308 16748 57980 16776
rect 25590 16708 25596 16720
rect 10376 16680 17264 16708
rect 17328 16680 25596 16708
rect 10376 16668 10382 16680
rect 2958 16600 2964 16652
rect 3016 16640 3022 16652
rect 17034 16640 17040 16652
rect 3016 16612 17040 16640
rect 3016 16600 3022 16612
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 17126 16600 17132 16652
rect 17184 16640 17190 16652
rect 17328 16640 17356 16680
rect 25590 16668 25596 16680
rect 25648 16668 25654 16720
rect 26970 16668 26976 16720
rect 27028 16708 27034 16720
rect 27525 16711 27583 16717
rect 27525 16708 27537 16711
rect 27028 16680 27537 16708
rect 27028 16668 27034 16680
rect 27525 16677 27537 16680
rect 27571 16677 27583 16711
rect 28810 16708 28816 16720
rect 27525 16671 27583 16677
rect 27816 16680 28672 16708
rect 28771 16680 28816 16708
rect 20990 16640 20996 16652
rect 17184 16612 17356 16640
rect 17420 16612 20996 16640
rect 17184 16600 17190 16612
rect 16390 16464 16396 16516
rect 16448 16504 16454 16516
rect 17420 16504 17448 16612
rect 20990 16600 20996 16612
rect 21048 16640 21054 16652
rect 25682 16640 25688 16652
rect 21048 16612 25688 16640
rect 21048 16600 21054 16612
rect 25682 16600 25688 16612
rect 25740 16600 25746 16652
rect 25869 16643 25927 16649
rect 25869 16609 25881 16643
rect 25915 16640 25927 16643
rect 27816 16640 27844 16680
rect 27982 16640 27988 16652
rect 25915 16612 27844 16640
rect 27943 16612 27988 16640
rect 25915 16609 25927 16612
rect 25869 16603 25927 16609
rect 27982 16600 27988 16612
rect 28040 16600 28046 16652
rect 28644 16640 28672 16680
rect 28810 16668 28816 16680
rect 28868 16668 28874 16720
rect 28902 16668 28908 16720
rect 28960 16708 28966 16720
rect 35802 16708 35808 16720
rect 28960 16680 35808 16708
rect 28960 16668 28966 16680
rect 35802 16668 35808 16680
rect 35860 16668 35866 16720
rect 35894 16668 35900 16720
rect 35952 16708 35958 16720
rect 40034 16708 40040 16720
rect 35952 16680 40040 16708
rect 35952 16668 35958 16680
rect 40034 16668 40040 16680
rect 40092 16668 40098 16720
rect 40954 16668 40960 16720
rect 41012 16708 41018 16720
rect 41138 16708 41144 16720
rect 41012 16680 41144 16708
rect 41012 16668 41018 16680
rect 41138 16668 41144 16680
rect 41196 16708 41202 16720
rect 46308 16708 46336 16748
rect 57974 16736 57980 16748
rect 58032 16736 58038 16788
rect 58526 16736 58532 16788
rect 58584 16776 58590 16788
rect 58710 16776 58716 16788
rect 58584 16748 58716 16776
rect 58584 16736 58590 16748
rect 58710 16736 58716 16748
rect 58768 16736 58774 16788
rect 67913 16779 67971 16785
rect 67913 16776 67925 16779
rect 60706 16748 67925 16776
rect 41196 16680 41276 16708
rect 41196 16668 41202 16680
rect 30466 16640 30472 16652
rect 28644 16612 30472 16640
rect 30466 16600 30472 16612
rect 30524 16600 30530 16652
rect 30558 16600 30564 16652
rect 30616 16640 30622 16652
rect 34238 16640 34244 16652
rect 30616 16612 34244 16640
rect 30616 16600 30622 16612
rect 34238 16600 34244 16612
rect 34296 16600 34302 16652
rect 35618 16600 35624 16652
rect 35676 16640 35682 16652
rect 40402 16640 40408 16652
rect 35676 16612 40408 16640
rect 35676 16600 35682 16612
rect 40402 16600 40408 16612
rect 40460 16600 40466 16652
rect 41046 16640 41052 16652
rect 40959 16612 41052 16640
rect 41046 16600 41052 16612
rect 41104 16600 41110 16652
rect 41248 16640 41276 16680
rect 41524 16680 46336 16708
rect 41417 16643 41475 16649
rect 41417 16640 41429 16643
rect 41248 16612 41429 16640
rect 41417 16609 41429 16612
rect 41463 16609 41475 16643
rect 41417 16603 41475 16609
rect 24118 16572 24124 16584
rect 16448 16476 17448 16504
rect 17512 16544 24124 16572
rect 16448 16464 16454 16476
rect 17218 16396 17224 16448
rect 17276 16436 17282 16448
rect 17512 16436 17540 16544
rect 24118 16532 24124 16544
rect 24176 16532 24182 16584
rect 26122 16532 26128 16584
rect 26180 16581 26186 16584
rect 26180 16575 26197 16581
rect 26185 16541 26197 16575
rect 26180 16535 26197 16541
rect 26180 16532 26186 16535
rect 26510 16532 26516 16584
rect 26568 16572 26574 16584
rect 41064 16572 41092 16600
rect 41524 16572 41552 16680
rect 46382 16668 46388 16720
rect 46440 16708 46446 16720
rect 52822 16708 52828 16720
rect 46440 16680 52828 16708
rect 46440 16668 46446 16680
rect 52822 16668 52828 16680
rect 52880 16668 52886 16720
rect 57146 16708 57152 16720
rect 55876 16680 56916 16708
rect 57107 16680 57152 16708
rect 42426 16600 42432 16652
rect 42484 16640 42490 16652
rect 42484 16612 46152 16640
rect 42484 16600 42490 16612
rect 26568 16544 36400 16572
rect 41064 16544 41552 16572
rect 26568 16532 26574 16544
rect 18322 16464 18328 16516
rect 18380 16504 18386 16516
rect 25682 16504 25688 16516
rect 18380 16476 25688 16504
rect 18380 16464 18386 16476
rect 25682 16464 25688 16476
rect 25740 16464 25746 16516
rect 36262 16504 36268 16516
rect 26896 16476 36268 16504
rect 17276 16408 17540 16436
rect 17276 16396 17282 16408
rect 17770 16396 17776 16448
rect 17828 16436 17834 16448
rect 26896 16436 26924 16476
rect 36262 16464 36268 16476
rect 36320 16464 36326 16516
rect 36372 16504 36400 16544
rect 44818 16532 44824 16584
rect 44876 16572 44882 16584
rect 45278 16572 45284 16584
rect 44876 16544 45284 16572
rect 44876 16532 44882 16544
rect 45278 16532 45284 16544
rect 45336 16532 45342 16584
rect 46124 16572 46152 16612
rect 46934 16600 46940 16652
rect 46992 16640 46998 16652
rect 55876 16640 55904 16680
rect 46992 16612 55904 16640
rect 46992 16600 46998 16612
rect 56502 16600 56508 16652
rect 56560 16640 56566 16652
rect 56781 16643 56839 16649
rect 56781 16640 56793 16643
rect 56560 16612 56793 16640
rect 56560 16600 56566 16612
rect 56781 16609 56793 16612
rect 56827 16609 56839 16643
rect 56888 16640 56916 16680
rect 57146 16668 57152 16680
rect 57204 16668 57210 16720
rect 57514 16668 57520 16720
rect 57572 16708 57578 16720
rect 60090 16708 60096 16720
rect 57572 16680 60096 16708
rect 57572 16668 57578 16680
rect 60090 16668 60096 16680
rect 60148 16708 60154 16720
rect 60706 16708 60734 16748
rect 67913 16745 67925 16748
rect 67959 16745 67971 16779
rect 67913 16739 67971 16745
rect 69382 16736 69388 16788
rect 69440 16776 69446 16788
rect 69842 16776 69848 16788
rect 69440 16748 69848 16776
rect 69440 16736 69446 16748
rect 69842 16736 69848 16748
rect 69900 16736 69906 16788
rect 70366 16748 80054 16776
rect 60148 16680 60734 16708
rect 60148 16668 60154 16680
rect 61286 16668 61292 16720
rect 61344 16708 61350 16720
rect 61838 16708 61844 16720
rect 61344 16680 61844 16708
rect 61344 16668 61350 16680
rect 61838 16668 61844 16680
rect 61896 16668 61902 16720
rect 70366 16708 70394 16748
rect 65536 16680 70394 16708
rect 65536 16640 65564 16680
rect 71958 16668 71964 16720
rect 72016 16708 72022 16720
rect 78490 16708 78496 16720
rect 72016 16680 78496 16708
rect 72016 16668 72022 16680
rect 78490 16668 78496 16680
rect 78548 16668 78554 16720
rect 80026 16708 80054 16748
rect 84473 16711 84531 16717
rect 84473 16708 84485 16711
rect 80026 16680 84485 16708
rect 84473 16677 84485 16680
rect 84519 16677 84531 16711
rect 84473 16671 84531 16677
rect 67726 16640 67732 16652
rect 56888 16612 65564 16640
rect 67687 16612 67732 16640
rect 56781 16603 56839 16609
rect 67726 16600 67732 16612
rect 67784 16640 67790 16652
rect 69026 16643 69084 16649
rect 69026 16640 69038 16643
rect 67784 16612 69038 16640
rect 67784 16600 67790 16612
rect 69026 16609 69038 16612
rect 69072 16609 69084 16643
rect 69026 16603 69084 16609
rect 69293 16643 69351 16649
rect 69293 16609 69305 16643
rect 69339 16640 69351 16643
rect 69750 16640 69756 16652
rect 69339 16612 69756 16640
rect 69339 16609 69351 16612
rect 69293 16603 69351 16609
rect 69750 16600 69756 16612
rect 69808 16600 69814 16652
rect 72970 16600 72976 16652
rect 73028 16640 73034 16652
rect 84105 16643 84163 16649
rect 84105 16640 84117 16643
rect 73028 16612 84117 16640
rect 73028 16600 73034 16612
rect 84105 16609 84117 16612
rect 84151 16609 84163 16643
rect 84105 16603 84163 16609
rect 46566 16572 46572 16584
rect 46124 16544 46572 16572
rect 46566 16532 46572 16544
rect 46624 16532 46630 16584
rect 49142 16532 49148 16584
rect 49200 16572 49206 16584
rect 53742 16572 53748 16584
rect 49200 16544 53748 16572
rect 49200 16532 49206 16544
rect 53742 16532 53748 16544
rect 53800 16532 53806 16584
rect 53834 16532 53840 16584
rect 53892 16572 53898 16584
rect 53892 16544 56364 16572
rect 53892 16532 53898 16544
rect 56042 16504 56048 16516
rect 36372 16476 56048 16504
rect 56042 16464 56048 16476
rect 56100 16464 56106 16516
rect 56336 16504 56364 16544
rect 58066 16532 58072 16584
rect 58124 16572 58130 16584
rect 59078 16572 59084 16584
rect 58124 16544 59084 16572
rect 58124 16532 58130 16544
rect 59078 16532 59084 16544
rect 59136 16532 59142 16584
rect 59170 16532 59176 16584
rect 59228 16572 59234 16584
rect 65058 16572 65064 16584
rect 59228 16544 65064 16572
rect 59228 16532 59234 16544
rect 65058 16532 65064 16544
rect 65116 16532 65122 16584
rect 65242 16532 65248 16584
rect 65300 16572 65306 16584
rect 66162 16572 66168 16584
rect 65300 16544 66168 16572
rect 65300 16532 65306 16544
rect 66162 16532 66168 16544
rect 66220 16532 66226 16584
rect 94038 16504 94044 16516
rect 56336 16476 68048 16504
rect 17828 16408 26924 16436
rect 17828 16396 17834 16408
rect 27338 16396 27344 16448
rect 27396 16436 27402 16448
rect 31754 16436 31760 16448
rect 27396 16408 31760 16436
rect 27396 16396 27402 16408
rect 31754 16396 31760 16408
rect 31812 16396 31818 16448
rect 31938 16396 31944 16448
rect 31996 16436 32002 16448
rect 65518 16436 65524 16448
rect 31996 16408 65524 16436
rect 31996 16396 32002 16408
rect 65518 16396 65524 16408
rect 65576 16396 65582 16448
rect 68020 16436 68048 16476
rect 70366 16476 94044 16504
rect 70366 16436 70394 16476
rect 94038 16464 94044 16476
rect 94096 16464 94102 16516
rect 68020 16408 70394 16436
rect 70762 16396 70768 16448
rect 70820 16436 70826 16448
rect 72694 16436 72700 16448
rect 70820 16408 72700 16436
rect 70820 16396 70826 16408
rect 72694 16396 72700 16408
rect 72752 16396 72758 16448
rect 85482 16396 85488 16448
rect 85540 16436 85546 16448
rect 92014 16436 92020 16448
rect 85540 16408 92020 16436
rect 85540 16396 85546 16408
rect 92014 16396 92020 16408
rect 92072 16436 92078 16448
rect 92382 16436 92388 16448
rect 92072 16408 92388 16436
rect 92072 16396 92078 16408
rect 92382 16396 92388 16408
rect 92440 16396 92446 16448
rect 1104 16346 98808 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 65686 16346
rect 65738 16294 65750 16346
rect 65802 16294 65814 16346
rect 65866 16294 65878 16346
rect 65930 16294 96406 16346
rect 96458 16294 96470 16346
rect 96522 16294 96534 16346
rect 96586 16294 96598 16346
rect 96650 16294 98808 16346
rect 1104 16272 98808 16294
rect 6730 16232 6736 16244
rect 6691 16204 6736 16232
rect 6730 16192 6736 16204
rect 6788 16232 6794 16244
rect 7009 16235 7067 16241
rect 7009 16232 7021 16235
rect 6788 16204 7021 16232
rect 6788 16192 6794 16204
rect 7009 16201 7021 16204
rect 7055 16201 7067 16235
rect 7009 16195 7067 16201
rect 9858 16192 9864 16244
rect 9916 16232 9922 16244
rect 17218 16232 17224 16244
rect 9916 16204 17224 16232
rect 9916 16192 9922 16204
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 17328 16204 22094 16232
rect 14550 16124 14556 16176
rect 14608 16164 14614 16176
rect 17328 16164 17356 16204
rect 18322 16164 18328 16176
rect 14608 16136 17356 16164
rect 17420 16136 18328 16164
rect 14608 16124 14614 16136
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 10594 16096 10600 16108
rect 5592 16068 10600 16096
rect 5592 16056 5598 16068
rect 10594 16056 10600 16068
rect 10652 16056 10658 16108
rect 17420 16028 17448 16136
rect 18322 16124 18328 16136
rect 18380 16124 18386 16176
rect 22066 16164 22094 16204
rect 23474 16192 23480 16244
rect 23532 16232 23538 16244
rect 24394 16232 24400 16244
rect 23532 16204 24400 16232
rect 23532 16192 23538 16204
rect 24394 16192 24400 16204
rect 24452 16192 24458 16244
rect 25774 16192 25780 16244
rect 25832 16232 25838 16244
rect 25869 16235 25927 16241
rect 25869 16232 25881 16235
rect 25832 16204 25881 16232
rect 25832 16192 25838 16204
rect 25869 16201 25881 16204
rect 25915 16201 25927 16235
rect 25869 16195 25927 16201
rect 26694 16192 26700 16244
rect 26752 16232 26758 16244
rect 26752 16204 27476 16232
rect 26752 16192 26758 16204
rect 27338 16164 27344 16176
rect 22066 16136 27344 16164
rect 27338 16124 27344 16136
rect 27396 16124 27402 16176
rect 27448 16164 27476 16204
rect 29638 16192 29644 16244
rect 29696 16232 29702 16244
rect 31386 16232 31392 16244
rect 29696 16204 31392 16232
rect 29696 16192 29702 16204
rect 31386 16192 31392 16204
rect 31444 16192 31450 16244
rect 31573 16235 31631 16241
rect 31573 16201 31585 16235
rect 31619 16232 31631 16235
rect 31619 16204 31708 16232
rect 31619 16201 31631 16204
rect 31573 16195 31631 16201
rect 31297 16167 31355 16173
rect 31297 16164 31309 16167
rect 27448 16136 31309 16164
rect 31297 16133 31309 16136
rect 31343 16133 31355 16167
rect 31297 16127 31355 16133
rect 17770 16096 17776 16108
rect 17731 16068 17776 16096
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 31386 16096 31392 16108
rect 19306 16068 31392 16096
rect 19306 16040 19334 16068
rect 31386 16056 31392 16068
rect 31444 16056 31450 16108
rect 31570 16056 31576 16108
rect 31628 16096 31634 16108
rect 31680 16096 31708 16204
rect 32766 16192 32772 16244
rect 32824 16232 32830 16244
rect 39298 16232 39304 16244
rect 32824 16204 39304 16232
rect 32824 16192 32830 16204
rect 39298 16192 39304 16204
rect 39356 16192 39362 16244
rect 40218 16192 40224 16244
rect 40276 16232 40282 16244
rect 41138 16232 41144 16244
rect 40276 16204 41144 16232
rect 40276 16192 40282 16204
rect 41138 16192 41144 16204
rect 41196 16192 41202 16244
rect 48866 16232 48872 16244
rect 43456 16204 48872 16232
rect 31754 16124 31760 16176
rect 31812 16164 31818 16176
rect 32490 16164 32496 16176
rect 31812 16136 32496 16164
rect 31812 16124 31818 16136
rect 31628 16068 31708 16096
rect 31628 16056 31634 16068
rect 17524 16031 17582 16037
rect 17524 16028 17536 16031
rect 17420 16000 17536 16028
rect 17524 15997 17536 16000
rect 17570 15997 17582 16031
rect 17524 15991 17582 15997
rect 17681 16031 17739 16037
rect 17681 15997 17693 16031
rect 17727 15997 17739 16031
rect 17862 16028 17868 16040
rect 17824 16000 17868 16028
rect 17681 15991 17739 15997
rect 17313 15963 17371 15969
rect 17313 15929 17325 15963
rect 17359 15960 17371 15963
rect 17696 15960 17724 15991
rect 17862 15988 17868 16000
rect 17920 15988 17926 16040
rect 18046 16028 18052 16040
rect 18007 16000 18052 16028
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 19242 15988 19248 16040
rect 19300 16000 19334 16040
rect 19300 15988 19306 16000
rect 25682 15988 25688 16040
rect 25740 16028 25746 16040
rect 31018 16028 31024 16040
rect 25740 16000 31024 16028
rect 25740 15988 25746 16000
rect 31018 15988 31024 16000
rect 31076 15988 31082 16040
rect 31864 16037 31892 16136
rect 32490 16124 32496 16136
rect 32548 16124 32554 16176
rect 34054 16164 34060 16176
rect 34015 16136 34060 16164
rect 34054 16124 34060 16136
rect 34112 16124 34118 16176
rect 35802 16124 35808 16176
rect 35860 16164 35866 16176
rect 38194 16164 38200 16176
rect 35860 16136 38200 16164
rect 35860 16124 35866 16136
rect 38194 16124 38200 16136
rect 38252 16124 38258 16176
rect 32030 16056 32036 16108
rect 32088 16096 32094 16108
rect 43456 16096 43484 16204
rect 48866 16192 48872 16204
rect 48924 16192 48930 16244
rect 53742 16192 53748 16244
rect 53800 16232 53806 16244
rect 58986 16232 58992 16244
rect 53800 16204 58992 16232
rect 53800 16192 53806 16204
rect 58986 16192 58992 16204
rect 59044 16192 59050 16244
rect 62390 16192 62396 16244
rect 62448 16232 62454 16244
rect 64138 16232 64144 16244
rect 62448 16204 64144 16232
rect 62448 16192 62454 16204
rect 64138 16192 64144 16204
rect 64196 16192 64202 16244
rect 65426 16192 65432 16244
rect 65484 16232 65490 16244
rect 66162 16232 66168 16244
rect 65484 16204 66168 16232
rect 65484 16192 65490 16204
rect 66162 16192 66168 16204
rect 66220 16192 66226 16244
rect 66254 16192 66260 16244
rect 66312 16232 66318 16244
rect 76929 16235 76987 16241
rect 76929 16232 76941 16235
rect 66312 16204 76941 16232
rect 66312 16192 66318 16204
rect 76929 16201 76941 16204
rect 76975 16201 76987 16235
rect 76929 16195 76987 16201
rect 44266 16124 44272 16176
rect 44324 16164 44330 16176
rect 44324 16136 55904 16164
rect 44324 16124 44330 16136
rect 32088 16068 43484 16096
rect 32088 16056 32094 16068
rect 44082 16056 44088 16108
rect 44140 16096 44146 16108
rect 44140 16068 53696 16096
rect 44140 16056 44146 16068
rect 31711 16031 31769 16037
rect 31711 16028 31723 16031
rect 31404 16000 31723 16028
rect 31404 15972 31432 16000
rect 31711 15997 31723 16000
rect 31757 15997 31769 16031
rect 31711 15991 31769 15997
rect 31849 16031 31907 16037
rect 31849 15997 31861 16031
rect 31895 15997 31907 16031
rect 32122 16028 32128 16040
rect 32083 16000 32128 16028
rect 31849 15991 31907 15997
rect 32122 15988 32128 16000
rect 32180 15988 32186 16040
rect 34698 15988 34704 16040
rect 34756 16028 34762 16040
rect 37274 16028 37280 16040
rect 34756 16000 37280 16028
rect 34756 15988 34762 16000
rect 37274 15988 37280 16000
rect 37332 16028 37338 16040
rect 53282 16028 53288 16040
rect 37332 16000 53288 16028
rect 37332 15988 37338 16000
rect 53282 15988 53288 16000
rect 53340 15988 53346 16040
rect 53668 16028 53696 16068
rect 53742 16056 53748 16108
rect 53800 16096 53806 16108
rect 53926 16096 53932 16108
rect 53800 16068 53932 16096
rect 53800 16056 53806 16068
rect 53926 16056 53932 16068
rect 53984 16056 53990 16108
rect 54018 16056 54024 16108
rect 54076 16096 54082 16108
rect 55766 16096 55772 16108
rect 54076 16068 55772 16096
rect 54076 16056 54082 16068
rect 55766 16056 55772 16068
rect 55824 16056 55830 16108
rect 55876 16096 55904 16136
rect 56042 16124 56048 16176
rect 56100 16164 56106 16176
rect 62666 16164 62672 16176
rect 56100 16136 62672 16164
rect 56100 16124 56106 16136
rect 62666 16124 62672 16136
rect 62724 16124 62730 16176
rect 65518 16124 65524 16176
rect 65576 16164 65582 16176
rect 70854 16164 70860 16176
rect 65576 16136 70860 16164
rect 65576 16124 65582 16136
rect 70854 16124 70860 16136
rect 70912 16124 70918 16176
rect 63218 16096 63224 16108
rect 55876 16068 63224 16096
rect 63218 16056 63224 16068
rect 63276 16056 63282 16108
rect 65334 16056 65340 16108
rect 65392 16096 65398 16108
rect 72513 16099 72571 16105
rect 72513 16096 72525 16099
rect 65392 16068 72525 16096
rect 65392 16056 65398 16068
rect 72513 16065 72525 16068
rect 72559 16096 72571 16099
rect 73338 16096 73344 16108
rect 72559 16068 73344 16096
rect 72559 16065 72571 16068
rect 72513 16059 72571 16065
rect 73338 16056 73344 16068
rect 73396 16056 73402 16108
rect 75549 16099 75607 16105
rect 75549 16065 75561 16099
rect 75595 16096 75607 16099
rect 80054 16096 80060 16108
rect 75595 16068 80060 16096
rect 75595 16065 75607 16068
rect 75549 16059 75607 16065
rect 80054 16056 80060 16068
rect 80112 16096 80118 16108
rect 85482 16096 85488 16108
rect 80112 16068 85488 16096
rect 80112 16056 80118 16068
rect 85482 16056 85488 16068
rect 85540 16056 85546 16108
rect 56042 16028 56048 16040
rect 53668 16000 56048 16028
rect 56042 15988 56048 16000
rect 56100 15988 56106 16040
rect 56318 16028 56324 16040
rect 56279 16000 56324 16028
rect 56318 15988 56324 16000
rect 56376 15988 56382 16040
rect 56502 15988 56508 16040
rect 56560 16028 56566 16040
rect 59170 16028 59176 16040
rect 56560 16000 59176 16028
rect 56560 15988 56566 16000
rect 59170 15988 59176 16000
rect 59228 15988 59234 16040
rect 59354 15988 59360 16040
rect 59412 16028 59418 16040
rect 66165 16031 66223 16037
rect 66165 16028 66177 16031
rect 59412 16000 66177 16028
rect 59412 15988 59418 16000
rect 66165 15997 66177 16000
rect 66211 15997 66223 16031
rect 66165 15991 66223 15997
rect 69750 15988 69756 16040
rect 69808 16028 69814 16040
rect 70857 16031 70915 16037
rect 70857 16028 70869 16031
rect 69808 16000 70869 16028
rect 69808 15988 69814 16000
rect 70857 15997 70869 16000
rect 70903 15997 70915 16031
rect 71133 16031 71191 16037
rect 71133 16028 71145 16031
rect 70857 15991 70915 15997
rect 70964 16000 71145 16028
rect 18138 15960 18144 15972
rect 17359 15932 17540 15960
rect 17696 15932 18144 15960
rect 17359 15929 17371 15932
rect 17313 15923 17371 15929
rect 17218 15892 17224 15904
rect 17179 15864 17224 15892
rect 17218 15852 17224 15864
rect 17276 15852 17282 15904
rect 17512 15892 17540 15932
rect 18138 15920 18144 15932
rect 18196 15920 18202 15972
rect 31202 15960 31208 15972
rect 19306 15932 31208 15960
rect 19306 15892 19334 15932
rect 31202 15920 31208 15932
rect 31260 15920 31266 15972
rect 31386 15920 31392 15972
rect 31444 15920 31450 15972
rect 31941 15963 31999 15969
rect 31941 15960 31953 15963
rect 31496 15932 31953 15960
rect 17512 15864 19334 15892
rect 21450 15852 21456 15904
rect 21508 15892 21514 15904
rect 26878 15892 26884 15904
rect 21508 15864 26884 15892
rect 21508 15852 21514 15864
rect 26878 15852 26884 15864
rect 26936 15852 26942 15904
rect 31297 15895 31355 15901
rect 31297 15861 31309 15895
rect 31343 15892 31355 15895
rect 31496 15892 31524 15932
rect 31941 15929 31953 15932
rect 31987 15929 31999 15963
rect 31941 15923 31999 15929
rect 32030 15920 32036 15972
rect 32088 15960 32094 15972
rect 70964 15960 70992 16000
rect 71133 15997 71145 16000
rect 71179 15997 71191 16031
rect 71133 15991 71191 15997
rect 73798 15988 73804 16040
rect 73856 16028 73862 16040
rect 75825 16031 75883 16037
rect 75825 16028 75837 16031
rect 73856 16000 75837 16028
rect 73856 15988 73862 16000
rect 75825 15997 75837 16000
rect 75871 15997 75883 16031
rect 75825 15991 75883 15997
rect 32088 15932 70992 15960
rect 32088 15920 32094 15932
rect 93118 15920 93124 15972
rect 93176 15960 93182 15972
rect 97166 15960 97172 15972
rect 93176 15932 97172 15960
rect 93176 15920 93182 15932
rect 97166 15920 97172 15932
rect 97224 15920 97230 15972
rect 31343 15864 31524 15892
rect 31343 15861 31355 15864
rect 31297 15855 31355 15861
rect 31754 15852 31760 15904
rect 31812 15892 31818 15904
rect 65334 15892 65340 15904
rect 31812 15864 65340 15892
rect 31812 15852 31818 15864
rect 65334 15852 65340 15864
rect 65392 15852 65398 15904
rect 65426 15852 65432 15904
rect 65484 15892 65490 15904
rect 70762 15892 70768 15904
rect 65484 15864 70768 15892
rect 65484 15852 65490 15864
rect 70762 15852 70768 15864
rect 70820 15852 70826 15904
rect 70854 15852 70860 15904
rect 70912 15892 70918 15904
rect 72602 15892 72608 15904
rect 70912 15864 72608 15892
rect 70912 15852 70918 15864
rect 72602 15852 72608 15864
rect 72660 15852 72666 15904
rect 75914 15852 75920 15904
rect 75972 15892 75978 15904
rect 77110 15892 77116 15904
rect 75972 15864 77116 15892
rect 75972 15852 75978 15864
rect 77110 15852 77116 15864
rect 77168 15892 77174 15904
rect 84746 15892 84752 15904
rect 77168 15864 84752 15892
rect 77168 15852 77174 15864
rect 84746 15852 84752 15864
rect 84804 15852 84810 15904
rect 91738 15852 91744 15904
rect 91796 15892 91802 15904
rect 97350 15892 97356 15904
rect 91796 15864 97356 15892
rect 91796 15852 91802 15864
rect 97350 15852 97356 15864
rect 97408 15852 97414 15904
rect 1104 15802 98808 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 50326 15802
rect 50378 15750 50390 15802
rect 50442 15750 50454 15802
rect 50506 15750 50518 15802
rect 50570 15750 81046 15802
rect 81098 15750 81110 15802
rect 81162 15750 81174 15802
rect 81226 15750 81238 15802
rect 81290 15750 98808 15802
rect 1104 15728 98808 15750
rect 17494 15648 17500 15700
rect 17552 15688 17558 15700
rect 17862 15688 17868 15700
rect 17552 15660 17868 15688
rect 17552 15648 17558 15660
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 24394 15648 24400 15700
rect 24452 15688 24458 15700
rect 36078 15688 36084 15700
rect 24452 15660 36084 15688
rect 24452 15648 24458 15660
rect 36078 15648 36084 15660
rect 36136 15648 36142 15700
rect 36262 15648 36268 15700
rect 36320 15688 36326 15700
rect 41046 15688 41052 15700
rect 36320 15660 41052 15688
rect 36320 15648 36326 15660
rect 41046 15648 41052 15660
rect 41104 15648 41110 15700
rect 41322 15648 41328 15700
rect 41380 15648 41386 15700
rect 41782 15688 41788 15700
rect 41524 15660 41788 15688
rect 2958 15580 2964 15632
rect 3016 15620 3022 15632
rect 40218 15620 40224 15632
rect 3016 15592 40224 15620
rect 3016 15580 3022 15592
rect 40218 15580 40224 15592
rect 40276 15580 40282 15632
rect 40310 15580 40316 15632
rect 40368 15620 40374 15632
rect 40957 15623 41015 15629
rect 40957 15620 40969 15623
rect 40368 15592 40969 15620
rect 40368 15580 40374 15592
rect 40957 15589 40969 15592
rect 41003 15589 41015 15623
rect 40957 15583 41015 15589
rect 17037 15555 17095 15561
rect 17037 15521 17049 15555
rect 17083 15552 17095 15555
rect 17310 15552 17316 15564
rect 17083 15524 17316 15552
rect 17083 15521 17095 15524
rect 17037 15515 17095 15521
rect 17310 15512 17316 15524
rect 17368 15512 17374 15564
rect 17586 15552 17592 15564
rect 17547 15524 17592 15552
rect 17586 15512 17592 15524
rect 17644 15512 17650 15564
rect 17678 15512 17684 15564
rect 17736 15552 17742 15564
rect 17862 15552 17868 15564
rect 17736 15524 17781 15552
rect 17823 15524 17868 15552
rect 17736 15512 17742 15524
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 18414 15552 18420 15564
rect 18375 15524 18420 15552
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 18782 15552 18788 15564
rect 18743 15524 18788 15552
rect 18782 15512 18788 15524
rect 18840 15512 18846 15564
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 24026 15552 24032 15564
rect 19392 15524 24032 15552
rect 19392 15512 19398 15524
rect 24026 15512 24032 15524
rect 24084 15512 24090 15564
rect 24118 15512 24124 15564
rect 24176 15552 24182 15564
rect 30190 15552 30196 15564
rect 24176 15524 30196 15552
rect 24176 15512 24182 15524
rect 30190 15512 30196 15524
rect 30248 15552 30254 15564
rect 32122 15552 32128 15564
rect 30248 15524 32128 15552
rect 30248 15512 30254 15524
rect 32122 15512 32128 15524
rect 32180 15512 32186 15564
rect 38654 15552 38660 15564
rect 36004 15524 38660 15552
rect 7190 15444 7196 15496
rect 7248 15484 7254 15496
rect 16390 15484 16396 15496
rect 7248 15456 16396 15484
rect 7248 15444 7254 15456
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15453 17555 15487
rect 17497 15447 17555 15453
rect 8110 15376 8116 15428
rect 8168 15416 8174 15428
rect 16298 15416 16304 15428
rect 8168 15388 16304 15416
rect 8168 15376 8174 15388
rect 16298 15376 16304 15388
rect 16356 15376 16362 15428
rect 17512 15416 17540 15447
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 20438 15484 20444 15496
rect 19484 15456 20444 15484
rect 19484 15444 19490 15456
rect 20438 15444 20444 15456
rect 20496 15444 20502 15496
rect 22922 15444 22928 15496
rect 22980 15484 22986 15496
rect 36004 15484 36032 15524
rect 38654 15512 38660 15524
rect 38712 15552 38718 15564
rect 41340 15561 41368 15648
rect 41417 15623 41475 15629
rect 41417 15589 41429 15623
rect 41463 15620 41475 15623
rect 41524 15620 41552 15660
rect 41782 15648 41788 15660
rect 41840 15648 41846 15700
rect 54018 15688 54024 15700
rect 48884 15660 54024 15688
rect 41463 15592 41552 15620
rect 41463 15589 41475 15592
rect 41417 15583 41475 15589
rect 47486 15580 47492 15632
rect 47544 15620 47550 15632
rect 48884 15620 48912 15660
rect 54018 15648 54024 15660
rect 54076 15648 54082 15700
rect 55858 15648 55864 15700
rect 55916 15688 55922 15700
rect 55916 15660 58664 15688
rect 55916 15648 55922 15660
rect 47544 15592 48912 15620
rect 47544 15580 47550 15592
rect 41325 15555 41383 15561
rect 38712 15524 41276 15552
rect 38712 15512 38718 15524
rect 22980 15456 36032 15484
rect 22980 15444 22986 15456
rect 36078 15444 36084 15496
rect 36136 15484 36142 15496
rect 40402 15484 40408 15496
rect 36136 15456 40408 15484
rect 36136 15444 36142 15456
rect 40402 15444 40408 15456
rect 40460 15444 40466 15496
rect 41248 15484 41276 15524
rect 41325 15521 41337 15555
rect 41371 15521 41383 15555
rect 41506 15552 41512 15564
rect 41467 15524 41512 15552
rect 41325 15515 41383 15521
rect 41506 15512 41512 15524
rect 41564 15512 41570 15564
rect 41693 15555 41751 15561
rect 41693 15521 41705 15555
rect 41739 15552 41751 15555
rect 45370 15552 45376 15564
rect 41739 15524 45376 15552
rect 41739 15521 41751 15524
rect 41693 15515 41751 15521
rect 45370 15512 45376 15524
rect 45428 15512 45434 15564
rect 48774 15552 48780 15564
rect 48286 15524 48780 15552
rect 48286 15484 48314 15524
rect 48774 15512 48780 15524
rect 48832 15512 48838 15564
rect 48884 15561 48912 15592
rect 49053 15623 49111 15629
rect 49053 15589 49065 15623
rect 49099 15620 49111 15623
rect 53926 15620 53932 15632
rect 49099 15592 53932 15620
rect 49099 15589 49111 15592
rect 49053 15583 49111 15589
rect 53926 15580 53932 15592
rect 53984 15580 53990 15632
rect 54294 15580 54300 15632
rect 54352 15620 54358 15632
rect 54665 15623 54723 15629
rect 54665 15620 54677 15623
rect 54352 15592 54677 15620
rect 54352 15580 54358 15592
rect 54665 15589 54677 15592
rect 54711 15589 54723 15623
rect 54665 15583 54723 15589
rect 55766 15580 55772 15632
rect 55824 15620 55830 15632
rect 58066 15620 58072 15632
rect 55824 15592 58072 15620
rect 55824 15580 55830 15592
rect 58066 15580 58072 15592
rect 58124 15580 58130 15632
rect 48870 15555 48928 15561
rect 48870 15521 48882 15555
rect 48916 15521 48928 15555
rect 48870 15515 48928 15521
rect 49145 15555 49203 15561
rect 49145 15521 49157 15555
rect 49191 15521 49203 15555
rect 49145 15515 49203 15521
rect 49283 15555 49341 15561
rect 49283 15521 49295 15555
rect 49329 15552 49341 15555
rect 49602 15552 49608 15564
rect 49329 15524 49608 15552
rect 49329 15521 49341 15524
rect 49283 15515 49341 15521
rect 41248 15456 48314 15484
rect 26418 15416 26424 15428
rect 17512 15388 26424 15416
rect 26418 15376 26424 15388
rect 26476 15376 26482 15428
rect 26878 15376 26884 15428
rect 26936 15416 26942 15428
rect 49160 15416 49188 15515
rect 49602 15512 49608 15524
rect 49660 15512 49666 15564
rect 54478 15552 54484 15564
rect 49712 15524 54484 15552
rect 49712 15416 49740 15524
rect 54478 15512 54484 15524
rect 54536 15512 54542 15564
rect 54754 15552 54760 15564
rect 54715 15524 54760 15552
rect 54754 15512 54760 15524
rect 54812 15512 54818 15564
rect 54849 15555 54907 15561
rect 54849 15521 54861 15555
rect 54895 15552 54907 15555
rect 55122 15552 55128 15564
rect 54895 15524 55128 15552
rect 54895 15521 54907 15524
rect 54849 15515 54907 15521
rect 54864 15484 54892 15515
rect 55122 15512 55128 15524
rect 55180 15512 55186 15564
rect 55398 15512 55404 15564
rect 55456 15552 55462 15564
rect 56502 15552 56508 15564
rect 55456 15524 56508 15552
rect 55456 15512 55462 15524
rect 56502 15512 56508 15524
rect 56560 15512 56566 15564
rect 58526 15552 58532 15564
rect 58487 15524 58532 15552
rect 58526 15512 58532 15524
rect 58584 15512 58590 15564
rect 58636 15552 58664 15660
rect 58802 15648 58808 15700
rect 58860 15688 58866 15700
rect 58860 15660 58940 15688
rect 58860 15648 58866 15660
rect 58912 15620 58940 15660
rect 58986 15648 58992 15700
rect 59044 15688 59050 15700
rect 65426 15688 65432 15700
rect 59044 15660 65432 15688
rect 59044 15648 59050 15660
rect 65426 15648 65432 15660
rect 65484 15648 65490 15700
rect 72234 15688 72240 15700
rect 65536 15660 72240 15688
rect 65536 15620 65564 15660
rect 72234 15648 72240 15660
rect 72292 15648 72298 15700
rect 77294 15648 77300 15700
rect 77352 15688 77358 15700
rect 78214 15688 78220 15700
rect 77352 15660 78220 15688
rect 77352 15648 77358 15660
rect 78214 15648 78220 15660
rect 78272 15688 78278 15700
rect 78272 15660 80054 15688
rect 78272 15648 78278 15660
rect 58912 15592 65564 15620
rect 65610 15580 65616 15632
rect 65668 15620 65674 15632
rect 68462 15620 68468 15632
rect 65668 15592 68468 15620
rect 65668 15580 65674 15592
rect 68462 15580 68468 15592
rect 68520 15580 68526 15632
rect 69658 15620 69664 15632
rect 69032 15592 69520 15620
rect 69619 15592 69664 15620
rect 58636 15524 62528 15552
rect 26936 15388 49188 15416
rect 49298 15388 49740 15416
rect 54312 15456 54892 15484
rect 26936 15376 26942 15388
rect 17126 15348 17132 15360
rect 17087 15320 17132 15348
rect 17126 15308 17132 15320
rect 17184 15308 17190 15360
rect 17218 15308 17224 15360
rect 17276 15348 17282 15360
rect 18138 15348 18144 15360
rect 17276 15320 18144 15348
rect 17276 15308 17282 15320
rect 18138 15308 18144 15320
rect 18196 15348 18202 15360
rect 31478 15348 31484 15360
rect 18196 15320 31484 15348
rect 18196 15308 18202 15320
rect 31478 15308 31484 15320
rect 31536 15308 31542 15360
rect 32030 15308 32036 15360
rect 32088 15348 32094 15360
rect 35342 15348 35348 15360
rect 32088 15320 35348 15348
rect 32088 15308 32094 15320
rect 35342 15308 35348 15320
rect 35400 15308 35406 15360
rect 38010 15308 38016 15360
rect 38068 15348 38074 15360
rect 41141 15351 41199 15357
rect 41141 15348 41153 15351
rect 38068 15320 41153 15348
rect 38068 15308 38074 15320
rect 41141 15317 41153 15320
rect 41187 15317 41199 15351
rect 41141 15311 41199 15317
rect 41782 15308 41788 15360
rect 41840 15348 41846 15360
rect 41877 15351 41935 15357
rect 41877 15348 41889 15351
rect 41840 15320 41889 15348
rect 41840 15308 41846 15320
rect 41877 15317 41889 15320
rect 41923 15348 41935 15351
rect 47946 15348 47952 15360
rect 41923 15320 47952 15348
rect 41923 15317 41935 15320
rect 41877 15311 41935 15317
rect 47946 15308 47952 15320
rect 48004 15308 48010 15360
rect 48038 15308 48044 15360
rect 48096 15348 48102 15360
rect 49298 15348 49326 15388
rect 54312 15360 54340 15456
rect 55858 15444 55864 15496
rect 55916 15484 55922 15496
rect 58802 15484 58808 15496
rect 55916 15456 58808 15484
rect 55916 15444 55922 15456
rect 58802 15444 58808 15456
rect 58860 15444 58866 15496
rect 58986 15484 58992 15496
rect 58947 15456 58992 15484
rect 58986 15444 58992 15456
rect 59044 15444 59050 15496
rect 59170 15444 59176 15496
rect 59228 15484 59234 15496
rect 62390 15484 62396 15496
rect 59228 15456 62396 15484
rect 59228 15444 59234 15456
rect 62390 15444 62396 15456
rect 62448 15444 62454 15496
rect 62500 15484 62528 15524
rect 62942 15512 62948 15564
rect 63000 15552 63006 15564
rect 65426 15552 65432 15564
rect 63000 15524 65432 15552
rect 63000 15512 63006 15524
rect 65426 15512 65432 15524
rect 65484 15552 65490 15564
rect 69032 15552 69060 15592
rect 65484 15524 69060 15552
rect 69109 15555 69167 15561
rect 65484 15512 65490 15524
rect 69109 15521 69121 15555
rect 69155 15552 69167 15555
rect 69382 15552 69388 15564
rect 69155 15524 69388 15552
rect 69155 15521 69167 15524
rect 69109 15515 69167 15521
rect 69382 15512 69388 15524
rect 69440 15512 69446 15564
rect 69492 15552 69520 15592
rect 69658 15580 69664 15592
rect 69716 15580 69722 15632
rect 80026 15620 80054 15660
rect 84746 15648 84752 15700
rect 84804 15688 84810 15700
rect 84804 15660 89760 15688
rect 84804 15648 84810 15660
rect 80026 15592 84148 15620
rect 75914 15552 75920 15564
rect 69492 15524 75920 15552
rect 75914 15512 75920 15524
rect 75972 15512 75978 15564
rect 83918 15552 83924 15564
rect 83879 15524 83924 15552
rect 83918 15512 83924 15524
rect 83976 15512 83982 15564
rect 84120 15561 84148 15592
rect 89732 15561 89760 15660
rect 84105 15555 84163 15561
rect 84105 15521 84117 15555
rect 84151 15521 84163 15555
rect 84105 15515 84163 15521
rect 84289 15555 84347 15561
rect 84289 15521 84301 15555
rect 84335 15521 84347 15555
rect 84289 15515 84347 15521
rect 89717 15555 89775 15561
rect 89717 15521 89729 15555
rect 89763 15521 89775 15555
rect 90039 15555 90097 15561
rect 90039 15552 90051 15555
rect 89717 15515 89775 15521
rect 89824 15524 90051 15552
rect 84304 15484 84332 15515
rect 89254 15484 89260 15496
rect 62500 15456 84332 15484
rect 89215 15456 89260 15484
rect 89254 15444 89260 15456
rect 89312 15444 89318 15496
rect 55766 15376 55772 15428
rect 55824 15416 55830 15428
rect 62666 15416 62672 15428
rect 55824 15388 62672 15416
rect 55824 15376 55830 15388
rect 62666 15376 62672 15388
rect 62724 15376 62730 15428
rect 73614 15416 73620 15428
rect 62776 15388 73620 15416
rect 49418 15348 49424 15360
rect 48096 15320 49326 15348
rect 49379 15320 49424 15348
rect 48096 15308 48102 15320
rect 49418 15308 49424 15320
rect 49476 15308 49482 15360
rect 50154 15308 50160 15360
rect 50212 15348 50218 15360
rect 51074 15348 51080 15360
rect 50212 15320 51080 15348
rect 50212 15308 50218 15320
rect 51074 15308 51080 15320
rect 51132 15308 51138 15360
rect 54018 15348 54024 15360
rect 53979 15320 54024 15348
rect 54018 15308 54024 15320
rect 54076 15308 54082 15360
rect 54294 15348 54300 15360
rect 54255 15320 54300 15348
rect 54294 15308 54300 15320
rect 54352 15308 54358 15360
rect 55033 15351 55091 15357
rect 55033 15317 55045 15351
rect 55079 15348 55091 15351
rect 62776 15348 62804 15388
rect 73614 15376 73620 15388
rect 73672 15376 73678 15428
rect 83734 15416 83740 15428
rect 83695 15388 83740 15416
rect 83734 15376 83740 15388
rect 83792 15376 83798 15428
rect 89824 15360 89852 15524
rect 90039 15521 90051 15524
rect 90085 15521 90097 15555
rect 90174 15552 90180 15564
rect 90135 15524 90180 15552
rect 90039 15515 90097 15521
rect 90174 15512 90180 15524
rect 90232 15512 90238 15564
rect 55079 15320 62804 15348
rect 55079 15317 55091 15320
rect 55033 15311 55091 15317
rect 65058 15308 65064 15360
rect 65116 15348 65122 15360
rect 89806 15348 89812 15360
rect 65116 15320 89812 15348
rect 65116 15308 65122 15320
rect 89806 15308 89812 15320
rect 89864 15308 89870 15360
rect 1104 15258 98808 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 65686 15258
rect 65738 15206 65750 15258
rect 65802 15206 65814 15258
rect 65866 15206 65878 15258
rect 65930 15206 96406 15258
rect 96458 15206 96470 15258
rect 96522 15206 96534 15258
rect 96586 15206 96598 15258
rect 96650 15206 98808 15258
rect 1104 15184 98808 15206
rect 12250 15144 12256 15156
rect 12211 15116 12256 15144
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 19334 15144 19340 15156
rect 12406 15116 19340 15144
rect 7466 15036 7472 15088
rect 7524 15076 7530 15088
rect 12406 15076 12434 15116
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 19429 15147 19487 15153
rect 19429 15113 19441 15147
rect 19475 15144 19487 15147
rect 20254 15144 20260 15156
rect 19475 15116 20260 15144
rect 19475 15113 19487 15116
rect 19429 15107 19487 15113
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 24026 15104 24032 15156
rect 24084 15144 24090 15156
rect 52454 15144 52460 15156
rect 24084 15116 52460 15144
rect 24084 15104 24090 15116
rect 52454 15104 52460 15116
rect 52512 15104 52518 15156
rect 52549 15147 52607 15153
rect 52549 15113 52561 15147
rect 52595 15144 52607 15147
rect 53834 15144 53840 15156
rect 52595 15116 53840 15144
rect 52595 15113 52607 15116
rect 52549 15107 52607 15113
rect 53834 15104 53840 15116
rect 53892 15104 53898 15156
rect 55858 15104 55864 15156
rect 55916 15144 55922 15156
rect 62298 15144 62304 15156
rect 55916 15116 62304 15144
rect 55916 15104 55922 15116
rect 62298 15104 62304 15116
rect 62356 15144 62362 15156
rect 63402 15144 63408 15156
rect 62356 15116 63408 15144
rect 62356 15104 62362 15116
rect 63402 15104 63408 15116
rect 63460 15104 63466 15156
rect 68002 15104 68008 15156
rect 68060 15144 68066 15156
rect 68554 15144 68560 15156
rect 68060 15116 68560 15144
rect 68060 15104 68066 15116
rect 68554 15104 68560 15116
rect 68612 15104 68618 15156
rect 68664 15116 75040 15144
rect 7524 15048 12434 15076
rect 7524 15036 7530 15048
rect 19518 15036 19524 15088
rect 19576 15036 19582 15088
rect 19610 15036 19616 15088
rect 19668 15076 19674 15088
rect 19668 15048 19932 15076
rect 19668 15036 19674 15048
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 19536 15008 19564 15036
rect 19904 15017 19932 15048
rect 31478 15036 31484 15088
rect 31536 15076 31542 15088
rect 31938 15076 31944 15088
rect 31536 15048 31944 15076
rect 31536 15036 31542 15048
rect 31938 15036 31944 15048
rect 31996 15036 32002 15088
rect 32582 15036 32588 15088
rect 32640 15076 32646 15088
rect 37918 15076 37924 15088
rect 32640 15048 37924 15076
rect 32640 15036 32646 15048
rect 6788 14980 19564 15008
rect 19889 15011 19947 15017
rect 6788 14968 6794 14980
rect 19889 14977 19901 15011
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 20254 14968 20260 15020
rect 20312 14968 20318 15020
rect 20530 14968 20536 15020
rect 20588 15008 20594 15020
rect 33686 15008 33692 15020
rect 20588 14980 33692 15008
rect 20588 14968 20594 14980
rect 33686 14968 33692 14980
rect 33744 14968 33750 15020
rect 35912 15017 35940 15048
rect 37918 15036 37924 15048
rect 37976 15076 37982 15088
rect 41046 15076 41052 15088
rect 37976 15048 41052 15076
rect 37976 15036 37982 15048
rect 41046 15036 41052 15048
rect 41104 15036 41110 15088
rect 41138 15036 41144 15088
rect 41196 15076 41202 15088
rect 42886 15076 42892 15088
rect 41196 15048 42892 15076
rect 41196 15036 41202 15048
rect 42886 15036 42892 15048
rect 42944 15076 42950 15088
rect 45830 15076 45836 15088
rect 42944 15048 45836 15076
rect 42944 15036 42950 15048
rect 45830 15036 45836 15048
rect 45888 15076 45894 15088
rect 51166 15076 51172 15088
rect 45888 15048 51172 15076
rect 45888 15036 45894 15048
rect 51166 15036 51172 15048
rect 51224 15036 51230 15088
rect 51258 15036 51264 15088
rect 51316 15076 51322 15088
rect 55674 15076 55680 15088
rect 51316 15048 55680 15076
rect 51316 15036 51322 15048
rect 55674 15036 55680 15048
rect 55732 15036 55738 15088
rect 57946 15048 61976 15076
rect 35897 15011 35955 15017
rect 35897 14977 35909 15011
rect 35943 14977 35955 15011
rect 35897 14971 35955 14977
rect 36262 14968 36268 15020
rect 36320 15008 36326 15020
rect 51074 15008 51080 15020
rect 36320 14980 51080 15008
rect 36320 14968 36326 14980
rect 51074 14968 51080 14980
rect 51132 14968 51138 15020
rect 54754 14968 54760 15020
rect 54812 15008 54818 15020
rect 57946 15008 57974 15048
rect 54812 14980 57974 15008
rect 54812 14968 54818 14980
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14940 9459 14943
rect 9677 14943 9735 14949
rect 9677 14940 9689 14943
rect 9447 14912 9689 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 9677 14909 9689 14912
rect 9723 14940 9735 14943
rect 9858 14940 9864 14952
rect 9723 14912 9864 14940
rect 9723 14909 9735 14912
rect 9677 14903 9735 14909
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18417 14943 18475 14949
rect 18417 14940 18429 14943
rect 18012 14912 18429 14940
rect 18012 14900 18018 14912
rect 18417 14909 18429 14912
rect 18463 14909 18475 14943
rect 19521 14943 19579 14949
rect 19521 14940 19533 14943
rect 18417 14903 18475 14909
rect 18524 14912 19533 14940
rect 13078 14832 13084 14884
rect 13136 14872 13142 14884
rect 18524 14872 18552 14912
rect 19444 14884 19472 14912
rect 19521 14909 19533 14912
rect 19567 14909 19579 14943
rect 19702 14940 19708 14952
rect 19663 14912 19708 14940
rect 19521 14903 19579 14909
rect 19702 14900 19708 14912
rect 19760 14900 19766 14952
rect 19797 14943 19855 14949
rect 19797 14909 19809 14943
rect 19843 14909 19855 14943
rect 19797 14903 19855 14909
rect 20073 14943 20131 14949
rect 20073 14909 20085 14943
rect 20119 14940 20131 14943
rect 20272 14940 20300 14968
rect 22830 14940 22836 14952
rect 20119 14912 22836 14940
rect 20119 14909 20131 14912
rect 20073 14903 20131 14909
rect 18966 14872 18972 14884
rect 13136 14844 18552 14872
rect 18927 14844 18972 14872
rect 13136 14832 13142 14844
rect 18966 14832 18972 14844
rect 19024 14832 19030 14884
rect 19334 14872 19340 14884
rect 19076 14844 19340 14872
rect 9766 14764 9772 14816
rect 9824 14804 9830 14816
rect 19076 14804 19104 14844
rect 19334 14832 19340 14844
rect 19392 14832 19398 14884
rect 19426 14832 19432 14884
rect 19484 14832 19490 14884
rect 19610 14832 19616 14884
rect 19668 14832 19674 14884
rect 9824 14776 19104 14804
rect 9824 14764 9830 14776
rect 19150 14764 19156 14816
rect 19208 14804 19214 14816
rect 19628 14804 19656 14832
rect 19208 14776 19656 14804
rect 19812 14804 19840 14903
rect 22830 14900 22836 14912
rect 22888 14900 22894 14952
rect 33134 14940 33140 14952
rect 33095 14912 33140 14940
rect 33134 14900 33140 14912
rect 33192 14900 33198 14952
rect 33226 14900 33232 14952
rect 33284 14940 33290 14952
rect 34057 14943 34115 14949
rect 34057 14940 34069 14943
rect 33284 14912 34069 14940
rect 33284 14900 33290 14912
rect 34057 14909 34069 14912
rect 34103 14909 34115 14943
rect 34057 14903 34115 14909
rect 35526 14900 35532 14952
rect 35584 14940 35590 14952
rect 35712 14943 35770 14949
rect 35584 14912 35629 14940
rect 35584 14900 35590 14912
rect 35712 14909 35724 14943
rect 35758 14909 35770 14943
rect 35712 14903 35770 14909
rect 20257 14875 20315 14881
rect 20257 14841 20269 14875
rect 20303 14872 20315 14875
rect 26510 14872 26516 14884
rect 20303 14844 26516 14872
rect 20303 14841 20315 14844
rect 20257 14835 20315 14841
rect 26510 14832 26516 14844
rect 26568 14832 26574 14884
rect 26878 14832 26884 14884
rect 26936 14872 26942 14884
rect 35727 14872 35755 14903
rect 35802 14900 35808 14952
rect 35860 14940 35866 14952
rect 35860 14912 35905 14940
rect 35860 14900 35866 14912
rect 35986 14900 35992 14952
rect 36044 14940 36050 14952
rect 36081 14943 36139 14949
rect 36081 14940 36093 14943
rect 36044 14912 36093 14940
rect 36044 14900 36050 14912
rect 36081 14909 36093 14912
rect 36127 14909 36139 14943
rect 36081 14903 36139 14909
rect 36538 14900 36544 14952
rect 36596 14940 36602 14952
rect 36596 14912 41414 14940
rect 36596 14900 36602 14912
rect 26936 14844 35755 14872
rect 26936 14832 26942 14844
rect 20530 14804 20536 14816
rect 19812 14776 20536 14804
rect 19208 14764 19214 14776
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 20714 14764 20720 14816
rect 20772 14804 20778 14816
rect 36173 14807 36231 14813
rect 36173 14804 36185 14807
rect 20772 14776 36185 14804
rect 20772 14764 20778 14776
rect 36173 14773 36185 14776
rect 36219 14773 36231 14807
rect 41386 14804 41414 14912
rect 43806 14900 43812 14952
rect 43864 14940 43870 14952
rect 46106 14940 46112 14952
rect 43864 14912 46112 14940
rect 43864 14900 43870 14912
rect 46106 14900 46112 14912
rect 46164 14940 46170 14952
rect 48038 14940 48044 14952
rect 46164 14912 48044 14940
rect 46164 14900 46170 14912
rect 48038 14900 48044 14912
rect 48096 14900 48102 14952
rect 51166 14900 51172 14952
rect 51224 14940 51230 14952
rect 54294 14940 54300 14952
rect 51224 14912 54300 14940
rect 51224 14900 51230 14912
rect 54294 14900 54300 14912
rect 54352 14900 54358 14952
rect 57790 14900 57796 14952
rect 57848 14940 57854 14952
rect 58342 14940 58348 14952
rect 57848 14912 58348 14940
rect 57848 14900 57854 14912
rect 58342 14900 58348 14912
rect 58400 14900 58406 14952
rect 58434 14900 58440 14952
rect 58492 14940 58498 14952
rect 59262 14940 59268 14952
rect 58492 14912 59268 14940
rect 58492 14900 58498 14912
rect 59262 14900 59268 14912
rect 59320 14900 59326 14952
rect 59446 14900 59452 14952
rect 59504 14940 59510 14952
rect 60458 14940 60464 14952
rect 59504 14912 60464 14940
rect 59504 14900 59510 14912
rect 60458 14900 60464 14912
rect 60516 14900 60522 14952
rect 61286 14940 61292 14952
rect 60706 14912 61292 14940
rect 53650 14832 53656 14884
rect 53708 14872 53714 14884
rect 60706 14872 60734 14912
rect 61286 14900 61292 14912
rect 61344 14900 61350 14952
rect 61948 14940 61976 15048
rect 62114 15036 62120 15088
rect 62172 15076 62178 15088
rect 62758 15076 62764 15088
rect 62172 15048 62764 15076
rect 62172 15036 62178 15048
rect 62758 15036 62764 15048
rect 62816 15076 62822 15088
rect 68664 15076 68692 15116
rect 62816 15048 68692 15076
rect 69937 15079 69995 15085
rect 62816 15036 62822 15048
rect 69937 15045 69949 15079
rect 69983 15076 69995 15079
rect 70026 15076 70032 15088
rect 69983 15048 70032 15076
rect 69983 15045 69995 15048
rect 69937 15039 69995 15045
rect 70026 15036 70032 15048
rect 70084 15036 70090 15088
rect 75012 15076 75040 15116
rect 75086 15104 75092 15156
rect 75144 15144 75150 15156
rect 78490 15144 78496 15156
rect 75144 15116 78496 15144
rect 75144 15104 75150 15116
rect 78490 15104 78496 15116
rect 78548 15104 78554 15156
rect 92198 15144 92204 15156
rect 92159 15116 92204 15144
rect 92198 15104 92204 15116
rect 92256 15144 92262 15156
rect 92382 15144 92388 15156
rect 92256 15116 92388 15144
rect 92256 15104 92262 15116
rect 92382 15104 92388 15116
rect 92440 15104 92446 15156
rect 93854 15104 93860 15156
rect 93912 15144 93918 15156
rect 93949 15147 94007 15153
rect 93949 15144 93961 15147
rect 93912 15116 93961 15144
rect 93912 15104 93918 15116
rect 93949 15113 93961 15116
rect 93995 15113 94007 15147
rect 93949 15107 94007 15113
rect 77294 15076 77300 15088
rect 75012 15048 77300 15076
rect 77294 15036 77300 15048
rect 77352 15036 77358 15088
rect 62390 14968 62396 15020
rect 62448 15008 62454 15020
rect 97442 15008 97448 15020
rect 62448 14980 97448 15008
rect 62448 14968 62454 14980
rect 97442 14968 97448 14980
rect 97500 14968 97506 15020
rect 68002 14940 68008 14952
rect 61948 14912 68008 14940
rect 68002 14900 68008 14912
rect 68060 14900 68066 14952
rect 69750 14900 69756 14952
rect 69808 14940 69814 14952
rect 70029 14943 70087 14949
rect 70029 14940 70041 14943
rect 69808 14912 70041 14940
rect 69808 14900 69814 14912
rect 70029 14909 70041 14912
rect 70075 14909 70087 14943
rect 70302 14940 70308 14952
rect 70263 14912 70308 14940
rect 70029 14903 70087 14909
rect 70302 14900 70308 14912
rect 70360 14900 70366 14952
rect 71774 14900 71780 14952
rect 71832 14940 71838 14952
rect 72789 14943 72847 14949
rect 72789 14940 72801 14943
rect 71832 14912 72801 14940
rect 71832 14900 71838 14912
rect 72789 14909 72801 14912
rect 72835 14909 72847 14943
rect 92385 14943 92443 14949
rect 72789 14903 72847 14909
rect 72896 14912 80054 14940
rect 53708 14844 60734 14872
rect 61013 14875 61071 14881
rect 53708 14832 53714 14844
rect 61013 14841 61025 14875
rect 61059 14872 61071 14875
rect 62114 14872 62120 14884
rect 61059 14844 62120 14872
rect 61059 14841 61071 14844
rect 61013 14835 61071 14841
rect 62114 14832 62120 14844
rect 62172 14832 62178 14884
rect 71038 14832 71044 14884
rect 71096 14872 71102 14884
rect 71685 14875 71743 14881
rect 71685 14872 71697 14875
rect 71096 14844 71697 14872
rect 71096 14832 71102 14844
rect 71685 14841 71697 14844
rect 71731 14872 71743 14875
rect 72896 14872 72924 14912
rect 71731 14844 72924 14872
rect 73341 14875 73399 14881
rect 71731 14841 71743 14844
rect 71685 14835 71743 14841
rect 73341 14841 73353 14875
rect 73387 14872 73399 14875
rect 73430 14872 73436 14884
rect 73387 14844 73436 14872
rect 73387 14841 73399 14844
rect 73341 14835 73399 14841
rect 73430 14832 73436 14844
rect 73488 14832 73494 14884
rect 69658 14804 69664 14816
rect 41386 14776 69664 14804
rect 36173 14767 36231 14773
rect 69658 14764 69664 14776
rect 69716 14764 69722 14816
rect 80026 14804 80054 14912
rect 92385 14909 92397 14943
rect 92431 14909 92443 14943
rect 92385 14903 92443 14909
rect 92014 14832 92020 14884
rect 92072 14872 92078 14884
rect 92400 14872 92428 14903
rect 92474 14900 92480 14952
rect 92532 14940 92538 14952
rect 92661 14943 92719 14949
rect 92661 14940 92673 14943
rect 92532 14912 92673 14940
rect 92532 14900 92538 14912
rect 92661 14909 92673 14912
rect 92707 14909 92719 14943
rect 92661 14903 92719 14909
rect 92072 14844 92428 14872
rect 92072 14832 92078 14844
rect 94958 14804 94964 14816
rect 80026 14776 94964 14804
rect 94958 14764 94964 14776
rect 95016 14764 95022 14816
rect 1104 14714 98808 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 50326 14714
rect 50378 14662 50390 14714
rect 50442 14662 50454 14714
rect 50506 14662 50518 14714
rect 50570 14662 81046 14714
rect 81098 14662 81110 14714
rect 81162 14662 81174 14714
rect 81226 14662 81238 14714
rect 81290 14662 98808 14714
rect 1104 14640 98808 14662
rect 17310 14560 17316 14612
rect 17368 14600 17374 14612
rect 24578 14600 24584 14612
rect 17368 14572 24584 14600
rect 17368 14560 17374 14572
rect 24578 14560 24584 14572
rect 24636 14560 24642 14612
rect 31846 14600 31852 14612
rect 28966 14572 31754 14600
rect 31807 14572 31852 14600
rect 17678 14492 17684 14544
rect 17736 14532 17742 14544
rect 26878 14532 26884 14544
rect 17736 14504 26884 14532
rect 17736 14492 17742 14504
rect 26878 14492 26884 14504
rect 26936 14492 26942 14544
rect 5077 14467 5135 14473
rect 5077 14433 5089 14467
rect 5123 14464 5135 14467
rect 10229 14467 10287 14473
rect 5123 14436 8248 14464
rect 5123 14433 5135 14436
rect 5077 14427 5135 14433
rect 8220 14408 8248 14436
rect 10229 14433 10241 14467
rect 10275 14464 10287 14467
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 10275 14436 10425 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 10413 14433 10425 14436
rect 10459 14464 10471 14467
rect 10597 14467 10655 14473
rect 10597 14464 10609 14467
rect 10459 14436 10609 14464
rect 10459 14433 10471 14436
rect 10413 14427 10471 14433
rect 10597 14433 10609 14436
rect 10643 14464 10655 14467
rect 10781 14467 10839 14473
rect 10781 14464 10793 14467
rect 10643 14436 10793 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 10781 14433 10793 14436
rect 10827 14464 10839 14467
rect 10827 14436 11192 14464
rect 10827 14433 10839 14436
rect 10781 14427 10839 14433
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14396 5411 14399
rect 5442 14396 5448 14408
rect 5399 14368 5448 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 8202 14356 8208 14408
rect 8260 14396 8266 14408
rect 11164 14405 11192 14436
rect 18966 14424 18972 14476
rect 19024 14464 19030 14476
rect 20254 14464 20260 14476
rect 19024 14436 20260 14464
rect 19024 14424 19030 14436
rect 20254 14424 20260 14436
rect 20312 14464 20318 14476
rect 28966 14464 28994 14572
rect 30466 14464 30472 14476
rect 20312 14436 28994 14464
rect 30427 14436 30472 14464
rect 20312 14424 20318 14436
rect 30466 14424 30472 14436
rect 30524 14424 30530 14476
rect 31726 14464 31754 14572
rect 31846 14560 31852 14572
rect 31904 14560 31910 14612
rect 34698 14560 34704 14612
rect 34756 14600 34762 14612
rect 35802 14600 35808 14612
rect 34756 14572 35808 14600
rect 34756 14560 34762 14572
rect 35802 14560 35808 14572
rect 35860 14560 35866 14612
rect 37642 14560 37648 14612
rect 37700 14600 37706 14612
rect 41049 14603 41107 14609
rect 41049 14600 41061 14603
rect 37700 14572 41061 14600
rect 37700 14560 37706 14572
rect 41049 14569 41061 14572
rect 41095 14569 41107 14603
rect 41049 14563 41107 14569
rect 41138 14560 41144 14612
rect 41196 14600 41202 14612
rect 55858 14600 55864 14612
rect 41196 14572 55864 14600
rect 41196 14560 41202 14572
rect 55858 14560 55864 14572
rect 55916 14560 55922 14612
rect 56226 14560 56232 14612
rect 56284 14600 56290 14612
rect 60274 14600 60280 14612
rect 56284 14572 60136 14600
rect 60235 14572 60280 14600
rect 56284 14560 56290 14572
rect 43898 14532 43904 14544
rect 38120 14504 43904 14532
rect 38010 14464 38016 14476
rect 31726 14436 38016 14464
rect 38010 14424 38016 14436
rect 38068 14424 38074 14476
rect 10873 14399 10931 14405
rect 10873 14396 10885 14399
rect 8260 14368 10885 14396
rect 8260 14356 8266 14368
rect 10873 14365 10885 14368
rect 10919 14365 10931 14399
rect 10873 14359 10931 14365
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14396 11207 14399
rect 11195 14368 11836 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 6638 14260 6644 14272
rect 6599 14232 6644 14260
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 10888 14260 10916 14359
rect 11146 14260 11152 14272
rect 10888 14232 11152 14260
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 11808 14260 11836 14368
rect 23658 14356 23664 14408
rect 23716 14396 23722 14408
rect 30745 14399 30803 14405
rect 30745 14396 30757 14399
rect 23716 14368 30757 14396
rect 23716 14356 23722 14368
rect 30745 14365 30757 14368
rect 30791 14365 30803 14399
rect 38120 14396 38148 14504
rect 43898 14492 43904 14504
rect 43956 14492 43962 14544
rect 46382 14492 46388 14544
rect 46440 14532 46446 14544
rect 51074 14532 51080 14544
rect 46440 14504 51080 14532
rect 46440 14492 46446 14504
rect 51074 14492 51080 14504
rect 51132 14492 51138 14544
rect 52546 14532 52552 14544
rect 51184 14504 52552 14532
rect 40770 14464 40776 14476
rect 40731 14436 40776 14464
rect 40770 14424 40776 14436
rect 40828 14464 40834 14476
rect 42162 14467 42220 14473
rect 42162 14464 42174 14467
rect 40828 14436 42174 14464
rect 40828 14424 40834 14436
rect 42162 14433 42174 14436
rect 42208 14433 42220 14467
rect 42162 14427 42220 14433
rect 43162 14424 43168 14476
rect 43220 14464 43226 14476
rect 51184 14464 51212 14504
rect 52546 14492 52552 14504
rect 52604 14492 52610 14544
rect 53282 14492 53288 14544
rect 53340 14532 53346 14544
rect 53340 14504 55352 14532
rect 53340 14492 53346 14504
rect 43220 14436 51212 14464
rect 43220 14424 43226 14436
rect 51258 14424 51264 14476
rect 51316 14464 51322 14476
rect 54754 14464 54760 14476
rect 51316 14436 54760 14464
rect 51316 14424 51322 14436
rect 54754 14424 54760 14436
rect 54812 14424 54818 14476
rect 54938 14424 54944 14476
rect 54996 14464 55002 14476
rect 55324 14464 55352 14504
rect 57238 14492 57244 14544
rect 57296 14532 57302 14544
rect 57790 14532 57796 14544
rect 57296 14504 57796 14532
rect 57296 14492 57302 14504
rect 57790 14492 57796 14504
rect 57848 14532 57854 14544
rect 60108 14532 60136 14572
rect 60274 14560 60280 14572
rect 60332 14560 60338 14612
rect 63402 14560 63408 14612
rect 63460 14600 63466 14612
rect 81894 14600 81900 14612
rect 63460 14572 81900 14600
rect 63460 14560 63466 14572
rect 81894 14560 81900 14572
rect 81952 14560 81958 14612
rect 57848 14504 60044 14532
rect 60108 14504 70348 14532
rect 57848 14492 57854 14504
rect 55490 14464 55496 14476
rect 54996 14436 55260 14464
rect 55324 14436 55496 14464
rect 54996 14424 55002 14436
rect 30745 14359 30803 14365
rect 31726 14368 38148 14396
rect 42429 14399 42487 14405
rect 12437 14331 12495 14337
rect 12437 14297 12449 14331
rect 12483 14328 12495 14331
rect 12483 14300 22094 14328
rect 12483 14297 12495 14300
rect 12437 14291 12495 14297
rect 12713 14263 12771 14269
rect 12713 14260 12725 14263
rect 11808 14232 12725 14260
rect 12713 14229 12725 14232
rect 12759 14260 12771 14263
rect 12897 14263 12955 14269
rect 12897 14260 12909 14263
rect 12759 14232 12909 14260
rect 12759 14229 12771 14232
rect 12713 14223 12771 14229
rect 12897 14229 12909 14232
rect 12943 14260 12955 14263
rect 13078 14260 13084 14272
rect 12943 14232 13084 14260
rect 12943 14229 12955 14232
rect 12897 14223 12955 14229
rect 13078 14220 13084 14232
rect 13136 14220 13142 14272
rect 22066 14260 22094 14300
rect 31726 14260 31754 14368
rect 42429 14365 42441 14399
rect 42475 14396 42487 14399
rect 43530 14396 43536 14408
rect 42475 14368 43536 14396
rect 42475 14365 42487 14368
rect 42429 14359 42487 14365
rect 43530 14356 43536 14368
rect 43588 14356 43594 14408
rect 49050 14356 49056 14408
rect 49108 14396 49114 14408
rect 55122 14396 55128 14408
rect 49108 14368 55128 14396
rect 49108 14356 49114 14368
rect 55122 14356 55128 14368
rect 55180 14356 55186 14408
rect 55232 14396 55260 14436
rect 55490 14424 55496 14436
rect 55548 14464 55554 14476
rect 58710 14464 58716 14476
rect 55548 14436 58716 14464
rect 55548 14424 55554 14436
rect 58710 14424 58716 14436
rect 58768 14424 58774 14476
rect 59630 14464 59636 14476
rect 59591 14436 59636 14464
rect 59630 14424 59636 14436
rect 59688 14424 59694 14476
rect 59722 14424 59728 14476
rect 59780 14473 59786 14476
rect 60016 14473 60044 14504
rect 59780 14467 59839 14473
rect 59780 14433 59793 14467
rect 59827 14433 59839 14467
rect 59780 14427 59839 14433
rect 60001 14467 60059 14473
rect 60001 14433 60013 14467
rect 60047 14433 60059 14467
rect 60182 14464 60188 14476
rect 60143 14436 60188 14464
rect 60001 14427 60059 14433
rect 59780 14424 59786 14427
rect 60182 14424 60188 14436
rect 60240 14424 60246 14476
rect 60734 14424 60740 14476
rect 60792 14464 60798 14476
rect 63494 14464 63500 14476
rect 60792 14436 63500 14464
rect 60792 14424 60798 14436
rect 63494 14424 63500 14436
rect 63552 14424 63558 14476
rect 63678 14424 63684 14476
rect 63736 14464 63742 14476
rect 63736 14436 67634 14464
rect 63736 14424 63742 14436
rect 59909 14399 59967 14405
rect 59909 14396 59921 14399
rect 55232 14368 59921 14396
rect 59909 14365 59921 14368
rect 59955 14365 59967 14399
rect 67450 14396 67456 14408
rect 59909 14359 59967 14365
rect 61028 14368 67456 14396
rect 35250 14288 35256 14340
rect 35308 14328 35314 14340
rect 35308 14300 38654 14328
rect 35308 14288 35314 14300
rect 22066 14232 31754 14260
rect 38626 14260 38654 14300
rect 42444 14300 51396 14328
rect 42444 14260 42472 14300
rect 38626 14232 42472 14260
rect 43070 14220 43076 14272
rect 43128 14260 43134 14272
rect 43714 14260 43720 14272
rect 43128 14232 43720 14260
rect 43128 14220 43134 14232
rect 43714 14220 43720 14232
rect 43772 14220 43778 14272
rect 43898 14220 43904 14272
rect 43956 14260 43962 14272
rect 51258 14260 51264 14272
rect 43956 14232 51264 14260
rect 43956 14220 43962 14232
rect 51258 14220 51264 14232
rect 51316 14220 51322 14272
rect 51368 14260 51396 14300
rect 52454 14288 52460 14340
rect 52512 14328 52518 14340
rect 55582 14328 55588 14340
rect 52512 14300 55588 14328
rect 52512 14288 52518 14300
rect 55582 14288 55588 14300
rect 55640 14328 55646 14340
rect 60274 14328 60280 14340
rect 55640 14300 60280 14328
rect 55640 14288 55646 14300
rect 60274 14288 60280 14300
rect 60332 14288 60338 14340
rect 60458 14288 60464 14340
rect 60516 14328 60522 14340
rect 61028 14328 61056 14368
rect 67450 14356 67456 14368
rect 67508 14356 67514 14408
rect 67606 14396 67634 14436
rect 69842 14424 69848 14476
rect 69900 14464 69906 14476
rect 70213 14467 70271 14473
rect 70213 14464 70225 14467
rect 69900 14436 70225 14464
rect 69900 14424 69906 14436
rect 70213 14433 70225 14436
rect 70259 14433 70271 14467
rect 70320 14464 70348 14504
rect 70394 14492 70400 14544
rect 70452 14532 70458 14544
rect 75362 14532 75368 14544
rect 70452 14504 70497 14532
rect 70872 14504 75368 14532
rect 70452 14492 70458 14504
rect 70489 14467 70547 14473
rect 70489 14464 70501 14467
rect 70320 14436 70501 14464
rect 70213 14427 70271 14433
rect 70489 14433 70501 14436
rect 70535 14433 70547 14467
rect 70489 14427 70547 14433
rect 70633 14467 70691 14473
rect 70633 14433 70645 14467
rect 70679 14464 70691 14467
rect 70762 14464 70768 14476
rect 70679 14436 70768 14464
rect 70679 14433 70691 14436
rect 70633 14427 70691 14433
rect 70762 14424 70768 14436
rect 70820 14424 70826 14476
rect 70872 14396 70900 14504
rect 75362 14492 75368 14504
rect 75420 14492 75426 14544
rect 91922 14492 91928 14544
rect 91980 14532 91986 14544
rect 91980 14504 97028 14532
rect 91980 14492 91986 14504
rect 97000 14473 97028 14504
rect 96985 14467 97043 14473
rect 67606 14368 70900 14396
rect 72436 14436 96936 14464
rect 60516 14300 61056 14328
rect 60516 14288 60522 14300
rect 61102 14288 61108 14340
rect 61160 14328 61166 14340
rect 72436 14328 72464 14436
rect 75362 14356 75368 14408
rect 75420 14396 75426 14408
rect 96246 14396 96252 14408
rect 75420 14368 96252 14396
rect 75420 14356 75426 14368
rect 96246 14356 96252 14368
rect 96304 14356 96310 14408
rect 96706 14396 96712 14408
rect 96667 14368 96712 14396
rect 96706 14356 96712 14368
rect 96764 14356 96770 14408
rect 96908 14396 96936 14436
rect 96985 14433 96997 14467
rect 97031 14433 97043 14467
rect 96985 14427 97043 14433
rect 97166 14424 97172 14476
rect 97224 14464 97230 14476
rect 97537 14467 97595 14473
rect 97537 14464 97549 14467
rect 97224 14436 97269 14464
rect 97368 14436 97549 14464
rect 97224 14424 97230 14436
rect 97368 14396 97396 14436
rect 97537 14433 97549 14436
rect 97583 14433 97595 14467
rect 97537 14427 97595 14433
rect 96908 14368 97396 14396
rect 97445 14399 97503 14405
rect 97445 14365 97457 14399
rect 97491 14365 97503 14399
rect 97445 14359 97503 14365
rect 61160 14300 72464 14328
rect 61160 14288 61166 14300
rect 81710 14288 81716 14340
rect 81768 14328 81774 14340
rect 97460 14328 97488 14359
rect 81768 14300 97488 14328
rect 81768 14288 81774 14300
rect 60734 14260 60740 14272
rect 51368 14232 60740 14260
rect 60734 14220 60740 14232
rect 60792 14220 60798 14272
rect 60826 14220 60832 14272
rect 60884 14260 60890 14272
rect 70578 14260 70584 14272
rect 60884 14232 70584 14260
rect 60884 14220 60890 14232
rect 70578 14220 70584 14232
rect 70636 14220 70642 14272
rect 70670 14220 70676 14272
rect 70728 14260 70734 14272
rect 70765 14263 70823 14269
rect 70765 14260 70777 14263
rect 70728 14232 70777 14260
rect 70728 14220 70734 14232
rect 70765 14229 70777 14232
rect 70811 14229 70823 14263
rect 70765 14223 70823 14229
rect 72694 14220 72700 14272
rect 72752 14260 72758 14272
rect 81894 14260 81900 14272
rect 72752 14232 81900 14260
rect 72752 14220 72758 14232
rect 81894 14220 81900 14232
rect 81952 14220 81958 14272
rect 89806 14220 89812 14272
rect 89864 14260 89870 14272
rect 97258 14260 97264 14272
rect 89864 14232 97264 14260
rect 89864 14220 89870 14232
rect 97258 14220 97264 14232
rect 97316 14220 97322 14272
rect 1104 14170 98808 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 65686 14170
rect 65738 14118 65750 14170
rect 65802 14118 65814 14170
rect 65866 14118 65878 14170
rect 65930 14118 96406 14170
rect 96458 14118 96470 14170
rect 96522 14118 96534 14170
rect 96586 14118 96598 14170
rect 96650 14118 98808 14170
rect 1104 14096 98808 14118
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 31202 14056 31208 14068
rect 13136 14028 31208 14056
rect 13136 14016 13142 14028
rect 31202 14016 31208 14028
rect 31260 14016 31266 14068
rect 33962 14016 33968 14068
rect 34020 14056 34026 14068
rect 40402 14056 40408 14068
rect 34020 14028 40408 14056
rect 34020 14016 34026 14028
rect 40402 14016 40408 14028
rect 40460 14016 40466 14068
rect 40862 14056 40868 14068
rect 40823 14028 40868 14056
rect 40862 14016 40868 14028
rect 40920 14016 40926 14068
rect 44085 14059 44143 14065
rect 44085 14025 44097 14059
rect 44131 14056 44143 14059
rect 66898 14056 66904 14068
rect 44131 14028 66904 14056
rect 44131 14025 44143 14028
rect 44085 14019 44143 14025
rect 66898 14016 66904 14028
rect 66956 14016 66962 14068
rect 70578 14016 70584 14068
rect 70636 14056 70642 14068
rect 72694 14056 72700 14068
rect 70636 14028 72700 14056
rect 70636 14016 70642 14028
rect 72694 14016 72700 14028
rect 72752 14016 72758 14068
rect 73893 14059 73951 14065
rect 73893 14025 73905 14059
rect 73939 14056 73951 14059
rect 76190 14056 76196 14068
rect 73939 14028 76196 14056
rect 73939 14025 73951 14028
rect 73893 14019 73951 14025
rect 76190 14016 76196 14028
rect 76248 14016 76254 14068
rect 86218 14016 86224 14068
rect 86276 14056 86282 14068
rect 86276 14028 97028 14056
rect 86276 14016 86282 14028
rect 6638 13948 6644 14000
rect 6696 13988 6702 14000
rect 13538 13988 13544 14000
rect 6696 13960 13544 13988
rect 6696 13948 6702 13960
rect 13538 13948 13544 13960
rect 13596 13948 13602 14000
rect 32490 13948 32496 14000
rect 32548 13988 32554 14000
rect 41138 13988 41144 14000
rect 32548 13960 41144 13988
rect 32548 13948 32554 13960
rect 41138 13948 41144 13960
rect 41196 13948 41202 14000
rect 47026 13988 47032 14000
rect 41248 13960 47032 13988
rect 10318 13920 10324 13932
rect 10279 13892 10324 13920
rect 10318 13880 10324 13892
rect 10376 13880 10382 13932
rect 10594 13880 10600 13932
rect 10652 13920 10658 13932
rect 24118 13920 24124 13932
rect 10652 13892 24124 13920
rect 10652 13880 10658 13892
rect 24118 13880 24124 13892
rect 24176 13880 24182 13932
rect 40402 13880 40408 13932
rect 40460 13920 40466 13932
rect 41248 13920 41276 13960
rect 43806 13920 43812 13932
rect 40460 13892 41276 13920
rect 43548 13892 43812 13920
rect 40460 13880 40466 13892
rect 9766 13852 9772 13864
rect 9727 13824 9772 13852
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 9858 13812 9864 13864
rect 9916 13852 9922 13864
rect 42978 13852 42984 13864
rect 9916 13824 40908 13852
rect 9916 13812 9922 13824
rect 5074 13744 5080 13796
rect 5132 13784 5138 13796
rect 17218 13784 17224 13796
rect 5132 13756 17224 13784
rect 5132 13744 5138 13756
rect 17218 13744 17224 13756
rect 17276 13744 17282 13796
rect 22094 13744 22100 13796
rect 22152 13784 22158 13796
rect 22738 13784 22744 13796
rect 22152 13756 22744 13784
rect 22152 13744 22158 13756
rect 22738 13744 22744 13756
rect 22796 13744 22802 13796
rect 27338 13744 27344 13796
rect 27396 13784 27402 13796
rect 31386 13784 31392 13796
rect 27396 13756 31392 13784
rect 27396 13744 27402 13756
rect 31386 13744 31392 13756
rect 31444 13744 31450 13796
rect 36906 13744 36912 13796
rect 36964 13784 36970 13796
rect 40402 13784 40408 13796
rect 36964 13756 40408 13784
rect 36964 13744 36970 13756
rect 40402 13744 40408 13756
rect 40460 13744 40466 13796
rect 40880 13784 40908 13824
rect 41524 13824 42984 13852
rect 41524 13784 41552 13824
rect 42978 13812 42984 13824
rect 43036 13812 43042 13864
rect 43548 13861 43576 13892
rect 43806 13880 43812 13892
rect 43864 13880 43870 13932
rect 43533 13855 43591 13861
rect 43533 13821 43545 13855
rect 43579 13821 43591 13855
rect 43714 13852 43720 13864
rect 43675 13824 43720 13852
rect 43533 13815 43591 13821
rect 40880 13756 41552 13784
rect 42518 13744 42524 13796
rect 42576 13784 42582 13796
rect 43548 13784 43576 13815
rect 43714 13812 43720 13824
rect 43772 13812 43778 13864
rect 43968 13861 43996 13960
rect 47026 13948 47032 13960
rect 47084 13948 47090 14000
rect 50798 13948 50804 14000
rect 50856 13988 50862 14000
rect 58621 13991 58679 13997
rect 58621 13988 58633 13991
rect 50856 13960 58633 13988
rect 50856 13948 50862 13960
rect 58621 13957 58633 13960
rect 58667 13957 58679 13991
rect 58621 13951 58679 13957
rect 58710 13948 58716 14000
rect 58768 13988 58774 14000
rect 60826 13988 60832 14000
rect 58768 13960 60832 13988
rect 58768 13948 58774 13960
rect 60826 13948 60832 13960
rect 60884 13948 60890 14000
rect 60936 13960 73384 13988
rect 44082 13880 44088 13932
rect 44140 13920 44146 13932
rect 53098 13920 53104 13932
rect 44140 13892 53104 13920
rect 44140 13880 44146 13892
rect 53098 13880 53104 13892
rect 53156 13880 53162 13932
rect 56505 13923 56563 13929
rect 56505 13889 56517 13923
rect 56551 13889 56563 13923
rect 56505 13883 56563 13889
rect 43953 13855 44011 13861
rect 43953 13821 43965 13855
rect 43999 13821 44011 13855
rect 43953 13815 44011 13821
rect 46014 13812 46020 13864
rect 46072 13852 46078 13864
rect 46382 13852 46388 13864
rect 46072 13824 46388 13852
rect 46072 13812 46078 13824
rect 46382 13812 46388 13824
rect 46440 13812 46446 13864
rect 49510 13852 49516 13864
rect 49471 13824 49516 13852
rect 49510 13812 49516 13824
rect 49568 13812 49574 13864
rect 55401 13855 55459 13861
rect 55401 13821 55413 13855
rect 55447 13821 55459 13855
rect 55401 13815 55459 13821
rect 42576 13756 43576 13784
rect 42576 13744 42582 13756
rect 43622 13744 43628 13796
rect 43680 13784 43686 13796
rect 43809 13787 43867 13793
rect 43809 13784 43821 13787
rect 43680 13756 43821 13784
rect 43680 13744 43686 13756
rect 43809 13753 43821 13756
rect 43855 13753 43867 13787
rect 43809 13747 43867 13753
rect 45186 13744 45192 13796
rect 45244 13784 45250 13796
rect 48314 13784 48320 13796
rect 45244 13756 48320 13784
rect 45244 13744 45250 13756
rect 48314 13744 48320 13756
rect 48372 13744 48378 13796
rect 49326 13744 49332 13796
rect 49384 13784 49390 13796
rect 49602 13784 49608 13796
rect 49384 13756 49608 13784
rect 49384 13744 49390 13756
rect 49602 13744 49608 13756
rect 49660 13784 49666 13796
rect 54846 13784 54852 13796
rect 49660 13756 54852 13784
rect 49660 13744 49666 13756
rect 54846 13744 54852 13756
rect 54904 13744 54910 13796
rect 55416 13784 55444 13815
rect 55674 13812 55680 13864
rect 55732 13852 55738 13864
rect 55953 13855 56011 13861
rect 55953 13852 55965 13855
rect 55732 13824 55965 13852
rect 55732 13812 55738 13824
rect 55953 13821 55965 13824
rect 55999 13821 56011 13855
rect 55953 13815 56011 13821
rect 56042 13812 56048 13864
rect 56100 13852 56106 13864
rect 56229 13855 56287 13861
rect 56229 13852 56241 13855
rect 56100 13824 56241 13852
rect 56100 13812 56106 13824
rect 56229 13821 56241 13824
rect 56275 13821 56287 13855
rect 56229 13815 56287 13821
rect 56520 13796 56548 13883
rect 56870 13880 56876 13932
rect 56928 13920 56934 13932
rect 60936 13920 60964 13960
rect 65978 13920 65984 13932
rect 56928 13892 60964 13920
rect 65939 13892 65984 13920
rect 56928 13880 56934 13892
rect 65978 13880 65984 13892
rect 66036 13880 66042 13932
rect 66254 13880 66260 13932
rect 66312 13920 66318 13932
rect 66312 13892 66668 13920
rect 66312 13880 66318 13892
rect 58621 13855 58679 13861
rect 58621 13821 58633 13855
rect 58667 13852 58679 13855
rect 66165 13855 66223 13861
rect 66165 13852 66177 13855
rect 58667 13824 66177 13852
rect 58667 13821 58679 13824
rect 58621 13815 58679 13821
rect 66165 13821 66177 13824
rect 66211 13821 66223 13855
rect 66165 13815 66223 13821
rect 66441 13855 66499 13861
rect 66441 13821 66453 13855
rect 66487 13852 66499 13855
rect 66530 13852 66536 13864
rect 66487 13824 66536 13852
rect 66487 13821 66499 13824
rect 66441 13815 66499 13821
rect 66530 13812 66536 13824
rect 66588 13812 66594 13864
rect 66640 13852 66668 13892
rect 66898 13880 66904 13932
rect 66956 13920 66962 13932
rect 71866 13920 71872 13932
rect 66956 13892 71872 13920
rect 66956 13880 66962 13892
rect 71866 13880 71872 13892
rect 71924 13880 71930 13932
rect 72050 13880 72056 13932
rect 72108 13920 72114 13932
rect 73356 13929 73384 13960
rect 96246 13948 96252 14000
rect 96304 13988 96310 14000
rect 96433 13991 96491 13997
rect 96433 13988 96445 13991
rect 96304 13960 96445 13988
rect 96304 13948 96310 13960
rect 96433 13957 96445 13960
rect 96479 13988 96491 13991
rect 96479 13960 96844 13988
rect 96479 13957 96491 13960
rect 96433 13951 96491 13957
rect 73341 13923 73399 13929
rect 72108 13892 73108 13920
rect 72108 13880 72114 13892
rect 66640 13824 66760 13852
rect 55766 13784 55772 13796
rect 55416 13756 55772 13784
rect 55766 13744 55772 13756
rect 55824 13744 55830 13796
rect 56502 13744 56508 13796
rect 56560 13744 56566 13796
rect 57974 13744 57980 13796
rect 58032 13784 58038 13796
rect 65518 13784 65524 13796
rect 58032 13756 65524 13784
rect 58032 13744 58038 13756
rect 65518 13744 65524 13756
rect 65576 13744 65582 13796
rect 66625 13787 66683 13793
rect 66625 13784 66637 13787
rect 65628 13756 66637 13784
rect 10226 13676 10232 13728
rect 10284 13716 10290 13728
rect 62114 13716 62120 13728
rect 10284 13688 62120 13716
rect 10284 13676 10290 13688
rect 62114 13676 62120 13688
rect 62172 13676 62178 13728
rect 63678 13676 63684 13728
rect 63736 13716 63742 13728
rect 65628 13716 65656 13756
rect 66625 13753 66637 13756
rect 66671 13753 66683 13787
rect 66732 13784 66760 13824
rect 69014 13812 69020 13864
rect 69072 13852 69078 13864
rect 69937 13855 69995 13861
rect 69072 13824 69888 13852
rect 69072 13812 69078 13824
rect 69750 13784 69756 13796
rect 66732 13756 69756 13784
rect 66625 13747 66683 13753
rect 69750 13744 69756 13756
rect 69808 13744 69814 13796
rect 69860 13784 69888 13824
rect 69937 13821 69949 13855
rect 69983 13852 69995 13855
rect 70026 13852 70032 13864
rect 69983 13824 70032 13852
rect 69983 13821 69995 13824
rect 69937 13815 69995 13821
rect 70026 13812 70032 13824
rect 70084 13812 70090 13864
rect 72694 13852 72700 13864
rect 72655 13824 72700 13852
rect 72694 13812 72700 13824
rect 72752 13812 72758 13864
rect 72878 13852 72884 13864
rect 72839 13824 72884 13852
rect 72878 13812 72884 13824
rect 72936 13812 72942 13864
rect 73080 13861 73108 13892
rect 73341 13889 73353 13923
rect 73387 13889 73399 13923
rect 73341 13883 73399 13889
rect 79870 13880 79876 13932
rect 79928 13920 79934 13932
rect 96816 13929 96844 13960
rect 96801 13923 96859 13929
rect 79928 13892 82860 13920
rect 79928 13880 79934 13892
rect 73065 13855 73123 13861
rect 73065 13821 73077 13855
rect 73111 13821 73123 13855
rect 73065 13815 73123 13821
rect 73433 13855 73491 13861
rect 73433 13821 73445 13855
rect 73479 13821 73491 13855
rect 73433 13815 73491 13821
rect 81989 13855 82047 13861
rect 81989 13821 82001 13855
rect 82035 13852 82047 13855
rect 82722 13852 82728 13864
rect 82035 13824 82728 13852
rect 82035 13821 82047 13824
rect 81989 13815 82047 13821
rect 73448 13784 73476 13815
rect 82722 13812 82728 13824
rect 82780 13812 82786 13864
rect 82832 13861 82860 13892
rect 96801 13889 96813 13923
rect 96847 13889 96859 13923
rect 96801 13883 96859 13889
rect 97000 13861 97028 14028
rect 97442 14016 97448 14068
rect 97500 14056 97506 14068
rect 97813 14059 97871 14065
rect 97813 14056 97825 14059
rect 97500 14028 97825 14056
rect 97500 14016 97506 14028
rect 97813 14025 97825 14028
rect 97859 14025 97871 14059
rect 97813 14019 97871 14025
rect 97258 13920 97264 13932
rect 97219 13892 97264 13920
rect 97258 13880 97264 13892
rect 97316 13880 97322 13932
rect 82817 13855 82875 13861
rect 82817 13821 82829 13855
rect 82863 13852 82875 13855
rect 96617 13855 96675 13861
rect 96617 13852 96629 13855
rect 82863 13824 96629 13852
rect 82863 13821 82875 13824
rect 82817 13815 82875 13821
rect 96617 13821 96629 13824
rect 96663 13821 96675 13855
rect 96617 13815 96675 13821
rect 96985 13855 97043 13861
rect 96985 13821 96997 13855
rect 97031 13821 97043 13855
rect 97350 13852 97356 13864
rect 97311 13824 97356 13852
rect 96985 13815 97043 13821
rect 97350 13812 97356 13824
rect 97408 13812 97414 13864
rect 69860 13756 73476 13784
rect 63736 13688 65656 13716
rect 63736 13676 63742 13688
rect 65978 13676 65984 13728
rect 66036 13716 66042 13728
rect 66257 13719 66315 13725
rect 66257 13716 66269 13719
rect 66036 13688 66269 13716
rect 66036 13676 66042 13688
rect 66257 13685 66269 13688
rect 66303 13685 66315 13719
rect 66257 13679 66315 13685
rect 81342 13676 81348 13728
rect 81400 13716 81406 13728
rect 88518 13716 88524 13728
rect 81400 13688 88524 13716
rect 81400 13676 81406 13688
rect 88518 13676 88524 13688
rect 88576 13676 88582 13728
rect 1104 13626 98808 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 50326 13626
rect 50378 13574 50390 13626
rect 50442 13574 50454 13626
rect 50506 13574 50518 13626
rect 50570 13574 81046 13626
rect 81098 13574 81110 13626
rect 81162 13574 81174 13626
rect 81226 13574 81238 13626
rect 81290 13574 98808 13626
rect 1104 13552 98808 13574
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13538 13512 13544 13524
rect 13320 13484 13544 13512
rect 13320 13472 13326 13484
rect 13538 13472 13544 13484
rect 13596 13512 13602 13524
rect 45186 13512 45192 13524
rect 13596 13484 45192 13512
rect 13596 13472 13602 13484
rect 45186 13472 45192 13484
rect 45244 13512 45250 13524
rect 48222 13512 48228 13524
rect 45244 13484 48228 13512
rect 45244 13472 45250 13484
rect 48222 13472 48228 13484
rect 48280 13472 48286 13524
rect 49786 13472 49792 13524
rect 49844 13512 49850 13524
rect 96706 13512 96712 13524
rect 49844 13484 96712 13512
rect 49844 13472 49850 13484
rect 96706 13472 96712 13484
rect 96764 13472 96770 13524
rect 3602 13404 3608 13456
rect 3660 13444 3666 13456
rect 20438 13444 20444 13456
rect 3660 13416 20444 13444
rect 3660 13404 3666 13416
rect 20438 13404 20444 13416
rect 20496 13444 20502 13456
rect 22462 13444 22468 13456
rect 20496 13416 22468 13444
rect 20496 13404 20502 13416
rect 22462 13404 22468 13416
rect 22520 13404 22526 13456
rect 27157 13447 27215 13453
rect 27157 13413 27169 13447
rect 27203 13444 27215 13447
rect 27203 13416 27476 13444
rect 27203 13413 27215 13416
rect 27157 13407 27215 13413
rect 26786 13336 26792 13388
rect 26844 13376 26850 13388
rect 26881 13379 26939 13385
rect 26881 13376 26893 13379
rect 26844 13348 26893 13376
rect 26844 13336 26850 13348
rect 26881 13345 26893 13348
rect 26927 13345 26939 13379
rect 27062 13376 27068 13388
rect 27023 13348 27068 13376
rect 26881 13339 26939 13345
rect 27062 13336 27068 13348
rect 27120 13336 27126 13388
rect 27246 13376 27252 13388
rect 27207 13348 27252 13376
rect 27246 13336 27252 13348
rect 27304 13336 27310 13388
rect 27448 13376 27476 13416
rect 27706 13404 27712 13456
rect 27764 13444 27770 13456
rect 39022 13444 39028 13456
rect 27764 13416 39028 13444
rect 27764 13404 27770 13416
rect 39022 13404 39028 13416
rect 39080 13444 39086 13456
rect 39080 13416 42012 13444
rect 39080 13404 39086 13416
rect 33778 13376 33784 13388
rect 27448 13348 33784 13376
rect 33778 13336 33784 13348
rect 33836 13336 33842 13388
rect 36722 13336 36728 13388
rect 36780 13376 36786 13388
rect 39390 13376 39396 13388
rect 36780 13348 39396 13376
rect 36780 13336 36786 13348
rect 39390 13336 39396 13348
rect 39448 13376 39454 13388
rect 39758 13376 39764 13388
rect 39448 13348 39764 13376
rect 39448 13336 39454 13348
rect 39758 13336 39764 13348
rect 39816 13336 39822 13388
rect 41984 13376 42012 13416
rect 45922 13404 45928 13456
rect 45980 13444 45986 13456
rect 62574 13444 62580 13456
rect 45980 13416 62580 13444
rect 45980 13404 45986 13416
rect 62574 13404 62580 13416
rect 62632 13444 62638 13456
rect 65978 13444 65984 13456
rect 62632 13416 65984 13444
rect 62632 13404 62638 13416
rect 65978 13404 65984 13416
rect 66036 13404 66042 13456
rect 66162 13404 66168 13456
rect 66220 13444 66226 13456
rect 66220 13416 75224 13444
rect 66220 13404 66226 13416
rect 41984 13348 65104 13376
rect 12986 13268 12992 13320
rect 13044 13308 13050 13320
rect 16942 13308 16948 13320
rect 13044 13280 16948 13308
rect 13044 13268 13050 13280
rect 16942 13268 16948 13280
rect 17000 13308 17006 13320
rect 42794 13308 42800 13320
rect 17000 13280 42800 13308
rect 17000 13268 17006 13280
rect 42794 13268 42800 13280
rect 42852 13308 42858 13320
rect 64966 13308 64972 13320
rect 42852 13280 64972 13308
rect 42852 13268 42858 13280
rect 64966 13268 64972 13280
rect 65024 13268 65030 13320
rect 65076 13308 65104 13348
rect 65518 13336 65524 13388
rect 65576 13376 65582 13388
rect 71774 13376 71780 13388
rect 65576 13348 71780 13376
rect 65576 13336 65582 13348
rect 71774 13336 71780 13348
rect 71832 13336 71838 13388
rect 72786 13376 72792 13388
rect 72747 13348 72792 13376
rect 72786 13336 72792 13348
rect 72844 13336 72850 13388
rect 72970 13336 72976 13388
rect 73028 13376 73034 13388
rect 73157 13379 73215 13385
rect 73157 13376 73169 13379
rect 73028 13348 73169 13376
rect 73028 13336 73034 13348
rect 73157 13345 73169 13348
rect 73203 13345 73215 13379
rect 75196 13376 75224 13416
rect 75362 13404 75368 13456
rect 75420 13444 75426 13456
rect 85666 13444 85672 13456
rect 75420 13416 85672 13444
rect 75420 13404 75426 13416
rect 85666 13404 85672 13416
rect 85724 13404 85730 13456
rect 83090 13385 83096 13388
rect 83047 13379 83096 13385
rect 75196 13348 80054 13376
rect 73157 13339 73215 13345
rect 69106 13308 69112 13320
rect 65076 13280 69112 13308
rect 69106 13268 69112 13280
rect 69164 13268 69170 13320
rect 70118 13268 70124 13320
rect 70176 13308 70182 13320
rect 75730 13308 75736 13320
rect 70176 13280 75736 13308
rect 70176 13268 70182 13280
rect 75730 13268 75736 13280
rect 75788 13268 75794 13320
rect 80026 13308 80054 13348
rect 83047 13345 83059 13379
rect 83093 13345 83096 13379
rect 83047 13339 83096 13345
rect 83090 13336 83096 13339
rect 83148 13336 83154 13388
rect 83277 13311 83335 13317
rect 83277 13308 83289 13311
rect 80026 13280 83289 13308
rect 83277 13277 83289 13280
rect 83323 13277 83335 13311
rect 83277 13271 83335 13277
rect 83366 13268 83372 13320
rect 83424 13308 83430 13320
rect 95237 13311 95295 13317
rect 95237 13308 95249 13311
rect 83424 13280 95249 13308
rect 83424 13268 83430 13280
rect 95237 13277 95249 13280
rect 95283 13277 95295 13311
rect 95237 13271 95295 13277
rect 13078 13200 13084 13252
rect 13136 13240 13142 13252
rect 44634 13240 44640 13252
rect 13136 13212 44640 13240
rect 13136 13200 13142 13212
rect 44634 13200 44640 13212
rect 44692 13200 44698 13252
rect 49234 13200 49240 13252
rect 49292 13240 49298 13252
rect 49786 13240 49792 13252
rect 49292 13212 49792 13240
rect 49292 13200 49298 13212
rect 49786 13200 49792 13212
rect 49844 13200 49850 13252
rect 54294 13200 54300 13252
rect 54352 13240 54358 13252
rect 81342 13240 81348 13252
rect 54352 13212 81348 13240
rect 54352 13200 54358 13212
rect 81342 13200 81348 13212
rect 81400 13200 81406 13252
rect 81544 13212 82952 13240
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 16022 13172 16028 13184
rect 12952 13144 16028 13172
rect 12952 13132 12958 13144
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 20530 13132 20536 13184
rect 20588 13172 20594 13184
rect 27433 13175 27491 13181
rect 27433 13172 27445 13175
rect 20588 13144 27445 13172
rect 20588 13132 20594 13144
rect 27433 13141 27445 13144
rect 27479 13141 27491 13175
rect 27433 13135 27491 13141
rect 28626 13132 28632 13184
rect 28684 13172 28690 13184
rect 36722 13172 36728 13184
rect 28684 13144 36728 13172
rect 28684 13132 28690 13144
rect 36722 13132 36728 13144
rect 36780 13132 36786 13184
rect 36998 13132 37004 13184
rect 37056 13172 37062 13184
rect 46382 13172 46388 13184
rect 37056 13144 46388 13172
rect 37056 13132 37062 13144
rect 46382 13132 46388 13144
rect 46440 13132 46446 13184
rect 52089 13175 52147 13181
rect 52089 13141 52101 13175
rect 52135 13172 52147 13175
rect 81544 13172 81572 13212
rect 52135 13144 81572 13172
rect 81621 13175 81679 13181
rect 52135 13141 52147 13144
rect 52089 13135 52147 13141
rect 81621 13141 81633 13175
rect 81667 13172 81679 13175
rect 82078 13172 82084 13184
rect 81667 13144 82084 13172
rect 81667 13141 81679 13144
rect 81621 13135 81679 13141
rect 82078 13132 82084 13144
rect 82136 13132 82142 13184
rect 82924 13172 82952 13212
rect 93946 13172 93952 13184
rect 82924 13144 93952 13172
rect 93946 13132 93952 13144
rect 94004 13132 94010 13184
rect 1104 13082 98808 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 65686 13082
rect 65738 13030 65750 13082
rect 65802 13030 65814 13082
rect 65866 13030 65878 13082
rect 65930 13030 96406 13082
rect 96458 13030 96470 13082
rect 96522 13030 96534 13082
rect 96586 13030 96598 13082
rect 96650 13030 98808 13082
rect 1104 13008 98808 13030
rect 22094 12968 22100 12980
rect 13096 12940 22100 12968
rect 7926 12832 7932 12844
rect 7887 12804 7932 12832
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 13096 12841 13124 12940
rect 22094 12928 22100 12940
rect 22152 12928 22158 12980
rect 22370 12968 22376 12980
rect 22331 12940 22376 12968
rect 22370 12928 22376 12940
rect 22428 12968 22434 12980
rect 23014 12968 23020 12980
rect 22428 12940 23020 12968
rect 22428 12928 22434 12940
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 30374 12928 30380 12980
rect 30432 12968 30438 12980
rect 40402 12968 40408 12980
rect 30432 12940 40408 12968
rect 30432 12928 30438 12940
rect 40402 12928 40408 12940
rect 40460 12928 40466 12980
rect 41386 12940 51074 12968
rect 17218 12860 17224 12912
rect 17276 12900 17282 12912
rect 28626 12900 28632 12912
rect 17276 12872 28632 12900
rect 17276 12860 17282 12872
rect 28626 12860 28632 12872
rect 28684 12860 28690 12912
rect 31386 12860 31392 12912
rect 31444 12900 31450 12912
rect 41386 12900 41414 12940
rect 31444 12872 41414 12900
rect 51046 12900 51074 12940
rect 52822 12928 52828 12980
rect 52880 12968 52886 12980
rect 54846 12968 54852 12980
rect 52880 12940 54852 12968
rect 52880 12928 52886 12940
rect 54846 12928 54852 12940
rect 54904 12928 54910 12980
rect 55122 12928 55128 12980
rect 55180 12968 55186 12980
rect 75362 12968 75368 12980
rect 55180 12940 75368 12968
rect 55180 12928 55186 12940
rect 75362 12928 75368 12940
rect 75420 12928 75426 12980
rect 75454 12928 75460 12980
rect 75512 12968 75518 12980
rect 75512 12940 75776 12968
rect 75512 12928 75518 12940
rect 60458 12900 60464 12912
rect 51046 12872 60464 12900
rect 31444 12860 31450 12872
rect 60458 12860 60464 12872
rect 60516 12860 60522 12912
rect 65058 12860 65064 12912
rect 65116 12900 65122 12912
rect 65242 12900 65248 12912
rect 65116 12872 65248 12900
rect 65116 12860 65122 12872
rect 65242 12860 65248 12872
rect 65300 12860 65306 12912
rect 66438 12860 66444 12912
rect 66496 12900 66502 12912
rect 67174 12900 67180 12912
rect 66496 12872 67180 12900
rect 66496 12860 66502 12872
rect 67174 12860 67180 12872
rect 67232 12860 67238 12912
rect 69750 12860 69756 12912
rect 69808 12900 69814 12912
rect 75748 12900 75776 12940
rect 79686 12928 79692 12980
rect 79744 12968 79750 12980
rect 79744 12940 93854 12968
rect 79744 12928 79750 12940
rect 85574 12900 85580 12912
rect 69808 12872 71360 12900
rect 75748 12872 85580 12900
rect 69808 12860 69814 12872
rect 12621 12835 12679 12841
rect 12621 12801 12633 12835
rect 12667 12832 12679 12835
rect 13081 12835 13139 12841
rect 12667 12804 12940 12832
rect 12667 12801 12679 12804
rect 12621 12795 12679 12801
rect 7650 12764 7656 12776
rect 7563 12736 7656 12764
rect 7650 12724 7656 12736
rect 7708 12764 7714 12776
rect 8202 12764 8208 12776
rect 7708 12736 8208 12764
rect 7708 12724 7714 12736
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 12710 12724 12716 12776
rect 12768 12724 12774 12776
rect 12912 12773 12940 12804
rect 13081 12801 13093 12835
rect 13127 12801 13139 12835
rect 17402 12832 17408 12844
rect 13081 12795 13139 12801
rect 13280 12804 17408 12832
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12764 12955 12767
rect 12986 12764 12992 12776
rect 12943 12736 12992 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 13280 12773 13308 12804
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 39114 12832 39120 12844
rect 22066 12804 39120 12832
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12733 13231 12767
rect 13173 12727 13231 12733
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12733 13323 12767
rect 13265 12727 13323 12733
rect 13449 12767 13507 12773
rect 13449 12733 13461 12767
rect 13495 12764 13507 12767
rect 22066 12764 22094 12804
rect 39114 12792 39120 12804
rect 39172 12792 39178 12844
rect 39666 12792 39672 12844
rect 39724 12832 39730 12844
rect 43162 12832 43168 12844
rect 39724 12804 43168 12832
rect 39724 12792 39730 12804
rect 43162 12792 43168 12804
rect 43220 12792 43226 12844
rect 43441 12835 43499 12841
rect 43441 12801 43453 12835
rect 43487 12832 43499 12835
rect 43806 12832 43812 12844
rect 43487 12804 43812 12832
rect 43487 12801 43499 12804
rect 43441 12795 43499 12801
rect 43806 12792 43812 12804
rect 43864 12792 43870 12844
rect 46382 12792 46388 12844
rect 46440 12832 46446 12844
rect 63678 12832 63684 12844
rect 46440 12804 63684 12832
rect 46440 12792 46446 12804
rect 63678 12792 63684 12804
rect 63736 12792 63742 12844
rect 71332 12841 71360 12872
rect 85574 12860 85580 12872
rect 85632 12860 85638 12912
rect 86926 12872 89714 12900
rect 71317 12835 71375 12841
rect 65536 12804 70348 12832
rect 13495 12736 22094 12764
rect 13495 12733 13507 12736
rect 13449 12727 13507 12733
rect 9309 12699 9367 12705
rect 9309 12665 9321 12699
rect 9355 12696 9367 12699
rect 12728 12696 12756 12724
rect 13078 12696 13084 12708
rect 9355 12668 13084 12696
rect 9355 12665 9367 12668
rect 9309 12659 9367 12665
rect 13078 12656 13084 12668
rect 13136 12656 13142 12708
rect 13188 12696 13216 12727
rect 22554 12724 22560 12776
rect 22612 12764 22618 12776
rect 22741 12767 22799 12773
rect 22741 12764 22753 12767
rect 22612 12736 22753 12764
rect 22612 12724 22618 12736
rect 22741 12733 22753 12736
rect 22787 12733 22799 12767
rect 23014 12764 23020 12776
rect 22975 12736 23020 12764
rect 22741 12727 22799 12733
rect 23014 12724 23020 12736
rect 23072 12724 23078 12776
rect 39574 12764 39580 12776
rect 23860 12736 39580 12764
rect 23860 12696 23888 12736
rect 39574 12724 39580 12736
rect 39632 12724 39638 12776
rect 39758 12724 39764 12776
rect 39816 12764 39822 12776
rect 39816 12736 41414 12764
rect 39816 12724 39822 12736
rect 13188 12668 23888 12696
rect 31018 12656 31024 12708
rect 31076 12696 31082 12708
rect 40310 12696 40316 12708
rect 31076 12668 40316 12696
rect 31076 12656 31082 12668
rect 40310 12656 40316 12668
rect 40368 12656 40374 12708
rect 41386 12696 41414 12736
rect 42426 12724 42432 12776
rect 42484 12764 42490 12776
rect 43530 12764 43536 12776
rect 42484 12736 43536 12764
rect 42484 12724 42490 12736
rect 43530 12724 43536 12736
rect 43588 12724 43594 12776
rect 43640 12736 46152 12764
rect 43640 12696 43668 12736
rect 41386 12668 43668 12696
rect 12713 12631 12771 12637
rect 12713 12597 12725 12631
rect 12759 12628 12771 12631
rect 13814 12628 13820 12640
rect 12759 12600 13820 12628
rect 12759 12597 12771 12600
rect 12713 12591 12771 12597
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 17218 12628 17224 12640
rect 16908 12600 17224 12628
rect 16908 12588 16914 12600
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 21542 12588 21548 12640
rect 21600 12628 21606 12640
rect 24210 12628 24216 12640
rect 21600 12600 24216 12628
rect 21600 12588 21606 12600
rect 24210 12588 24216 12600
rect 24268 12588 24274 12640
rect 39114 12588 39120 12640
rect 39172 12628 39178 12640
rect 42242 12628 42248 12640
rect 39172 12600 42248 12628
rect 39172 12588 39178 12600
rect 42242 12588 42248 12600
rect 42300 12588 42306 12640
rect 44634 12588 44640 12640
rect 44692 12628 44698 12640
rect 44913 12631 44971 12637
rect 44913 12628 44925 12631
rect 44692 12600 44925 12628
rect 44692 12588 44698 12600
rect 44913 12597 44925 12600
rect 44959 12597 44971 12631
rect 46124 12628 46152 12736
rect 48222 12724 48228 12776
rect 48280 12764 48286 12776
rect 48280 12736 54616 12764
rect 48280 12724 48286 12736
rect 46566 12656 46572 12708
rect 46624 12696 46630 12708
rect 54294 12696 54300 12708
rect 46624 12668 54300 12696
rect 46624 12656 46630 12668
rect 54294 12656 54300 12668
rect 54352 12656 54358 12708
rect 54588 12696 54616 12736
rect 55766 12724 55772 12776
rect 55824 12764 55830 12776
rect 65536 12764 65564 12804
rect 66162 12764 66168 12776
rect 55824 12736 65564 12764
rect 65904 12736 66168 12764
rect 55824 12724 55830 12736
rect 58618 12696 58624 12708
rect 54588 12668 58624 12696
rect 58618 12656 58624 12668
rect 58676 12656 58682 12708
rect 60550 12656 60556 12708
rect 60608 12696 60614 12708
rect 61746 12696 61752 12708
rect 60608 12668 61752 12696
rect 60608 12656 60614 12668
rect 61746 12656 61752 12668
rect 61804 12656 61810 12708
rect 61838 12656 61844 12708
rect 61896 12696 61902 12708
rect 65426 12696 65432 12708
rect 61896 12668 65432 12696
rect 61896 12656 61902 12668
rect 65426 12656 65432 12668
rect 65484 12696 65490 12708
rect 65904 12696 65932 12736
rect 66162 12724 66168 12736
rect 66220 12724 66226 12776
rect 66438 12764 66444 12776
rect 66399 12736 66444 12764
rect 66438 12724 66444 12736
rect 66496 12724 66502 12776
rect 65484 12668 65932 12696
rect 65484 12656 65490 12668
rect 65978 12656 65984 12708
rect 66036 12696 66042 12708
rect 66809 12699 66867 12705
rect 66809 12696 66821 12699
rect 66036 12668 66821 12696
rect 66036 12656 66042 12668
rect 66809 12665 66821 12668
rect 66855 12696 66867 12699
rect 69842 12696 69848 12708
rect 66855 12668 69848 12696
rect 66855 12665 66867 12668
rect 66809 12659 66867 12665
rect 69842 12656 69848 12668
rect 69900 12656 69906 12708
rect 70210 12628 70216 12640
rect 46124 12600 70216 12628
rect 44913 12591 44971 12597
rect 70210 12588 70216 12600
rect 70268 12588 70274 12640
rect 70320 12628 70348 12804
rect 71317 12801 71329 12835
rect 71363 12801 71375 12835
rect 71317 12795 71375 12801
rect 85209 12835 85267 12841
rect 85209 12801 85221 12835
rect 85255 12832 85267 12835
rect 85761 12835 85819 12841
rect 85761 12832 85773 12835
rect 85255 12804 85773 12832
rect 85255 12801 85267 12804
rect 85209 12795 85267 12801
rect 85761 12801 85773 12804
rect 85807 12832 85819 12835
rect 86313 12835 86371 12841
rect 86313 12832 86325 12835
rect 85807 12804 86325 12832
rect 85807 12801 85819 12804
rect 85761 12795 85819 12801
rect 86313 12801 86325 12804
rect 86359 12832 86371 12835
rect 86926 12832 86954 12872
rect 86359 12804 86954 12832
rect 86359 12801 86371 12804
rect 86313 12795 86371 12801
rect 71590 12764 71596 12776
rect 71551 12736 71596 12764
rect 71590 12724 71596 12736
rect 71648 12724 71654 12776
rect 71682 12724 71688 12776
rect 71740 12764 71746 12776
rect 71740 12736 72280 12764
rect 71740 12724 71746 12736
rect 72252 12696 72280 12736
rect 72418 12724 72424 12776
rect 72476 12764 72482 12776
rect 75454 12764 75460 12776
rect 72476 12736 75460 12764
rect 72476 12724 72482 12736
rect 75454 12724 75460 12736
rect 75512 12724 75518 12776
rect 75641 12767 75699 12773
rect 75641 12733 75653 12767
rect 75687 12733 75699 12767
rect 75641 12727 75699 12733
rect 75656 12696 75684 12727
rect 81894 12724 81900 12776
rect 81952 12764 81958 12776
rect 85485 12767 85543 12773
rect 85485 12764 85497 12767
rect 81952 12736 85497 12764
rect 81952 12724 81958 12736
rect 85485 12733 85497 12736
rect 85531 12733 85543 12767
rect 85485 12727 85543 12733
rect 85574 12724 85580 12776
rect 85632 12764 85638 12776
rect 85669 12767 85727 12773
rect 85669 12764 85681 12767
rect 85632 12736 85681 12764
rect 85632 12724 85638 12736
rect 85669 12733 85681 12736
rect 85715 12733 85727 12767
rect 85850 12764 85856 12776
rect 85811 12736 85856 12764
rect 85669 12727 85727 12733
rect 85850 12724 85856 12736
rect 85908 12724 85914 12776
rect 86034 12764 86040 12776
rect 85995 12736 86040 12764
rect 86034 12724 86040 12736
rect 86092 12724 86098 12776
rect 72252 12668 75684 12696
rect 75730 12656 75736 12708
rect 75788 12696 75794 12708
rect 86221 12699 86279 12705
rect 86221 12696 86233 12699
rect 75788 12668 86233 12696
rect 75788 12656 75794 12668
rect 86221 12665 86233 12668
rect 86267 12665 86279 12699
rect 86221 12659 86279 12665
rect 72697 12631 72755 12637
rect 72697 12628 72709 12631
rect 70320 12600 72709 12628
rect 72697 12597 72709 12600
rect 72743 12597 72755 12631
rect 75454 12628 75460 12640
rect 75415 12600 75460 12628
rect 72697 12591 72755 12597
rect 75454 12588 75460 12600
rect 75512 12588 75518 12640
rect 75914 12588 75920 12640
rect 75972 12628 75978 12640
rect 85209 12631 85267 12637
rect 85209 12628 85221 12631
rect 75972 12600 85221 12628
rect 75972 12588 75978 12600
rect 85209 12597 85221 12600
rect 85255 12597 85267 12631
rect 85390 12628 85396 12640
rect 85303 12600 85396 12628
rect 85209 12591 85267 12597
rect 85390 12588 85396 12600
rect 85448 12628 85454 12640
rect 85666 12628 85672 12640
rect 85448 12600 85672 12628
rect 85448 12588 85454 12600
rect 85666 12588 85672 12600
rect 85724 12628 85730 12640
rect 85850 12628 85856 12640
rect 85724 12600 85856 12628
rect 85724 12588 85730 12600
rect 85850 12588 85856 12600
rect 85908 12588 85914 12640
rect 89686 12628 89714 12872
rect 93826 12764 93854 12940
rect 96525 12767 96583 12773
rect 96525 12764 96537 12767
rect 93826 12736 96537 12764
rect 96525 12733 96537 12736
rect 96571 12733 96583 12767
rect 96525 12727 96583 12733
rect 90634 12628 90640 12640
rect 89686 12600 90640 12628
rect 90634 12588 90640 12600
rect 90692 12588 90698 12640
rect 1104 12538 98808 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 50326 12538
rect 50378 12486 50390 12538
rect 50442 12486 50454 12538
rect 50506 12486 50518 12538
rect 50570 12486 81046 12538
rect 81098 12486 81110 12538
rect 81162 12486 81174 12538
rect 81226 12486 81238 12538
rect 81290 12486 98808 12538
rect 1104 12464 98808 12486
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 38194 12424 38200 12436
rect 7064 12396 38200 12424
rect 7064 12384 7070 12396
rect 38194 12384 38200 12396
rect 38252 12424 38258 12436
rect 38562 12424 38568 12436
rect 38252 12396 38568 12424
rect 38252 12384 38258 12396
rect 38562 12384 38568 12396
rect 38620 12384 38626 12436
rect 38948 12396 54800 12424
rect 10778 12316 10784 12368
rect 10836 12356 10842 12368
rect 20438 12356 20444 12368
rect 10836 12328 20444 12356
rect 10836 12316 10842 12328
rect 20438 12316 20444 12328
rect 20496 12316 20502 12368
rect 35342 12356 35348 12368
rect 22066 12328 35348 12356
rect 10597 12291 10655 12297
rect 10597 12257 10609 12291
rect 10643 12288 10655 12291
rect 10870 12288 10876 12300
rect 10643 12260 10876 12288
rect 10643 12257 10655 12260
rect 10597 12251 10655 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 17681 12291 17739 12297
rect 17681 12257 17693 12291
rect 17727 12288 17739 12291
rect 17954 12288 17960 12300
rect 17727 12260 17960 12288
rect 17727 12257 17739 12260
rect 17681 12251 17739 12257
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 18233 12223 18291 12229
rect 18233 12189 18245 12223
rect 18279 12220 18291 12223
rect 22066 12220 22094 12328
rect 35342 12316 35348 12328
rect 35400 12356 35406 12368
rect 37918 12356 37924 12368
rect 35400 12328 37924 12356
rect 35400 12316 35406 12328
rect 37918 12316 37924 12328
rect 37976 12316 37982 12368
rect 38010 12316 38016 12368
rect 38068 12356 38074 12368
rect 38948 12356 38976 12396
rect 42702 12356 42708 12368
rect 38068 12328 38976 12356
rect 42663 12328 42708 12356
rect 38068 12316 38074 12328
rect 42702 12316 42708 12328
rect 42760 12316 42766 12368
rect 42794 12316 42800 12368
rect 42852 12356 42858 12368
rect 42852 12328 42897 12356
rect 42852 12316 42858 12328
rect 47210 12316 47216 12368
rect 47268 12356 47274 12368
rect 54662 12356 54668 12368
rect 47268 12328 54668 12356
rect 47268 12316 47274 12328
rect 54662 12316 54668 12328
rect 54720 12316 54726 12368
rect 30742 12248 30748 12300
rect 30800 12288 30806 12300
rect 35894 12288 35900 12300
rect 30800 12260 35900 12288
rect 30800 12248 30806 12260
rect 35894 12248 35900 12260
rect 35952 12248 35958 12300
rect 36446 12248 36452 12300
rect 36504 12288 36510 12300
rect 42058 12288 42064 12300
rect 36504 12260 42064 12288
rect 36504 12248 36510 12260
rect 42058 12248 42064 12260
rect 42116 12288 42122 12300
rect 42242 12288 42248 12300
rect 42116 12260 42248 12288
rect 42116 12248 42122 12260
rect 42242 12248 42248 12260
rect 42300 12248 42306 12300
rect 42518 12288 42524 12300
rect 42479 12260 42524 12288
rect 42518 12248 42524 12260
rect 42576 12248 42582 12300
rect 42886 12288 42892 12300
rect 42847 12260 42892 12288
rect 42886 12248 42892 12260
rect 42944 12248 42950 12300
rect 44634 12248 44640 12300
rect 44692 12288 44698 12300
rect 44818 12288 44824 12300
rect 44692 12260 44824 12288
rect 44692 12248 44698 12260
rect 44818 12248 44824 12260
rect 44876 12248 44882 12300
rect 45646 12248 45652 12300
rect 45704 12288 45710 12300
rect 46477 12291 46535 12297
rect 46477 12288 46489 12291
rect 45704 12260 46489 12288
rect 45704 12248 45710 12260
rect 46477 12257 46489 12260
rect 46523 12257 46535 12291
rect 46477 12251 46535 12257
rect 47118 12248 47124 12300
rect 47176 12288 47182 12300
rect 54772 12288 54800 12396
rect 56042 12384 56048 12436
rect 56100 12424 56106 12436
rect 56100 12396 59216 12424
rect 56100 12384 56106 12396
rect 57422 12316 57428 12368
rect 57480 12356 57486 12368
rect 59188 12356 59216 12396
rect 59538 12384 59544 12436
rect 59596 12424 59602 12436
rect 59633 12427 59691 12433
rect 59633 12424 59645 12427
rect 59596 12396 59645 12424
rect 59596 12384 59602 12396
rect 59633 12393 59645 12396
rect 59679 12393 59691 12427
rect 59633 12387 59691 12393
rect 65426 12384 65432 12436
rect 65484 12424 65490 12436
rect 65797 12427 65855 12433
rect 65797 12424 65809 12427
rect 65484 12396 65809 12424
rect 65484 12384 65490 12396
rect 65797 12393 65809 12396
rect 65843 12393 65855 12427
rect 65797 12387 65855 12393
rect 65886 12384 65892 12436
rect 65944 12424 65950 12436
rect 91002 12424 91008 12436
rect 65944 12396 91008 12424
rect 65944 12384 65950 12396
rect 91002 12384 91008 12396
rect 91060 12384 91066 12436
rect 70762 12356 70768 12368
rect 57480 12328 59124 12356
rect 59188 12328 70768 12356
rect 57480 12316 57486 12328
rect 58345 12291 58403 12297
rect 58345 12288 58357 12291
rect 47176 12260 53144 12288
rect 54772 12260 58357 12288
rect 47176 12248 47182 12260
rect 18279 12192 22094 12220
rect 18279 12189 18291 12192
rect 18233 12183 18291 12189
rect 26418 12180 26424 12232
rect 26476 12220 26482 12232
rect 30466 12220 30472 12232
rect 26476 12192 30472 12220
rect 26476 12180 26482 12192
rect 30466 12180 30472 12192
rect 30524 12220 30530 12232
rect 32030 12220 32036 12232
rect 30524 12192 32036 12220
rect 30524 12180 30530 12192
rect 32030 12180 32036 12192
rect 32088 12180 32094 12232
rect 37550 12180 37556 12232
rect 37608 12220 37614 12232
rect 42426 12220 42432 12232
rect 37608 12192 42432 12220
rect 37608 12180 37614 12192
rect 42426 12180 42432 12192
rect 42484 12180 42490 12232
rect 46198 12220 46204 12232
rect 46159 12192 46204 12220
rect 46198 12180 46204 12192
rect 46256 12180 46262 12232
rect 46658 12180 46664 12232
rect 46716 12220 46722 12232
rect 47581 12223 47639 12229
rect 47581 12220 47593 12223
rect 46716 12192 47593 12220
rect 46716 12180 46722 12192
rect 47581 12189 47593 12192
rect 47627 12189 47639 12223
rect 47581 12183 47639 12189
rect 48038 12180 48044 12232
rect 48096 12220 48102 12232
rect 50062 12220 50068 12232
rect 48096 12192 50068 12220
rect 48096 12180 48102 12192
rect 50062 12180 50068 12192
rect 50120 12180 50126 12232
rect 53116 12220 53144 12260
rect 58345 12257 58357 12260
rect 58391 12257 58403 12291
rect 58345 12251 58403 12257
rect 58437 12291 58495 12297
rect 58437 12257 58449 12291
rect 58483 12288 58495 12291
rect 58802 12288 58808 12300
rect 58483 12260 58572 12288
rect 58763 12260 58808 12288
rect 58483 12257 58495 12260
rect 58437 12251 58495 12257
rect 58544 12232 58572 12260
rect 58802 12248 58808 12260
rect 58860 12248 58866 12300
rect 59096 12297 59124 12328
rect 70762 12316 70768 12328
rect 70820 12316 70826 12368
rect 75454 12356 75460 12368
rect 72436 12328 75460 12356
rect 59081 12291 59139 12297
rect 59081 12257 59093 12291
rect 59127 12257 59139 12291
rect 59081 12251 59139 12257
rect 59173 12291 59231 12297
rect 59173 12257 59185 12291
rect 59219 12257 59231 12291
rect 59173 12251 59231 12257
rect 55858 12220 55864 12232
rect 53116 12192 55864 12220
rect 55858 12180 55864 12192
rect 55916 12180 55922 12232
rect 55950 12180 55956 12232
rect 56008 12220 56014 12232
rect 58066 12220 58072 12232
rect 56008 12192 58072 12220
rect 56008 12180 56014 12192
rect 58066 12180 58072 12192
rect 58124 12180 58130 12232
rect 58526 12180 58532 12232
rect 58584 12180 58590 12232
rect 58897 12223 58955 12229
rect 58897 12189 58909 12223
rect 58943 12220 58955 12223
rect 58986 12220 58992 12232
rect 58943 12192 58992 12220
rect 58943 12189 58955 12192
rect 58897 12183 58955 12189
rect 58986 12180 58992 12192
rect 59044 12180 59050 12232
rect 3418 12112 3424 12164
rect 3476 12152 3482 12164
rect 30650 12152 30656 12164
rect 3476 12124 30656 12152
rect 3476 12112 3482 12124
rect 30650 12112 30656 12124
rect 30708 12112 30714 12164
rect 36538 12112 36544 12164
rect 36596 12152 36602 12164
rect 41690 12152 41696 12164
rect 36596 12124 41696 12152
rect 36596 12112 36602 12124
rect 41690 12112 41696 12124
rect 41748 12112 41754 12164
rect 42702 12112 42708 12164
rect 42760 12152 42766 12164
rect 46014 12152 46020 12164
rect 42760 12124 46020 12152
rect 42760 12112 42766 12124
rect 46014 12112 46020 12124
rect 46072 12112 46078 12164
rect 47302 12112 47308 12164
rect 47360 12152 47366 12164
rect 59188 12152 59216 12251
rect 59262 12248 59268 12300
rect 59320 12288 59326 12300
rect 62209 12291 62267 12297
rect 62209 12288 62221 12291
rect 59320 12260 62221 12288
rect 59320 12248 59326 12260
rect 62209 12257 62221 12260
rect 62255 12288 62267 12291
rect 64966 12288 64972 12300
rect 62255 12260 64972 12288
rect 62255 12257 62267 12260
rect 62209 12251 62267 12257
rect 64966 12248 64972 12260
rect 65024 12248 65030 12300
rect 65886 12288 65892 12300
rect 65076 12260 65892 12288
rect 62485 12223 62543 12229
rect 62485 12189 62497 12223
rect 62531 12220 62543 12223
rect 62666 12220 62672 12232
rect 62531 12192 62672 12220
rect 62531 12189 62543 12192
rect 62485 12183 62543 12189
rect 62666 12180 62672 12192
rect 62724 12180 62730 12232
rect 63954 12180 63960 12232
rect 64012 12220 64018 12232
rect 65076 12220 65104 12260
rect 65886 12248 65892 12260
rect 65944 12248 65950 12300
rect 65981 12291 66039 12297
rect 65981 12257 65993 12291
rect 66027 12288 66039 12291
rect 72436 12288 72464 12328
rect 75454 12316 75460 12328
rect 75512 12316 75518 12368
rect 85390 12316 85396 12368
rect 85448 12356 85454 12368
rect 85666 12356 85672 12368
rect 85448 12328 85672 12356
rect 85448 12316 85454 12328
rect 85666 12316 85672 12328
rect 85724 12316 85730 12368
rect 72602 12288 72608 12300
rect 66027 12260 72464 12288
rect 72563 12260 72608 12288
rect 66027 12257 66039 12260
rect 65981 12251 66039 12257
rect 72602 12248 72608 12260
rect 72660 12248 72666 12300
rect 64012 12192 65104 12220
rect 64012 12180 64018 12192
rect 65518 12180 65524 12232
rect 65576 12220 65582 12232
rect 93670 12220 93676 12232
rect 65576 12192 93676 12220
rect 65576 12180 65582 12192
rect 93670 12180 93676 12192
rect 93728 12180 93734 12232
rect 47360 12124 59216 12152
rect 47360 12112 47366 12124
rect 59262 12112 59268 12164
rect 59320 12152 59326 12164
rect 59320 12124 70394 12152
rect 59320 12112 59326 12124
rect 4433 12087 4491 12093
rect 4433 12053 4445 12087
rect 4479 12084 4491 12087
rect 31018 12084 31024 12096
rect 4479 12056 31024 12084
rect 4479 12053 4491 12056
rect 4433 12047 4491 12053
rect 31018 12044 31024 12056
rect 31076 12044 31082 12096
rect 32490 12044 32496 12096
rect 32548 12084 32554 12096
rect 39574 12084 39580 12096
rect 32548 12056 39580 12084
rect 32548 12044 32554 12056
rect 39574 12044 39580 12056
rect 39632 12044 39638 12096
rect 40494 12044 40500 12096
rect 40552 12084 40558 12096
rect 42978 12084 42984 12096
rect 40552 12056 42984 12084
rect 40552 12044 40558 12056
rect 42978 12044 42984 12056
rect 43036 12044 43042 12096
rect 43073 12087 43131 12093
rect 43073 12053 43085 12087
rect 43119 12084 43131 12087
rect 45462 12084 45468 12096
rect 43119 12056 45468 12084
rect 43119 12053 43131 12056
rect 43073 12047 43131 12053
rect 45462 12044 45468 12056
rect 45520 12044 45526 12096
rect 45646 12044 45652 12096
rect 45704 12084 45710 12096
rect 46658 12084 46664 12096
rect 45704 12056 46664 12084
rect 45704 12044 45710 12056
rect 46658 12044 46664 12056
rect 46716 12044 46722 12096
rect 46842 12044 46848 12096
rect 46900 12084 46906 12096
rect 49050 12084 49056 12096
rect 46900 12056 49056 12084
rect 46900 12044 46906 12056
rect 49050 12044 49056 12056
rect 49108 12044 49114 12096
rect 50062 12044 50068 12096
rect 50120 12084 50126 12096
rect 50706 12084 50712 12096
rect 50120 12056 50712 12084
rect 50120 12044 50126 12056
rect 50706 12044 50712 12056
rect 50764 12044 50770 12096
rect 54662 12044 54668 12096
rect 54720 12084 54726 12096
rect 56502 12084 56508 12096
rect 54720 12056 56508 12084
rect 54720 12044 54726 12056
rect 56502 12044 56508 12056
rect 56560 12044 56566 12096
rect 57698 12084 57704 12096
rect 57659 12056 57704 12084
rect 57698 12044 57704 12056
rect 57756 12044 57762 12096
rect 58345 12087 58403 12093
rect 58345 12053 58357 12087
rect 58391 12084 58403 12087
rect 61562 12084 61568 12096
rect 58391 12056 61568 12084
rect 58391 12053 58403 12056
rect 58345 12047 58403 12053
rect 61562 12044 61568 12056
rect 61620 12044 61626 12096
rect 65334 12084 65340 12096
rect 65295 12056 65340 12084
rect 65334 12044 65340 12056
rect 65392 12044 65398 12096
rect 67358 12084 67364 12096
rect 67319 12056 67364 12084
rect 67358 12044 67364 12056
rect 67416 12044 67422 12096
rect 70366 12084 70394 12124
rect 97534 12084 97540 12096
rect 70366 12056 97540 12084
rect 97534 12044 97540 12056
rect 97592 12044 97598 12096
rect 1104 11994 98808 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 65686 11994
rect 65738 11942 65750 11994
rect 65802 11942 65814 11994
rect 65866 11942 65878 11994
rect 65930 11942 96406 11994
rect 96458 11942 96470 11994
rect 96522 11942 96534 11994
rect 96586 11942 96598 11994
rect 96650 11942 98808 11994
rect 1104 11920 98808 11942
rect 2222 11840 2228 11892
rect 2280 11880 2286 11892
rect 38654 11880 38660 11892
rect 2280 11852 38660 11880
rect 2280 11840 2286 11852
rect 38654 11840 38660 11852
rect 38712 11840 38718 11892
rect 42058 11880 42064 11892
rect 38764 11852 42064 11880
rect 10318 11812 10324 11824
rect 10279 11784 10324 11812
rect 10318 11772 10324 11784
rect 10376 11772 10382 11824
rect 17126 11812 17132 11824
rect 11808 11784 17132 11812
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 11808 11744 11836 11784
rect 17126 11772 17132 11784
rect 17184 11772 17190 11824
rect 17954 11772 17960 11824
rect 18012 11812 18018 11824
rect 18012 11784 22094 11812
rect 18012 11772 18018 11784
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 7147 11716 11836 11744
rect 12406 11716 13001 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 6914 11676 6920 11688
rect 6871 11648 6920 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 9306 11568 9312 11620
rect 9364 11608 9370 11620
rect 12406 11608 12434 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 18414 11744 18420 11756
rect 12989 11707 13047 11713
rect 13556 11716 18420 11744
rect 12805 11679 12863 11685
rect 12805 11645 12817 11679
rect 12851 11676 12863 11679
rect 13556 11676 13584 11716
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 22066 11744 22094 11784
rect 26326 11772 26332 11824
rect 26384 11812 26390 11824
rect 27154 11812 27160 11824
rect 26384 11784 27160 11812
rect 26384 11772 26390 11784
rect 27154 11772 27160 11784
rect 27212 11772 27218 11824
rect 28092 11784 38572 11812
rect 28092 11756 28120 11784
rect 28074 11744 28080 11756
rect 22066 11716 28080 11744
rect 28074 11704 28080 11716
rect 28132 11704 28138 11756
rect 28626 11744 28632 11756
rect 28587 11716 28632 11744
rect 28626 11704 28632 11716
rect 28684 11704 28690 11756
rect 36354 11704 36360 11756
rect 36412 11744 36418 11756
rect 38544 11744 38572 11784
rect 38764 11744 38792 11852
rect 42058 11840 42064 11852
rect 42116 11840 42122 11892
rect 42242 11840 42248 11892
rect 42300 11880 42306 11892
rect 46842 11880 46848 11892
rect 42300 11852 46848 11880
rect 42300 11840 42306 11852
rect 46842 11840 46848 11852
rect 46900 11840 46906 11892
rect 47762 11840 47768 11892
rect 47820 11880 47826 11892
rect 57974 11880 57980 11892
rect 47820 11852 57980 11880
rect 47820 11840 47826 11852
rect 57974 11840 57980 11852
rect 58032 11840 58038 11892
rect 58066 11840 58072 11892
rect 58124 11880 58130 11892
rect 59262 11880 59268 11892
rect 58124 11852 59268 11880
rect 58124 11840 58130 11852
rect 59262 11840 59268 11852
rect 59320 11840 59326 11892
rect 62666 11840 62672 11892
rect 62724 11880 62730 11892
rect 70118 11880 70124 11892
rect 62724 11852 70124 11880
rect 62724 11840 62730 11852
rect 70118 11840 70124 11852
rect 70176 11840 70182 11892
rect 70302 11840 70308 11892
rect 70360 11880 70366 11892
rect 79686 11880 79692 11892
rect 70360 11852 79692 11880
rect 70360 11840 70366 11852
rect 79686 11840 79692 11852
rect 79744 11840 79750 11892
rect 97629 11883 97687 11889
rect 97629 11880 97641 11883
rect 80026 11852 97641 11880
rect 38838 11772 38844 11824
rect 38896 11812 38902 11824
rect 38896 11784 39160 11812
rect 38896 11772 38902 11784
rect 39022 11744 39028 11756
rect 36412 11716 37964 11744
rect 38544 11716 38792 11744
rect 38948 11716 39028 11744
rect 36412 11704 36418 11716
rect 37936 11688 37964 11716
rect 12851 11648 13584 11676
rect 15197 11679 15255 11685
rect 12851 11645 12863 11648
rect 12805 11639 12863 11645
rect 15197 11645 15209 11679
rect 15243 11676 15255 11679
rect 15243 11648 22094 11676
rect 15243 11645 15255 11648
rect 15197 11639 15255 11645
rect 9364 11580 12434 11608
rect 9364 11568 9370 11580
rect 12526 11568 12532 11620
rect 12584 11608 12590 11620
rect 12894 11608 12900 11620
rect 12584 11580 12900 11608
rect 12584 11568 12590 11580
rect 12894 11568 12900 11580
rect 12952 11568 12958 11620
rect 17310 11608 17316 11620
rect 14844 11580 17316 11608
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 7616 11512 8401 11540
rect 7616 11500 7622 11512
rect 8389 11509 8401 11512
rect 8435 11540 8447 11543
rect 14844 11540 14872 11580
rect 17310 11568 17316 11580
rect 17368 11568 17374 11620
rect 22066 11608 22094 11648
rect 27522 11636 27528 11688
rect 27580 11676 27586 11688
rect 27801 11679 27859 11685
rect 27801 11676 27813 11679
rect 27580 11648 27813 11676
rect 27580 11636 27586 11648
rect 27801 11645 27813 11648
rect 27847 11645 27859 11679
rect 35069 11679 35127 11685
rect 35069 11676 35081 11679
rect 27801 11639 27859 11645
rect 31726 11648 35081 11676
rect 25222 11608 25228 11620
rect 22066 11580 25228 11608
rect 25222 11568 25228 11580
rect 25280 11608 25286 11620
rect 31726 11608 31754 11648
rect 35069 11645 35081 11648
rect 35115 11645 35127 11679
rect 35069 11639 35127 11645
rect 37918 11636 37924 11688
rect 37976 11676 37982 11688
rect 38197 11679 38255 11685
rect 38197 11676 38209 11679
rect 37976 11648 38209 11676
rect 37976 11636 37982 11648
rect 38197 11645 38209 11648
rect 38243 11645 38255 11679
rect 38197 11639 38255 11645
rect 25280 11580 31754 11608
rect 25280 11568 25286 11580
rect 15010 11540 15016 11552
rect 8435 11512 14872 11540
rect 14971 11512 15016 11540
rect 8435 11509 8447 11512
rect 8389 11503 8447 11509
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 28350 11540 28356 11552
rect 25556 11512 28356 11540
rect 25556 11500 25562 11512
rect 28350 11500 28356 11512
rect 28408 11540 28414 11552
rect 30374 11540 30380 11552
rect 28408 11512 30380 11540
rect 28408 11500 28414 11512
rect 30374 11500 30380 11512
rect 30432 11500 30438 11552
rect 32030 11500 32036 11552
rect 32088 11540 32094 11552
rect 34885 11543 34943 11549
rect 34885 11540 34897 11543
rect 32088 11512 34897 11540
rect 32088 11500 32094 11512
rect 34885 11509 34897 11512
rect 34931 11540 34943 11543
rect 37550 11540 37556 11552
rect 34931 11512 37556 11540
rect 34931 11509 34943 11512
rect 34885 11503 34943 11509
rect 37550 11500 37556 11512
rect 37608 11500 37614 11552
rect 37642 11500 37648 11552
rect 37700 11540 37706 11552
rect 38010 11540 38016 11552
rect 37700 11512 38016 11540
rect 37700 11500 37706 11512
rect 38010 11500 38016 11512
rect 38068 11500 38074 11552
rect 38212 11540 38240 11639
rect 38375 11636 38381 11688
rect 38433 11676 38439 11688
rect 38562 11676 38568 11688
rect 38433 11648 38478 11676
rect 38523 11648 38568 11676
rect 38433 11636 38439 11648
rect 38562 11636 38568 11648
rect 38620 11636 38626 11688
rect 38654 11636 38660 11688
rect 38712 11676 38718 11688
rect 38948 11685 38976 11716
rect 39022 11704 39028 11716
rect 39080 11704 39086 11756
rect 39132 11744 39160 11784
rect 39390 11772 39396 11824
rect 39448 11812 39454 11824
rect 45646 11812 45652 11824
rect 39448 11784 45652 11812
rect 39448 11772 39454 11784
rect 45646 11772 45652 11784
rect 45704 11772 45710 11824
rect 46198 11772 46204 11824
rect 46256 11812 46262 11824
rect 56594 11812 56600 11824
rect 46256 11784 56600 11812
rect 46256 11772 46262 11784
rect 56594 11772 56600 11784
rect 56652 11772 56658 11824
rect 58986 11772 58992 11824
rect 59044 11812 59050 11824
rect 65518 11812 65524 11824
rect 59044 11784 65524 11812
rect 59044 11772 59050 11784
rect 65518 11772 65524 11784
rect 65576 11772 65582 11824
rect 39758 11744 39764 11756
rect 39132 11716 39764 11744
rect 39758 11704 39764 11716
rect 39816 11744 39822 11756
rect 41966 11744 41972 11756
rect 39816 11716 41972 11744
rect 39816 11704 39822 11716
rect 41966 11704 41972 11716
rect 42024 11704 42030 11756
rect 42058 11704 42064 11756
rect 42116 11744 42122 11756
rect 69474 11744 69480 11756
rect 42116 11716 69480 11744
rect 42116 11704 42122 11716
rect 69474 11704 69480 11716
rect 69532 11744 69538 11756
rect 75546 11744 75552 11756
rect 69532 11716 70394 11744
rect 75507 11716 75552 11744
rect 69532 11704 69538 11716
rect 38795 11679 38853 11685
rect 38712 11648 38757 11676
rect 38712 11636 38718 11648
rect 38795 11645 38807 11679
rect 38841 11645 38853 11679
rect 38795 11639 38853 11645
rect 38933 11679 38991 11685
rect 38933 11645 38945 11679
rect 38979 11645 38991 11679
rect 62666 11676 62672 11688
rect 38933 11639 38991 11645
rect 39040 11648 62672 11676
rect 38810 11608 38838 11639
rect 38672 11580 38838 11608
rect 38672 11540 38700 11580
rect 38212 11512 38700 11540
rect 38746 11500 38752 11552
rect 38804 11540 38810 11552
rect 39040 11540 39068 11648
rect 62666 11636 62672 11648
rect 62724 11636 62730 11688
rect 70366 11676 70394 11716
rect 75546 11704 75552 11716
rect 75604 11704 75610 11756
rect 75089 11679 75147 11685
rect 75089 11676 75101 11679
rect 70366 11648 75101 11676
rect 75089 11645 75101 11648
rect 75135 11645 75147 11679
rect 75089 11639 75147 11645
rect 39117 11611 39175 11617
rect 39117 11577 39129 11611
rect 39163 11577 39175 11611
rect 39117 11571 39175 11577
rect 38804 11512 39068 11540
rect 39132 11540 39160 11571
rect 39574 11568 39580 11620
rect 39632 11608 39638 11620
rect 67266 11608 67272 11620
rect 39632 11580 67272 11608
rect 39632 11568 39638 11580
rect 67266 11568 67272 11580
rect 67324 11568 67330 11620
rect 69474 11568 69480 11620
rect 69532 11608 69538 11620
rect 80026 11608 80054 11852
rect 97629 11849 97641 11852
rect 97675 11849 97687 11883
rect 97629 11843 97687 11849
rect 85482 11812 85488 11824
rect 85443 11784 85488 11812
rect 85482 11772 85488 11784
rect 85540 11772 85546 11824
rect 91002 11812 91008 11824
rect 90963 11784 91008 11812
rect 91002 11772 91008 11784
rect 91060 11772 91066 11824
rect 85669 11679 85727 11685
rect 85669 11645 85681 11679
rect 85715 11645 85727 11679
rect 85669 11639 85727 11645
rect 85684 11608 85712 11639
rect 69532 11580 80054 11608
rect 81912 11580 85712 11608
rect 69532 11568 69538 11580
rect 67634 11540 67640 11552
rect 39132 11512 67640 11540
rect 38804 11500 38810 11512
rect 67634 11500 67640 11512
rect 67692 11500 67698 11552
rect 75454 11500 75460 11552
rect 75512 11540 75518 11552
rect 81912 11540 81940 11580
rect 75512 11512 81940 11540
rect 75512 11500 75518 11512
rect 92566 11500 92572 11552
rect 92624 11540 92630 11552
rect 96706 11540 96712 11552
rect 92624 11512 96712 11540
rect 92624 11500 92630 11512
rect 96706 11500 96712 11512
rect 96764 11500 96770 11552
rect 1104 11450 98808 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 50326 11450
rect 50378 11398 50390 11450
rect 50442 11398 50454 11450
rect 50506 11398 50518 11450
rect 50570 11398 81046 11450
rect 81098 11398 81110 11450
rect 81162 11398 81174 11450
rect 81226 11398 81238 11450
rect 81290 11398 98808 11450
rect 1104 11376 98808 11398
rect 12161 11339 12219 11345
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 12526 11336 12532 11348
rect 12207 11308 12532 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 14185 11339 14243 11345
rect 14185 11305 14197 11339
rect 14231 11336 14243 11339
rect 36538 11336 36544 11348
rect 14231 11308 36544 11336
rect 14231 11305 14243 11308
rect 14185 11299 14243 11305
rect 36538 11296 36544 11308
rect 36596 11296 36602 11348
rect 38194 11296 38200 11348
rect 38252 11336 38258 11348
rect 38252 11308 38332 11336
rect 38252 11296 38258 11308
rect 13357 11271 13415 11277
rect 13357 11268 13369 11271
rect 13188 11240 13369 11268
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 12342 11200 12348 11212
rect 6503 11172 6868 11200
rect 12303 11172 12348 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 6730 11132 6736 11144
rect 6691 11104 6736 11132
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 6840 11132 6868 11172
rect 12342 11160 12348 11172
rect 12400 11160 12406 11212
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 12584 11172 12633 11200
rect 12584 11160 12590 11172
rect 12621 11169 12633 11172
rect 12667 11169 12679 11203
rect 12621 11163 12679 11169
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13078 11209 13084 11212
rect 13025 11203 13084 11209
rect 12952 11172 12997 11200
rect 12952 11160 12958 11172
rect 13025 11169 13037 11203
rect 13071 11169 13084 11203
rect 13025 11163 13084 11169
rect 13078 11160 13084 11163
rect 13136 11160 13142 11212
rect 13188 11209 13216 11240
rect 13357 11237 13369 11240
rect 13403 11268 13415 11271
rect 26786 11268 26792 11280
rect 13403 11240 26792 11268
rect 13403 11237 13415 11240
rect 13357 11231 13415 11237
rect 26786 11228 26792 11240
rect 26844 11228 26850 11280
rect 28350 11268 28356 11280
rect 28311 11240 28356 11268
rect 28350 11228 28356 11240
rect 28408 11228 28414 11280
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 21453 11203 21511 11209
rect 21453 11169 21465 11203
rect 21499 11200 21511 11203
rect 21726 11200 21732 11212
rect 21499 11172 21732 11200
rect 21499 11169 21511 11172
rect 21453 11163 21511 11169
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 25409 11203 25467 11209
rect 25409 11169 25421 11203
rect 25455 11200 25467 11203
rect 26326 11200 26332 11212
rect 25455 11172 26332 11200
rect 25455 11169 25467 11172
rect 25409 11163 25467 11169
rect 26326 11160 26332 11172
rect 26384 11160 26390 11212
rect 26605 11203 26663 11209
rect 26605 11169 26617 11203
rect 26651 11200 26663 11203
rect 26651 11172 27108 11200
rect 26651 11169 26663 11172
rect 26605 11163 26663 11169
rect 6914 11132 6920 11144
rect 6840 11104 6920 11132
rect 6914 11092 6920 11104
rect 6972 11132 6978 11144
rect 7650 11132 7656 11144
rect 6972 11104 7656 11132
rect 6972 11092 6978 11104
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8159 11104 12664 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 12636 11064 12664 11104
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 12860 11104 14197 11132
rect 12860 11092 12866 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 26418 11092 26424 11144
rect 26476 11132 26482 11144
rect 26697 11135 26755 11141
rect 26697 11132 26709 11135
rect 26476 11104 26709 11132
rect 26476 11092 26482 11104
rect 26697 11101 26709 11104
rect 26743 11101 26755 11135
rect 26697 11095 26755 11101
rect 26878 11092 26884 11144
rect 26936 11132 26942 11144
rect 26973 11135 27031 11141
rect 26973 11132 26985 11135
rect 26936 11104 26985 11132
rect 26936 11092 26942 11104
rect 26973 11101 26985 11104
rect 27019 11101 27031 11135
rect 27080 11132 27108 11172
rect 27246 11160 27252 11212
rect 27304 11200 27310 11212
rect 36446 11200 36452 11212
rect 27304 11172 36452 11200
rect 27304 11160 27310 11172
rect 36446 11160 36452 11172
rect 36504 11160 36510 11212
rect 37274 11160 37280 11212
rect 37332 11200 37338 11212
rect 38197 11203 38255 11209
rect 38197 11200 38209 11203
rect 37332 11172 38209 11200
rect 37332 11160 37338 11172
rect 38197 11169 38209 11172
rect 38243 11169 38255 11203
rect 38304 11200 38332 11308
rect 38378 11296 38384 11348
rect 38436 11296 38442 11348
rect 38562 11296 38568 11348
rect 38620 11336 38626 11348
rect 38620 11308 38700 11336
rect 38620 11296 38626 11308
rect 38396 11268 38424 11296
rect 38672 11268 38700 11308
rect 41966 11296 41972 11348
rect 42024 11336 42030 11348
rect 55858 11336 55864 11348
rect 42024 11308 55864 11336
rect 42024 11296 42030 11308
rect 55858 11296 55864 11308
rect 55916 11296 55922 11348
rect 60366 11296 60372 11348
rect 60424 11336 60430 11348
rect 60424 11308 67220 11336
rect 60424 11296 60430 11308
rect 38396 11240 38608 11268
rect 38672 11240 38792 11268
rect 38580 11212 38608 11240
rect 38381 11203 38439 11209
rect 38381 11200 38393 11203
rect 38304 11172 38393 11200
rect 38197 11163 38255 11169
rect 38381 11169 38393 11172
rect 38427 11169 38439 11203
rect 38381 11163 38439 11169
rect 38562 11160 38568 11212
rect 38620 11200 38626 11212
rect 38764 11200 38792 11240
rect 38838 11228 38844 11280
rect 38896 11268 38902 11280
rect 38896 11240 39160 11268
rect 38896 11228 38902 11240
rect 39132 11209 39160 11240
rect 39224 11240 42932 11268
rect 38933 11203 38991 11209
rect 38933 11200 38945 11203
rect 38620 11172 38713 11200
rect 38764 11172 38945 11200
rect 38620 11160 38626 11172
rect 38933 11169 38945 11172
rect 38979 11169 38991 11203
rect 38933 11163 38991 11169
rect 39117 11203 39175 11209
rect 39117 11169 39129 11203
rect 39163 11169 39175 11203
rect 39117 11163 39175 11169
rect 37737 11135 37795 11141
rect 27080 11104 31754 11132
rect 26973 11095 27031 11101
rect 26605 11067 26663 11073
rect 26605 11064 26617 11067
rect 7760 11036 7972 11064
rect 4890 10956 4896 11008
rect 4948 10996 4954 11008
rect 7760 10996 7788 11036
rect 4948 10968 7788 10996
rect 7944 10996 7972 11036
rect 11992 11036 12434 11064
rect 12636 11036 26617 11064
rect 11992 10996 12020 11036
rect 7944 10968 12020 10996
rect 12406 11008 12434 11036
rect 26605 11033 26617 11036
rect 26651 11033 26663 11067
rect 31726 11064 31754 11104
rect 37737 11101 37749 11135
rect 37783 11132 37795 11135
rect 39224 11132 39252 11240
rect 41598 11160 41604 11212
rect 41656 11200 41662 11212
rect 42613 11203 42671 11209
rect 42613 11200 42625 11203
rect 41656 11172 42625 11200
rect 41656 11160 41662 11172
rect 42613 11169 42625 11172
rect 42659 11169 42671 11203
rect 42904 11200 42932 11240
rect 42978 11228 42984 11280
rect 43036 11268 43042 11280
rect 67192 11277 67220 11308
rect 67450 11296 67456 11348
rect 67508 11336 67514 11348
rect 69017 11339 69075 11345
rect 69017 11336 69029 11339
rect 67508 11308 69029 11336
rect 67508 11296 67514 11308
rect 69017 11305 69029 11308
rect 69063 11305 69075 11339
rect 69017 11299 69075 11305
rect 69290 11296 69296 11348
rect 69348 11336 69354 11348
rect 69348 11308 69520 11336
rect 69348 11296 69354 11308
rect 67177 11271 67235 11277
rect 43036 11240 65196 11268
rect 43036 11228 43042 11240
rect 42904 11172 55628 11200
rect 42613 11163 42671 11169
rect 55490 11132 55496 11144
rect 37783 11104 39252 11132
rect 39316 11104 55496 11132
rect 37783 11101 37795 11104
rect 37737 11095 37795 11101
rect 39316 11064 39344 11104
rect 55490 11092 55496 11104
rect 55548 11092 55554 11144
rect 55600 11132 55628 11172
rect 55858 11160 55864 11212
rect 55916 11200 55922 11212
rect 62942 11200 62948 11212
rect 55916 11172 62948 11200
rect 55916 11160 55922 11172
rect 62942 11160 62948 11172
rect 63000 11160 63006 11212
rect 65168 11200 65196 11240
rect 67177 11237 67189 11271
rect 67223 11237 67235 11271
rect 67177 11231 67235 11237
rect 67818 11228 67824 11280
rect 67876 11268 67882 11280
rect 67913 11271 67971 11277
rect 67913 11268 67925 11271
rect 67876 11240 67925 11268
rect 67876 11228 67882 11240
rect 67913 11237 67925 11240
rect 67959 11237 67971 11271
rect 69385 11271 69443 11277
rect 69385 11268 69397 11271
rect 67913 11231 67971 11237
rect 68020 11240 69397 11268
rect 68020 11200 68048 11240
rect 69385 11237 69397 11240
rect 69431 11237 69443 11271
rect 69492 11268 69520 11308
rect 69842 11296 69848 11348
rect 69900 11336 69906 11348
rect 95973 11339 96031 11345
rect 95973 11336 95985 11339
rect 69900 11308 95985 11336
rect 69900 11296 69906 11308
rect 95973 11305 95985 11308
rect 96019 11305 96031 11339
rect 97534 11336 97540 11348
rect 97495 11308 97540 11336
rect 95973 11299 96031 11305
rect 97534 11296 97540 11308
rect 97592 11296 97598 11348
rect 69492 11240 97028 11268
rect 69385 11231 69443 11237
rect 65168 11172 68048 11200
rect 69017 11203 69075 11209
rect 69017 11169 69029 11203
rect 69063 11200 69075 11203
rect 69109 11203 69167 11209
rect 69109 11200 69121 11203
rect 69063 11172 69121 11200
rect 69063 11169 69075 11172
rect 69017 11163 69075 11169
rect 69109 11169 69121 11172
rect 69155 11169 69167 11203
rect 69109 11163 69167 11169
rect 69216 11172 70394 11200
rect 58066 11132 58072 11144
rect 55600 11104 58072 11132
rect 58066 11092 58072 11104
rect 58124 11092 58130 11144
rect 59722 11092 59728 11144
rect 59780 11132 59786 11144
rect 69216 11132 69244 11172
rect 59780 11104 69244 11132
rect 70366 11132 70394 11172
rect 72326 11160 72332 11212
rect 72384 11200 72390 11212
rect 73890 11200 73896 11212
rect 72384 11172 73896 11200
rect 72384 11160 72390 11172
rect 73890 11160 73896 11172
rect 73948 11160 73954 11212
rect 79778 11160 79784 11212
rect 79836 11200 79842 11212
rect 82630 11200 82636 11212
rect 79836 11172 82636 11200
rect 79836 11160 79842 11172
rect 82630 11160 82636 11172
rect 82688 11160 82694 11212
rect 95973 11203 96031 11209
rect 95973 11169 95985 11203
rect 96019 11200 96031 11203
rect 96341 11203 96399 11209
rect 96341 11200 96353 11203
rect 96019 11172 96353 11200
rect 96019 11169 96031 11172
rect 95973 11163 96031 11169
rect 96341 11169 96353 11172
rect 96387 11169 96399 11203
rect 96706 11200 96712 11212
rect 96667 11172 96712 11200
rect 96341 11163 96399 11169
rect 96706 11160 96712 11172
rect 96764 11160 96770 11212
rect 97000 11209 97028 11240
rect 96985 11203 97043 11209
rect 96985 11169 96997 11203
rect 97031 11169 97043 11203
rect 96985 11163 97043 11169
rect 97077 11203 97135 11209
rect 97077 11169 97089 11203
rect 97123 11169 97135 11203
rect 97077 11163 97135 11169
rect 96157 11135 96215 11141
rect 96157 11132 96169 11135
rect 70366 11104 96169 11132
rect 59780 11092 59786 11104
rect 96157 11101 96169 11104
rect 96203 11132 96215 11135
rect 96525 11135 96583 11141
rect 96525 11132 96537 11135
rect 96203 11104 96537 11132
rect 96203 11101 96215 11104
rect 96157 11095 96215 11101
rect 96525 11101 96537 11104
rect 96571 11101 96583 11135
rect 96525 11095 96583 11101
rect 31726 11036 39344 11064
rect 39393 11067 39451 11073
rect 26605 11027 26663 11033
rect 39393 11033 39405 11067
rect 39439 11064 39451 11067
rect 86494 11064 86500 11076
rect 39439 11036 86500 11064
rect 39439 11033 39451 11036
rect 39393 11027 39451 11033
rect 86494 11024 86500 11036
rect 86552 11024 86558 11076
rect 92658 11024 92664 11076
rect 92716 11064 92722 11076
rect 97092 11064 97120 11163
rect 92716 11036 97120 11064
rect 92716 11024 92722 11036
rect 12406 10968 12440 11008
rect 4948 10956 4954 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 25222 10996 25228 11008
rect 12584 10968 12629 10996
rect 25183 10968 25228 10996
rect 12584 10956 12590 10968
rect 25222 10956 25228 10968
rect 25280 10956 25286 11008
rect 26234 10956 26240 11008
rect 26292 10996 26298 11008
rect 28626 10996 28632 11008
rect 26292 10968 28632 10996
rect 26292 10956 26298 10968
rect 28626 10956 28632 10968
rect 28684 10956 28690 11008
rect 35802 10956 35808 11008
rect 35860 10996 35866 11008
rect 61470 10996 61476 11008
rect 35860 10968 61476 10996
rect 35860 10956 35866 10968
rect 61470 10956 61476 10968
rect 61528 10956 61534 11008
rect 61562 10956 61568 11008
rect 61620 10996 61626 11008
rect 62850 10996 62856 11008
rect 61620 10968 62856 10996
rect 61620 10956 61626 10968
rect 62850 10956 62856 10968
rect 62908 10956 62914 11008
rect 64322 10956 64328 11008
rect 64380 10996 64386 11008
rect 83090 10996 83096 11008
rect 64380 10968 83096 10996
rect 64380 10956 64386 10968
rect 83090 10956 83096 10968
rect 83148 10956 83154 11008
rect 1104 10906 98808 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 65686 10906
rect 65738 10854 65750 10906
rect 65802 10854 65814 10906
rect 65866 10854 65878 10906
rect 65930 10854 96406 10906
rect 96458 10854 96470 10906
rect 96522 10854 96534 10906
rect 96586 10854 96598 10906
rect 96650 10854 98808 10906
rect 1104 10832 98808 10854
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 28442 10792 28448 10804
rect 12492 10764 28448 10792
rect 12492 10752 12498 10764
rect 28442 10752 28448 10764
rect 28500 10752 28506 10804
rect 28626 10752 28632 10804
rect 28684 10792 28690 10804
rect 42886 10792 42892 10804
rect 28684 10764 42892 10792
rect 28684 10752 28690 10764
rect 42886 10752 42892 10764
rect 42944 10752 42950 10804
rect 44634 10752 44640 10804
rect 44692 10792 44698 10804
rect 44821 10795 44879 10801
rect 44821 10792 44833 10795
rect 44692 10764 44833 10792
rect 44692 10752 44698 10764
rect 44821 10761 44833 10764
rect 44867 10761 44879 10795
rect 44821 10755 44879 10761
rect 45094 10752 45100 10804
rect 45152 10792 45158 10804
rect 46382 10792 46388 10804
rect 45152 10764 46388 10792
rect 45152 10752 45158 10764
rect 46382 10752 46388 10764
rect 46440 10752 46446 10804
rect 57974 10752 57980 10804
rect 58032 10792 58038 10804
rect 91554 10792 91560 10804
rect 58032 10764 91560 10792
rect 58032 10752 58038 10764
rect 91554 10752 91560 10764
rect 91612 10752 91618 10804
rect 12250 10684 12256 10736
rect 12308 10724 12314 10736
rect 32766 10724 32772 10736
rect 12308 10696 32772 10724
rect 12308 10684 12314 10696
rect 32766 10684 32772 10696
rect 32824 10684 32830 10736
rect 33244 10696 33640 10724
rect 25958 10616 25964 10668
rect 26016 10656 26022 10668
rect 33244 10656 33272 10696
rect 26016 10628 33272 10656
rect 33612 10656 33640 10696
rect 36538 10684 36544 10736
rect 36596 10724 36602 10736
rect 44358 10724 44364 10736
rect 36596 10696 44364 10724
rect 36596 10684 36602 10696
rect 44358 10684 44364 10696
rect 44416 10684 44422 10736
rect 45370 10684 45376 10736
rect 45428 10724 45434 10736
rect 49418 10724 49424 10736
rect 45428 10696 49424 10724
rect 45428 10684 45434 10696
rect 49418 10684 49424 10696
rect 49476 10684 49482 10736
rect 51718 10684 51724 10736
rect 51776 10724 51782 10736
rect 61654 10724 61660 10736
rect 51776 10696 61660 10724
rect 51776 10684 51782 10696
rect 61654 10684 61660 10696
rect 61712 10684 61718 10736
rect 67266 10724 67272 10736
rect 67227 10696 67272 10724
rect 67266 10684 67272 10696
rect 67324 10684 67330 10736
rect 67376 10696 68968 10724
rect 41138 10656 41144 10668
rect 33612 10628 41144 10656
rect 26016 10616 26022 10628
rect 41138 10616 41144 10628
rect 41196 10616 41202 10668
rect 44375 10656 44403 10684
rect 44545 10659 44603 10665
rect 44545 10656 44557 10659
rect 44375 10628 44557 10656
rect 44545 10625 44557 10628
rect 44591 10625 44603 10659
rect 46290 10656 46296 10668
rect 44545 10619 44603 10625
rect 44652 10628 46296 10656
rect 20070 10548 20076 10600
rect 20128 10588 20134 10600
rect 27246 10588 27252 10600
rect 20128 10560 27252 10588
rect 20128 10548 20134 10560
rect 27246 10548 27252 10560
rect 27304 10548 27310 10600
rect 28353 10591 28411 10597
rect 28353 10557 28365 10591
rect 28399 10588 28411 10591
rect 33226 10588 33232 10600
rect 28399 10560 33232 10588
rect 28399 10557 28411 10560
rect 28353 10551 28411 10557
rect 33226 10548 33232 10560
rect 33284 10548 33290 10600
rect 33410 10548 33416 10600
rect 33468 10588 33474 10600
rect 36446 10588 36452 10600
rect 33468 10560 36452 10588
rect 33468 10548 33474 10560
rect 36446 10548 36452 10560
rect 36504 10548 36510 10600
rect 41782 10588 41788 10600
rect 36556 10560 41788 10588
rect 5442 10480 5448 10532
rect 5500 10520 5506 10532
rect 36556 10520 36584 10560
rect 41782 10548 41788 10560
rect 41840 10548 41846 10600
rect 44174 10588 44180 10600
rect 44135 10560 44180 10588
rect 44174 10548 44180 10560
rect 44232 10548 44238 10600
rect 44266 10548 44272 10600
rect 44324 10597 44330 10600
rect 44324 10591 44383 10597
rect 44324 10557 44337 10591
rect 44371 10557 44383 10591
rect 44324 10551 44383 10557
rect 44453 10591 44511 10597
rect 44453 10557 44465 10591
rect 44499 10588 44511 10591
rect 44652 10588 44680 10628
rect 46290 10616 46296 10628
rect 46348 10616 46354 10668
rect 46566 10616 46572 10668
rect 46624 10656 46630 10668
rect 61470 10656 61476 10668
rect 46624 10628 61476 10656
rect 46624 10616 46630 10628
rect 61470 10616 61476 10628
rect 61528 10616 61534 10668
rect 66349 10659 66407 10665
rect 66349 10656 66361 10659
rect 61580 10628 66361 10656
rect 44499 10560 44680 10588
rect 44729 10591 44787 10597
rect 44499 10557 44511 10560
rect 44453 10551 44511 10557
rect 44729 10557 44741 10591
rect 44775 10588 44787 10591
rect 45186 10588 45192 10600
rect 44775 10560 45192 10588
rect 44775 10557 44787 10560
rect 44729 10551 44787 10557
rect 44324 10548 44330 10551
rect 45186 10548 45192 10560
rect 45244 10548 45250 10600
rect 47762 10548 47768 10600
rect 47820 10588 47826 10600
rect 51718 10588 51724 10600
rect 47820 10560 51724 10588
rect 47820 10548 47826 10560
rect 51718 10548 51724 10560
rect 51776 10548 51782 10600
rect 51902 10548 51908 10600
rect 51960 10588 51966 10600
rect 58158 10588 58164 10600
rect 51960 10560 58164 10588
rect 51960 10548 51966 10560
rect 58158 10548 58164 10560
rect 58216 10548 58222 10600
rect 5500 10492 36584 10520
rect 5500 10480 5506 10492
rect 37918 10480 37924 10532
rect 37976 10520 37982 10532
rect 39666 10520 39672 10532
rect 37976 10492 39672 10520
rect 37976 10480 37982 10492
rect 39666 10480 39672 10492
rect 39724 10480 39730 10532
rect 41386 10492 51074 10520
rect 12526 10412 12532 10464
rect 12584 10452 12590 10464
rect 41386 10452 41414 10492
rect 12584 10424 41414 10452
rect 12584 10412 12590 10424
rect 41690 10412 41696 10464
rect 41748 10452 41754 10464
rect 50614 10452 50620 10464
rect 41748 10424 50620 10452
rect 41748 10412 41754 10424
rect 50614 10412 50620 10424
rect 50672 10412 50678 10464
rect 51046 10452 51074 10492
rect 57330 10480 57336 10532
rect 57388 10520 57394 10532
rect 61580 10520 61608 10628
rect 66349 10625 66361 10628
rect 66395 10625 66407 10659
rect 66349 10619 66407 10625
rect 61654 10548 61660 10600
rect 61712 10588 61718 10600
rect 61838 10588 61844 10600
rect 61712 10560 61844 10588
rect 61712 10548 61718 10560
rect 61838 10548 61844 10560
rect 61896 10548 61902 10600
rect 62117 10591 62175 10597
rect 62117 10588 62129 10591
rect 61948 10560 62129 10588
rect 61948 10520 61976 10560
rect 62117 10557 62129 10560
rect 62163 10557 62175 10591
rect 62117 10551 62175 10557
rect 64966 10548 64972 10600
rect 65024 10588 65030 10600
rect 65337 10591 65395 10597
rect 65337 10588 65349 10591
rect 65024 10560 65349 10588
rect 65024 10548 65030 10560
rect 65337 10557 65349 10560
rect 65383 10588 65395 10591
rect 67376 10588 67404 10696
rect 68940 10656 68968 10696
rect 69106 10684 69112 10736
rect 69164 10724 69170 10736
rect 87782 10724 87788 10736
rect 69164 10696 87788 10724
rect 69164 10684 69170 10696
rect 87782 10684 87788 10696
rect 87840 10684 87846 10736
rect 85942 10656 85948 10668
rect 65383 10560 67404 10588
rect 67606 10628 68876 10656
rect 68940 10628 85948 10656
rect 65383 10557 65395 10560
rect 65337 10551 65395 10557
rect 65242 10520 65248 10532
rect 57388 10492 61608 10520
rect 61672 10492 61976 10520
rect 62776 10492 63356 10520
rect 65203 10492 65248 10520
rect 57388 10480 57394 10492
rect 61672 10461 61700 10492
rect 61657 10455 61715 10461
rect 61657 10452 61669 10455
rect 51046 10424 61669 10452
rect 61657 10421 61669 10424
rect 61703 10421 61715 10455
rect 61657 10415 61715 10421
rect 62114 10412 62120 10464
rect 62172 10452 62178 10464
rect 62776 10452 62804 10492
rect 62172 10424 62804 10452
rect 62172 10412 62178 10424
rect 62942 10412 62948 10464
rect 63000 10452 63006 10464
rect 63218 10452 63224 10464
rect 63000 10424 63224 10452
rect 63000 10412 63006 10424
rect 63218 10412 63224 10424
rect 63276 10412 63282 10464
rect 63328 10452 63356 10492
rect 65242 10480 65248 10492
rect 65300 10480 65306 10532
rect 66349 10523 66407 10529
rect 66349 10489 66361 10523
rect 66395 10520 66407 10523
rect 67606 10520 67634 10628
rect 68646 10548 68652 10600
rect 68704 10588 68710 10600
rect 68741 10591 68799 10597
rect 68741 10588 68753 10591
rect 68704 10560 68753 10588
rect 68704 10548 68710 10560
rect 68741 10557 68753 10560
rect 68787 10557 68799 10591
rect 68848 10588 68876 10628
rect 85942 10616 85948 10628
rect 86000 10616 86006 10668
rect 75086 10588 75092 10600
rect 68848 10560 75092 10588
rect 68741 10551 68799 10557
rect 75086 10548 75092 10560
rect 75144 10548 75150 10600
rect 77938 10588 77944 10600
rect 75196 10560 77944 10588
rect 66395 10492 67634 10520
rect 66395 10489 66407 10492
rect 66349 10483 66407 10489
rect 71498 10480 71504 10532
rect 71556 10520 71562 10532
rect 75196 10520 75224 10560
rect 77938 10548 77944 10560
rect 77996 10548 78002 10600
rect 82630 10548 82636 10600
rect 82688 10588 82694 10600
rect 91005 10591 91063 10597
rect 91005 10588 91017 10591
rect 82688 10560 91017 10588
rect 82688 10548 82694 10560
rect 91005 10557 91017 10560
rect 91051 10557 91063 10591
rect 91005 10551 91063 10557
rect 71556 10492 75224 10520
rect 71556 10480 71562 10492
rect 75270 10480 75276 10532
rect 75328 10520 75334 10532
rect 91281 10523 91339 10529
rect 91281 10520 91293 10523
rect 75328 10492 91293 10520
rect 75328 10480 75334 10492
rect 91281 10489 91293 10492
rect 91327 10489 91339 10523
rect 91281 10483 91339 10489
rect 68278 10452 68284 10464
rect 63328 10424 68284 10452
rect 68278 10412 68284 10424
rect 68336 10412 68342 10464
rect 75178 10412 75184 10464
rect 75236 10452 75242 10464
rect 96062 10452 96068 10464
rect 75236 10424 96068 10452
rect 75236 10412 75242 10424
rect 96062 10412 96068 10424
rect 96120 10412 96126 10464
rect 1104 10362 98808 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 50326 10362
rect 50378 10310 50390 10362
rect 50442 10310 50454 10362
rect 50506 10310 50518 10362
rect 50570 10310 81046 10362
rect 81098 10310 81110 10362
rect 81162 10310 81174 10362
rect 81226 10310 81238 10362
rect 81290 10310 98808 10362
rect 1104 10288 98808 10310
rect 9766 10248 9772 10260
rect 6656 10220 9772 10248
rect 4890 10180 4896 10192
rect 4851 10152 4896 10180
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 6656 10121 6684 10220
rect 9766 10208 9772 10220
rect 9824 10248 9830 10260
rect 10870 10248 10876 10260
rect 9824 10220 10876 10248
rect 9824 10208 9830 10220
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 25774 10208 25780 10260
rect 25832 10248 25838 10260
rect 26234 10248 26240 10260
rect 25832 10220 26240 10248
rect 25832 10208 25838 10220
rect 26234 10208 26240 10220
rect 26292 10208 26298 10260
rect 26326 10208 26332 10260
rect 26384 10208 26390 10260
rect 27246 10248 27252 10260
rect 27207 10220 27252 10248
rect 27246 10208 27252 10220
rect 27304 10208 27310 10260
rect 28074 10248 28080 10260
rect 28035 10220 28080 10248
rect 28074 10208 28080 10220
rect 28132 10208 28138 10260
rect 29917 10251 29975 10257
rect 29917 10248 29929 10251
rect 28368 10220 29929 10248
rect 26344 10180 26372 10208
rect 28368 10180 28396 10220
rect 29917 10217 29929 10220
rect 29963 10217 29975 10251
rect 29917 10211 29975 10217
rect 32766 10208 32772 10260
rect 32824 10248 32830 10260
rect 46198 10248 46204 10260
rect 32824 10220 46204 10248
rect 32824 10208 32830 10220
rect 46198 10208 46204 10220
rect 46256 10208 46262 10260
rect 46474 10208 46480 10260
rect 46532 10248 46538 10260
rect 50706 10248 50712 10260
rect 46532 10220 50712 10248
rect 46532 10208 46538 10220
rect 50706 10208 50712 10220
rect 50764 10248 50770 10260
rect 57425 10251 57483 10257
rect 57425 10248 57437 10251
rect 50764 10220 57437 10248
rect 50764 10208 50770 10220
rect 57425 10217 57437 10220
rect 57471 10217 57483 10251
rect 57425 10211 57483 10217
rect 57517 10251 57575 10257
rect 57517 10217 57529 10251
rect 57563 10248 57575 10251
rect 65242 10248 65248 10260
rect 57563 10220 65248 10248
rect 57563 10217 57575 10220
rect 57517 10211 57575 10217
rect 65242 10208 65248 10220
rect 65300 10208 65306 10260
rect 67358 10208 67364 10260
rect 67416 10248 67422 10260
rect 75178 10248 75184 10260
rect 67416 10220 75184 10248
rect 67416 10208 67422 10220
rect 75178 10208 75184 10220
rect 75236 10208 75242 10260
rect 36538 10180 36544 10192
rect 22066 10152 26280 10180
rect 26344 10152 28396 10180
rect 28460 10152 36544 10180
rect 4341 10115 4399 10121
rect 4341 10081 4353 10115
rect 4387 10112 4399 10115
rect 6641 10115 6699 10121
rect 4387 10084 5672 10112
rect 4387 10081 4399 10084
rect 4341 10075 4399 10081
rect 5644 10044 5672 10084
rect 6641 10081 6653 10115
rect 6687 10081 6699 10115
rect 6641 10075 6699 10081
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10112 7343 10115
rect 18506 10112 18512 10124
rect 7331 10084 18512 10112
rect 7331 10081 7343 10084
rect 7285 10075 7343 10081
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 18782 10072 18788 10124
rect 18840 10112 18846 10124
rect 20070 10112 20076 10124
rect 18840 10084 20076 10112
rect 18840 10072 18846 10084
rect 20070 10072 20076 10084
rect 20128 10072 20134 10124
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 21174 10112 21180 10124
rect 20864 10084 21180 10112
rect 20864 10072 20870 10084
rect 21174 10072 21180 10084
rect 21232 10112 21238 10124
rect 22066 10112 22094 10152
rect 21232 10084 22094 10112
rect 21232 10072 21238 10084
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 26125 10115 26183 10121
rect 26125 10112 26137 10115
rect 23440 10084 26137 10112
rect 23440 10072 23446 10084
rect 26125 10081 26137 10084
rect 26171 10081 26183 10115
rect 26252 10112 26280 10152
rect 27062 10112 27068 10124
rect 26252 10084 27068 10112
rect 26125 10075 26183 10081
rect 27062 10072 27068 10084
rect 27120 10072 27126 10124
rect 27982 10112 27988 10124
rect 27943 10084 27988 10112
rect 27982 10072 27988 10084
rect 28040 10072 28046 10124
rect 28460 10112 28488 10152
rect 36538 10140 36544 10152
rect 36596 10140 36602 10192
rect 39206 10140 39212 10192
rect 39264 10180 39270 10192
rect 42426 10180 42432 10192
rect 39264 10152 42432 10180
rect 39264 10140 39270 10152
rect 42426 10140 42432 10152
rect 42484 10140 42490 10192
rect 42794 10140 42800 10192
rect 42852 10180 42858 10192
rect 45370 10180 45376 10192
rect 42852 10152 45376 10180
rect 42852 10140 42858 10152
rect 45370 10140 45376 10152
rect 45428 10140 45434 10192
rect 46290 10140 46296 10192
rect 46348 10180 46354 10192
rect 86770 10180 86776 10192
rect 46348 10152 86776 10180
rect 46348 10140 46354 10152
rect 86770 10140 86776 10152
rect 86828 10140 86834 10192
rect 28092 10084 28488 10112
rect 29917 10115 29975 10121
rect 9122 10044 9128 10056
rect 5644 10016 9128 10044
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 10502 10044 10508 10056
rect 9447 10016 10508 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 10502 10004 10508 10016
rect 10560 10044 10566 10056
rect 10873 10047 10931 10053
rect 10873 10044 10885 10047
rect 10560 10016 10885 10044
rect 10560 10004 10566 10016
rect 10873 10013 10885 10016
rect 10919 10013 10931 10047
rect 11146 10044 11152 10056
rect 11059 10016 11152 10044
rect 10873 10007 10931 10013
rect 11146 10004 11152 10016
rect 11204 10044 11210 10056
rect 15010 10044 15016 10056
rect 11204 10016 15016 10044
rect 11204 10004 11210 10016
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 18598 10004 18604 10056
rect 18656 10044 18662 10056
rect 18656 10016 20760 10044
rect 18656 10004 18662 10016
rect 6178 9936 6184 9988
rect 6236 9976 6242 9988
rect 7650 9976 7656 9988
rect 6236 9948 7656 9976
rect 6236 9936 6242 9948
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 18690 9936 18696 9988
rect 18748 9976 18754 9988
rect 20622 9976 20628 9988
rect 18748 9948 20628 9976
rect 18748 9936 18754 9948
rect 20622 9936 20628 9948
rect 20680 9936 20686 9988
rect 20732 9976 20760 10016
rect 24854 10004 24860 10056
rect 24912 10044 24918 10056
rect 25130 10044 25136 10056
rect 24912 10016 25136 10044
rect 24912 10004 24918 10016
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 25866 10044 25872 10056
rect 25827 10016 25872 10044
rect 25866 10004 25872 10016
rect 25924 10004 25930 10056
rect 26970 10004 26976 10056
rect 27028 10044 27034 10056
rect 28092 10044 28120 10084
rect 29917 10081 29929 10115
rect 29963 10112 29975 10115
rect 29963 10084 33640 10112
rect 29963 10081 29975 10084
rect 29917 10075 29975 10081
rect 27028 10016 28120 10044
rect 27028 10004 27034 10016
rect 28442 10004 28448 10056
rect 28500 10044 28506 10056
rect 33410 10044 33416 10056
rect 28500 10016 33416 10044
rect 28500 10004 28506 10016
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 33612 10044 33640 10084
rect 33962 10072 33968 10124
rect 34020 10112 34026 10124
rect 57517 10115 57575 10121
rect 57517 10112 57529 10115
rect 34020 10084 57529 10112
rect 34020 10072 34026 10084
rect 57517 10081 57529 10084
rect 57563 10112 57575 10115
rect 57701 10115 57759 10121
rect 57701 10112 57713 10115
rect 57563 10084 57713 10112
rect 57563 10081 57575 10084
rect 57517 10075 57575 10081
rect 57701 10081 57713 10084
rect 57747 10081 57759 10115
rect 57701 10075 57759 10081
rect 62666 10072 62672 10124
rect 62724 10112 62730 10124
rect 63402 10112 63408 10124
rect 62724 10084 63408 10112
rect 62724 10072 62730 10084
rect 63402 10072 63408 10084
rect 63460 10072 63466 10124
rect 63494 10072 63500 10124
rect 63552 10112 63558 10124
rect 63552 10084 71820 10112
rect 63552 10072 63558 10084
rect 37918 10044 37924 10056
rect 33612 10016 37924 10044
rect 37918 10004 37924 10016
rect 37976 10004 37982 10056
rect 38105 10047 38163 10053
rect 38105 10013 38117 10047
rect 38151 10013 38163 10047
rect 38105 10007 38163 10013
rect 38381 10047 38439 10053
rect 38381 10013 38393 10047
rect 38427 10044 38439 10047
rect 52730 10044 52736 10056
rect 38427 10016 52736 10044
rect 38427 10013 38439 10016
rect 38381 10007 38439 10013
rect 30374 9976 30380 9988
rect 20732 9948 25912 9976
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9769 9911 9827 9917
rect 9769 9908 9781 9911
rect 9732 9880 9781 9908
rect 9732 9868 9738 9880
rect 9769 9877 9781 9880
rect 9815 9908 9827 9911
rect 25774 9908 25780 9920
rect 9815 9880 25780 9908
rect 9815 9877 9827 9880
rect 9769 9871 9827 9877
rect 25774 9868 25780 9880
rect 25832 9868 25838 9920
rect 25884 9908 25912 9948
rect 26988 9948 30380 9976
rect 26988 9908 27016 9948
rect 30374 9936 30380 9948
rect 30432 9936 30438 9988
rect 31202 9936 31208 9988
rect 31260 9976 31266 9988
rect 31260 9948 36584 9976
rect 31260 9936 31266 9948
rect 25884 9880 27016 9908
rect 27062 9868 27068 9920
rect 27120 9908 27126 9920
rect 33962 9908 33968 9920
rect 27120 9880 33968 9908
rect 27120 9868 27126 9880
rect 33962 9868 33968 9880
rect 34020 9868 34026 9920
rect 36556 9908 36584 9948
rect 37550 9936 37556 9988
rect 37608 9976 37614 9988
rect 38120 9976 38148 10007
rect 52730 10004 52736 10016
rect 52788 10004 52794 10056
rect 57790 10004 57796 10056
rect 57848 10044 57854 10056
rect 57977 10047 58035 10053
rect 57977 10044 57989 10047
rect 57848 10016 57989 10044
rect 57848 10004 57854 10016
rect 57977 10013 57989 10016
rect 58023 10013 58035 10047
rect 57977 10007 58035 10013
rect 58158 10004 58164 10056
rect 58216 10044 58222 10056
rect 71498 10044 71504 10056
rect 58216 10016 71504 10044
rect 58216 10004 58222 10016
rect 71498 10004 71504 10016
rect 71556 10004 71562 10056
rect 71792 10044 71820 10084
rect 75086 10072 75092 10124
rect 75144 10112 75150 10124
rect 81161 10115 81219 10121
rect 81161 10112 81173 10115
rect 75144 10084 81173 10112
rect 75144 10072 75150 10084
rect 81161 10081 81173 10084
rect 81207 10081 81219 10115
rect 81710 10112 81716 10124
rect 81671 10084 81716 10112
rect 81161 10075 81219 10081
rect 81710 10072 81716 10084
rect 81768 10072 81774 10124
rect 95881 10047 95939 10053
rect 95881 10044 95893 10047
rect 71792 10016 80054 10044
rect 43990 9976 43996 9988
rect 37608 9948 38148 9976
rect 39040 9948 43996 9976
rect 37608 9936 37614 9948
rect 39040 9908 39068 9948
rect 43990 9936 43996 9948
rect 44048 9936 44054 9988
rect 44082 9936 44088 9988
rect 44140 9976 44146 9988
rect 53558 9976 53564 9988
rect 44140 9948 53564 9976
rect 44140 9936 44146 9948
rect 53558 9936 53564 9948
rect 53616 9936 53622 9988
rect 57425 9979 57483 9985
rect 57425 9945 57437 9979
rect 57471 9976 57483 9979
rect 66530 9976 66536 9988
rect 57471 9948 66536 9976
rect 57471 9945 57483 9948
rect 57425 9939 57483 9945
rect 66530 9936 66536 9948
rect 66588 9976 66594 9988
rect 75270 9976 75276 9988
rect 66588 9948 75276 9976
rect 66588 9936 66594 9948
rect 75270 9936 75276 9948
rect 75328 9936 75334 9988
rect 80026 9976 80054 10016
rect 89686 10016 95893 10044
rect 89686 9976 89714 10016
rect 95881 10013 95893 10016
rect 95927 10013 95939 10047
rect 95881 10007 95939 10013
rect 96890 9976 96896 9988
rect 80026 9948 89714 9976
rect 93826 9948 96896 9976
rect 39666 9908 39672 9920
rect 36556 9880 39068 9908
rect 39627 9880 39672 9908
rect 39666 9868 39672 9880
rect 39724 9868 39730 9920
rect 39850 9868 39856 9920
rect 39908 9908 39914 9920
rect 42794 9908 42800 9920
rect 39908 9880 42800 9908
rect 39908 9868 39914 9880
rect 42794 9868 42800 9880
rect 42852 9868 42858 9920
rect 42886 9868 42892 9920
rect 42944 9908 42950 9920
rect 50982 9908 50988 9920
rect 42944 9880 50988 9908
rect 42944 9868 42950 9880
rect 50982 9868 50988 9880
rect 51040 9868 51046 9920
rect 52457 9911 52515 9917
rect 52457 9877 52469 9911
rect 52503 9908 52515 9911
rect 55122 9908 55128 9920
rect 52503 9880 55128 9908
rect 52503 9877 52515 9880
rect 52457 9871 52515 9877
rect 55122 9868 55128 9880
rect 55180 9868 55186 9920
rect 59541 9911 59599 9917
rect 59541 9877 59553 9911
rect 59587 9908 59599 9911
rect 93826 9908 93854 9948
rect 96890 9936 96896 9948
rect 96948 9936 96954 9988
rect 59587 9880 93854 9908
rect 59587 9877 59599 9880
rect 59541 9871 59599 9877
rect 1104 9818 98808 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 65686 9818
rect 65738 9766 65750 9818
rect 65802 9766 65814 9818
rect 65866 9766 65878 9818
rect 65930 9766 96406 9818
rect 96458 9766 96470 9818
rect 96522 9766 96534 9818
rect 96586 9766 96598 9818
rect 96650 9766 98808 9818
rect 1104 9744 98808 9766
rect 12360 9676 13124 9704
rect 12360 9568 12388 9676
rect 12618 9596 12624 9648
rect 12676 9636 12682 9648
rect 12989 9639 13047 9645
rect 12989 9636 13001 9639
rect 12676 9608 13001 9636
rect 12676 9596 12682 9608
rect 12989 9605 13001 9608
rect 13035 9605 13047 9639
rect 13096 9636 13124 9676
rect 20180 9676 20484 9704
rect 14734 9636 14740 9648
rect 13096 9608 14740 9636
rect 12989 9599 13047 9605
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 18506 9596 18512 9648
rect 18564 9636 18570 9648
rect 20180 9636 20208 9676
rect 20346 9636 20352 9648
rect 18564 9608 20208 9636
rect 20307 9608 20352 9636
rect 18564 9596 18570 9608
rect 20346 9596 20352 9608
rect 20404 9596 20410 9648
rect 20456 9636 20484 9676
rect 20622 9664 20628 9716
rect 20680 9704 20686 9716
rect 62666 9704 62672 9716
rect 20680 9676 62672 9704
rect 20680 9664 20686 9676
rect 62666 9664 62672 9676
rect 62724 9664 62730 9716
rect 63402 9664 63408 9716
rect 63460 9704 63466 9716
rect 68278 9704 68284 9716
rect 63460 9676 68284 9704
rect 63460 9664 63466 9676
rect 68278 9664 68284 9676
rect 68336 9664 68342 9716
rect 68370 9664 68376 9716
rect 68428 9704 68434 9716
rect 73062 9704 73068 9716
rect 68428 9676 73068 9704
rect 68428 9664 68434 9676
rect 73062 9664 73068 9676
rect 73120 9664 73126 9716
rect 20456 9608 36860 9636
rect 13630 9568 13636 9580
rect 12360 9540 12480 9568
rect 3234 9500 3240 9512
rect 3195 9472 3240 9500
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 3418 9500 3424 9512
rect 3379 9472 3424 9500
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 3602 9500 3608 9512
rect 3563 9472 3608 9500
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 12452 9509 12480 9540
rect 12544 9540 13636 9568
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 3694 9432 3700 9444
rect 3655 9404 3700 9432
rect 3694 9392 3700 9404
rect 3752 9392 3758 9444
rect 5258 9392 5264 9444
rect 5316 9432 5322 9444
rect 12544 9432 12572 9540
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9568 18935 9571
rect 19242 9568 19248 9580
rect 18923 9540 19248 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 19242 9528 19248 9540
rect 19300 9568 19306 9580
rect 19337 9571 19395 9577
rect 19337 9568 19349 9571
rect 19300 9540 19349 9568
rect 19300 9528 19306 9540
rect 19337 9537 19349 9540
rect 19383 9537 19395 9571
rect 19337 9531 19395 9537
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9568 19487 9571
rect 31570 9568 31576 9580
rect 19475 9540 31576 9568
rect 19475 9537 19487 9540
rect 19429 9531 19487 9537
rect 31570 9528 31576 9540
rect 31628 9528 31634 9580
rect 35529 9571 35587 9577
rect 35529 9537 35541 9571
rect 35575 9568 35587 9571
rect 35802 9568 35808 9580
rect 35575 9540 35808 9568
rect 35575 9537 35587 9540
rect 35529 9531 35587 9537
rect 35802 9528 35808 9540
rect 35860 9528 35866 9580
rect 12710 9500 12716 9512
rect 12671 9472 12716 9500
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9500 12863 9503
rect 15102 9500 15108 9512
rect 12851 9472 15108 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 18782 9460 18788 9512
rect 18840 9500 18846 9512
rect 19153 9503 19211 9509
rect 19153 9500 19165 9503
rect 18840 9472 19165 9500
rect 18840 9460 18846 9472
rect 19153 9469 19165 9472
rect 19199 9469 19211 9503
rect 19518 9500 19524 9512
rect 19479 9472 19524 9500
rect 19153 9463 19211 9469
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 26878 9500 26884 9512
rect 19751 9472 26884 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 26878 9460 26884 9472
rect 26936 9460 26942 9512
rect 35986 9500 35992 9512
rect 35947 9472 35992 9500
rect 35986 9460 35992 9472
rect 36044 9460 36050 9512
rect 36262 9500 36268 9512
rect 36223 9472 36268 9500
rect 36262 9460 36268 9472
rect 36320 9460 36326 9512
rect 36357 9503 36415 9509
rect 36357 9469 36369 9503
rect 36403 9500 36415 9503
rect 36538 9500 36544 9512
rect 36403 9472 36544 9500
rect 36403 9469 36415 9472
rect 36357 9463 36415 9469
rect 36538 9460 36544 9472
rect 36596 9460 36602 9512
rect 36832 9509 36860 9608
rect 36906 9596 36912 9648
rect 36964 9636 36970 9648
rect 89714 9636 89720 9648
rect 36964 9608 89720 9636
rect 36964 9596 36970 9608
rect 89714 9596 89720 9608
rect 89772 9596 89778 9648
rect 37366 9528 37372 9580
rect 37424 9568 37430 9580
rect 50893 9571 50951 9577
rect 50893 9568 50905 9571
rect 37424 9540 50905 9568
rect 37424 9528 37430 9540
rect 50893 9537 50905 9540
rect 50939 9537 50951 9571
rect 54294 9568 54300 9580
rect 54255 9540 54300 9568
rect 50893 9531 50951 9537
rect 54294 9528 54300 9540
rect 54352 9528 54358 9580
rect 54754 9528 54760 9580
rect 54812 9568 54818 9580
rect 72970 9568 72976 9580
rect 54812 9540 72976 9568
rect 54812 9528 54818 9540
rect 72970 9528 72976 9540
rect 73028 9528 73034 9580
rect 78674 9528 78680 9580
rect 78732 9568 78738 9580
rect 82354 9568 82360 9580
rect 78732 9540 82360 9568
rect 78732 9528 78738 9540
rect 82354 9528 82360 9540
rect 82412 9568 82418 9580
rect 95510 9568 95516 9580
rect 82412 9540 95516 9568
rect 82412 9528 82418 9540
rect 95510 9528 95516 9540
rect 95568 9528 95574 9580
rect 36633 9503 36691 9509
rect 36633 9469 36645 9503
rect 36679 9469 36691 9503
rect 36633 9463 36691 9469
rect 36817 9503 36875 9509
rect 36817 9469 36829 9503
rect 36863 9469 36875 9503
rect 36817 9463 36875 9469
rect 12621 9435 12679 9441
rect 12621 9432 12633 9435
rect 5316 9404 6914 9432
rect 12544 9404 12633 9432
rect 5316 9392 5322 9404
rect 6886 9364 6914 9404
rect 12621 9401 12633 9404
rect 12667 9401 12679 9435
rect 36648 9432 36676 9463
rect 37274 9460 37280 9512
rect 37332 9500 37338 9512
rect 37332 9472 39344 9500
rect 37332 9460 37338 9472
rect 37826 9432 37832 9444
rect 12621 9395 12679 9401
rect 12912 9404 35848 9432
rect 36648 9404 37832 9432
rect 12912 9364 12940 9404
rect 6886 9336 12940 9364
rect 18969 9367 19027 9373
rect 18969 9333 18981 9367
rect 19015 9364 19027 9367
rect 23382 9364 23388 9376
rect 19015 9336 23388 9364
rect 19015 9333 19027 9336
rect 18969 9327 19027 9333
rect 23382 9324 23388 9336
rect 23440 9324 23446 9376
rect 25866 9324 25872 9376
rect 25924 9364 25930 9376
rect 26234 9364 26240 9376
rect 25924 9336 26240 9364
rect 25924 9324 25930 9336
rect 26234 9324 26240 9336
rect 26292 9324 26298 9376
rect 35820 9364 35848 9404
rect 37826 9392 37832 9404
rect 37884 9392 37890 9444
rect 39316 9432 39344 9472
rect 44910 9460 44916 9512
rect 44968 9500 44974 9512
rect 50617 9503 50675 9509
rect 50617 9500 50629 9503
rect 44968 9472 50629 9500
rect 44968 9460 44974 9472
rect 50617 9469 50629 9472
rect 50663 9469 50675 9503
rect 51074 9500 51080 9512
rect 51035 9472 51080 9500
rect 50617 9463 50675 9469
rect 51074 9460 51080 9472
rect 51132 9460 51138 9512
rect 51353 9503 51411 9509
rect 51353 9469 51365 9503
rect 51399 9500 51411 9503
rect 51534 9500 51540 9512
rect 51399 9472 51540 9500
rect 51399 9469 51411 9472
rect 51353 9463 51411 9469
rect 51534 9460 51540 9472
rect 51592 9460 51598 9512
rect 52273 9503 52331 9509
rect 52273 9469 52285 9503
rect 52319 9500 52331 9503
rect 53926 9500 53932 9512
rect 52319 9472 53932 9500
rect 52319 9469 52331 9472
rect 52273 9463 52331 9469
rect 53926 9460 53932 9472
rect 53984 9460 53990 9512
rect 54021 9503 54079 9509
rect 54021 9469 54033 9503
rect 54067 9500 54079 9503
rect 57330 9500 57336 9512
rect 54067 9472 57336 9500
rect 54067 9469 54079 9472
rect 54021 9463 54079 9469
rect 57330 9460 57336 9472
rect 57388 9460 57394 9512
rect 62390 9500 62396 9512
rect 60706 9472 62396 9500
rect 40494 9432 40500 9444
rect 39316 9404 40500 9432
rect 40494 9392 40500 9404
rect 40552 9392 40558 9444
rect 60706 9432 60734 9472
rect 62390 9460 62396 9472
rect 62448 9460 62454 9512
rect 62482 9460 62488 9512
rect 62540 9500 62546 9512
rect 63218 9500 63224 9512
rect 62540 9472 63224 9500
rect 62540 9460 62546 9472
rect 63218 9460 63224 9472
rect 63276 9460 63282 9512
rect 63310 9460 63316 9512
rect 63368 9500 63374 9512
rect 67174 9500 67180 9512
rect 63368 9472 67180 9500
rect 63368 9460 63374 9472
rect 67174 9460 67180 9472
rect 67232 9460 67238 9512
rect 67361 9503 67419 9509
rect 67361 9469 67373 9503
rect 67407 9500 67419 9503
rect 86954 9500 86960 9512
rect 67407 9472 86960 9500
rect 67407 9469 67419 9472
rect 67361 9463 67419 9469
rect 86954 9460 86960 9472
rect 87012 9460 87018 9512
rect 90726 9500 90732 9512
rect 90687 9472 90732 9500
rect 90726 9460 90732 9472
rect 90784 9460 90790 9512
rect 90818 9460 90824 9512
rect 90876 9500 90882 9512
rect 91005 9503 91063 9509
rect 90876 9472 90921 9500
rect 90876 9460 90882 9472
rect 91005 9469 91017 9503
rect 91051 9469 91063 9503
rect 91005 9463 91063 9469
rect 41432 9404 60734 9432
rect 41432 9364 41460 9404
rect 62850 9392 62856 9444
rect 62908 9432 62914 9444
rect 65334 9432 65340 9444
rect 62908 9404 65340 9432
rect 62908 9392 62914 9404
rect 65334 9392 65340 9404
rect 65392 9392 65398 9444
rect 65518 9392 65524 9444
rect 65576 9432 65582 9444
rect 68278 9432 68284 9444
rect 65576 9404 68284 9432
rect 65576 9392 65582 9404
rect 68278 9392 68284 9404
rect 68336 9432 68342 9444
rect 68738 9432 68744 9444
rect 68336 9404 68744 9432
rect 68336 9392 68342 9404
rect 68738 9392 68744 9404
rect 68796 9392 68802 9444
rect 73890 9392 73896 9444
rect 73948 9432 73954 9444
rect 91020 9432 91048 9463
rect 73948 9404 91048 9432
rect 73948 9392 73954 9404
rect 35820 9336 41460 9364
rect 41506 9324 41512 9376
rect 41564 9364 41570 9376
rect 49326 9364 49332 9376
rect 41564 9336 49332 9364
rect 41564 9324 41570 9336
rect 49326 9324 49332 9336
rect 49384 9324 49390 9376
rect 50617 9367 50675 9373
rect 50617 9333 50629 9367
rect 50663 9364 50675 9367
rect 50801 9367 50859 9373
rect 50801 9364 50813 9367
rect 50663 9336 50813 9364
rect 50663 9333 50675 9336
rect 50617 9327 50675 9333
rect 50801 9333 50813 9336
rect 50847 9364 50859 9367
rect 51261 9367 51319 9373
rect 51261 9364 51273 9367
rect 50847 9336 51273 9364
rect 50847 9333 50859 9336
rect 50801 9327 50859 9333
rect 51261 9333 51273 9336
rect 51307 9364 51319 9367
rect 71866 9364 71872 9376
rect 51307 9336 71872 9364
rect 51307 9333 51319 9336
rect 51261 9327 51319 9333
rect 71866 9324 71872 9336
rect 71924 9324 71930 9376
rect 85942 9324 85948 9376
rect 86000 9364 86006 9376
rect 91189 9367 91247 9373
rect 91189 9364 91201 9367
rect 86000 9336 91201 9364
rect 86000 9324 86006 9336
rect 91189 9333 91201 9336
rect 91235 9333 91247 9367
rect 91189 9327 91247 9333
rect 1104 9274 98808 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 50326 9274
rect 50378 9222 50390 9274
rect 50442 9222 50454 9274
rect 50506 9222 50518 9274
rect 50570 9222 81046 9274
rect 81098 9222 81110 9274
rect 81162 9222 81174 9274
rect 81226 9222 81238 9274
rect 81290 9222 98808 9274
rect 1104 9200 98808 9222
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 11425 9163 11483 9169
rect 11425 9160 11437 9163
rect 11020 9132 11437 9160
rect 11020 9120 11026 9132
rect 11425 9129 11437 9132
rect 11471 9160 11483 9163
rect 12250 9160 12256 9172
rect 11471 9132 12020 9160
rect 12211 9132 12256 9160
rect 11471 9129 11483 9132
rect 11425 9123 11483 9129
rect 5350 9052 5356 9104
rect 5408 9052 5414 9104
rect 5997 9095 6055 9101
rect 5997 9061 6009 9095
rect 6043 9092 6055 9095
rect 9030 9092 9036 9104
rect 6043 9064 9036 9092
rect 6043 9061 6055 9064
rect 5997 9055 6055 9061
rect 9030 9052 9036 9064
rect 9088 9052 9094 9104
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 9024 4767 9027
rect 4798 9024 4804 9036
rect 4755 8996 4804 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 5074 9024 5080 9036
rect 5035 8996 5080 9024
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5368 9024 5396 9052
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 5368 8996 5457 9024
rect 5445 8993 5457 8996
rect 5491 8993 5503 9027
rect 5445 8987 5503 8993
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 7466 9024 7472 9036
rect 5675 8996 7472 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 11606 9024 11612 9036
rect 11567 8996 11612 9024
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 11790 9024 11796 9036
rect 11751 8996 11796 9024
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 11992 9033 12020 9132
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 16666 9160 16672 9172
rect 16627 9132 16672 9160
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 19392 9132 22094 9160
rect 19392 9120 19398 9132
rect 22066 9092 22094 9132
rect 30374 9120 30380 9172
rect 30432 9160 30438 9172
rect 36906 9160 36912 9172
rect 30432 9132 36912 9160
rect 30432 9120 30438 9132
rect 36906 9120 36912 9132
rect 36964 9120 36970 9172
rect 49878 9120 49884 9172
rect 49936 9160 49942 9172
rect 50798 9160 50804 9172
rect 49936 9132 50804 9160
rect 49936 9120 49942 9132
rect 50798 9120 50804 9132
rect 50856 9160 50862 9172
rect 51074 9160 51080 9172
rect 50856 9132 51080 9160
rect 50856 9120 50862 9132
rect 51074 9120 51080 9132
rect 51132 9120 51138 9172
rect 54478 9120 54484 9172
rect 54536 9160 54542 9172
rect 54536 9132 70394 9160
rect 54536 9120 54542 9132
rect 36998 9092 37004 9104
rect 22066 9064 37004 9092
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 8993 12035 9027
rect 12158 9024 12164 9036
rect 12119 8996 12164 9024
rect 11977 8987 12035 8993
rect 12158 8984 12164 8996
rect 12216 9024 12222 9036
rect 12437 9027 12495 9033
rect 12437 9024 12449 9027
rect 12216 8996 12449 9024
rect 12216 8984 12222 8996
rect 12437 8993 12449 8996
rect 12483 8993 12495 9027
rect 12437 8987 12495 8993
rect 16390 8984 16396 9036
rect 16448 9024 16454 9036
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 16448 8996 16497 9024
rect 16448 8984 16454 8996
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 16761 9027 16819 9033
rect 16761 8993 16773 9027
rect 16807 9024 16819 9027
rect 35710 9024 35716 9036
rect 16807 8996 35716 9024
rect 16807 8993 16819 8996
rect 16761 8987 16819 8993
rect 35710 8984 35716 8996
rect 35768 8984 35774 9036
rect 36924 9033 36952 9064
rect 36998 9052 37004 9064
rect 37056 9052 37062 9104
rect 37274 9052 37280 9104
rect 37332 9092 37338 9104
rect 37642 9092 37648 9104
rect 37332 9064 37504 9092
rect 37332 9052 37338 9064
rect 36909 9027 36967 9033
rect 36909 8993 36921 9027
rect 36955 8993 36967 9027
rect 36909 8987 36967 8993
rect 37092 9027 37150 9033
rect 37092 8993 37104 9027
rect 37138 9024 37150 9027
rect 37366 9024 37372 9036
rect 37138 8996 37372 9024
rect 37138 8993 37150 8996
rect 37092 8987 37150 8993
rect 37366 8984 37372 8996
rect 37424 8984 37430 9036
rect 37476 9033 37504 9064
rect 37568 9064 37648 9092
rect 37461 9027 37519 9033
rect 37461 8993 37473 9027
rect 37507 8993 37519 9027
rect 37461 8987 37519 8993
rect 5166 8956 5172 8968
rect 5127 8928 5172 8956
rect 5166 8916 5172 8928
rect 5224 8956 5230 8968
rect 11885 8959 11943 8965
rect 5224 8928 6914 8956
rect 5224 8916 5230 8928
rect 6886 8820 6914 8928
rect 11885 8925 11897 8959
rect 11931 8925 11943 8959
rect 11885 8919 11943 8925
rect 11514 8848 11520 8900
rect 11572 8888 11578 8900
rect 11900 8888 11928 8919
rect 15010 8916 15016 8968
rect 15068 8956 15074 8968
rect 20809 8959 20867 8965
rect 20809 8956 20821 8959
rect 15068 8928 20821 8956
rect 15068 8916 15074 8928
rect 20809 8925 20821 8928
rect 20855 8925 20867 8959
rect 20809 8919 20867 8925
rect 21085 8959 21143 8965
rect 21085 8925 21097 8959
rect 21131 8956 21143 8959
rect 21266 8956 21272 8968
rect 21131 8928 21272 8956
rect 21131 8925 21143 8928
rect 21085 8919 21143 8925
rect 17678 8888 17684 8900
rect 11572 8860 11928 8888
rect 12406 8860 17684 8888
rect 11572 8848 11578 8860
rect 12406 8820 12434 8860
rect 17678 8848 17684 8860
rect 17736 8848 17742 8900
rect 6886 8792 12434 8820
rect 15654 8780 15660 8832
rect 15712 8820 15718 8832
rect 16301 8823 16359 8829
rect 16301 8820 16313 8823
rect 15712 8792 16313 8820
rect 15712 8780 15718 8792
rect 16301 8789 16313 8792
rect 16347 8789 16359 8823
rect 20824 8820 20852 8919
rect 21266 8916 21272 8928
rect 21324 8916 21330 8968
rect 35894 8916 35900 8968
rect 35952 8956 35958 8968
rect 37185 8959 37243 8965
rect 37185 8956 37197 8959
rect 35952 8928 37197 8956
rect 35952 8916 35958 8928
rect 37185 8925 37197 8928
rect 37231 8925 37243 8959
rect 37185 8919 37243 8925
rect 37277 8959 37335 8965
rect 37277 8925 37289 8959
rect 37323 8956 37335 8959
rect 37568 8956 37596 9064
rect 37642 9052 37648 9064
rect 37700 9052 37706 9104
rect 39758 9092 39764 9104
rect 39719 9064 39764 9092
rect 39758 9052 39764 9064
rect 39816 9052 39822 9104
rect 42610 9052 42616 9104
rect 42668 9092 42674 9104
rect 42668 9064 47808 9092
rect 42668 9052 42674 9064
rect 37734 8984 37740 9036
rect 37792 9024 37798 9036
rect 38381 9027 38439 9033
rect 38381 9024 38393 9027
rect 37792 8996 38393 9024
rect 37792 8984 37798 8996
rect 38381 8993 38393 8996
rect 38427 8993 38439 9027
rect 38381 8987 38439 8993
rect 40310 8984 40316 9036
rect 40368 9024 40374 9036
rect 44726 9024 44732 9036
rect 40368 8996 44732 9024
rect 40368 8984 40374 8996
rect 44726 8984 44732 8996
rect 44784 8984 44790 9036
rect 37323 8928 37596 8956
rect 37323 8925 37335 8928
rect 37277 8919 37335 8925
rect 37642 8916 37648 8968
rect 37700 8956 37706 8968
rect 38105 8959 38163 8965
rect 38105 8956 38117 8959
rect 37700 8928 38117 8956
rect 37700 8916 37706 8928
rect 38105 8925 38117 8928
rect 38151 8925 38163 8959
rect 38105 8919 38163 8925
rect 43070 8916 43076 8968
rect 43128 8956 43134 8968
rect 47780 8956 47808 9064
rect 56778 9052 56784 9104
rect 56836 9092 56842 9104
rect 59262 9092 59268 9104
rect 56836 9064 59268 9092
rect 56836 9052 56842 9064
rect 59262 9052 59268 9064
rect 59320 9052 59326 9104
rect 59446 9052 59452 9104
rect 59504 9092 59510 9104
rect 62850 9092 62856 9104
rect 59504 9064 62856 9092
rect 59504 9052 59510 9064
rect 62850 9052 62856 9064
rect 62908 9052 62914 9104
rect 63862 9052 63868 9104
rect 63920 9092 63926 9104
rect 67358 9092 67364 9104
rect 63920 9064 67364 9092
rect 63920 9052 63926 9064
rect 67358 9052 67364 9064
rect 67416 9052 67422 9104
rect 70366 9092 70394 9132
rect 74258 9120 74264 9172
rect 74316 9160 74322 9172
rect 74445 9163 74503 9169
rect 74445 9160 74457 9163
rect 74316 9132 74457 9160
rect 74316 9120 74322 9132
rect 74445 9129 74457 9132
rect 74491 9129 74503 9163
rect 74445 9123 74503 9129
rect 87046 9092 87052 9104
rect 70366 9064 87052 9092
rect 87046 9052 87052 9064
rect 87104 9052 87110 9104
rect 88518 9052 88524 9104
rect 88576 9092 88582 9104
rect 94130 9092 94136 9104
rect 88576 9064 89484 9092
rect 88576 9052 88582 9064
rect 48406 8984 48412 9036
rect 48464 9024 48470 9036
rect 63034 9024 63040 9036
rect 48464 8996 62896 9024
rect 62995 8996 63040 9024
rect 48464 8984 48470 8996
rect 62022 8956 62028 8968
rect 43128 8928 47716 8956
rect 47780 8928 62028 8956
rect 43128 8916 43134 8928
rect 26878 8848 26884 8900
rect 26936 8888 26942 8900
rect 47578 8888 47584 8900
rect 26936 8860 37688 8888
rect 26936 8848 26942 8860
rect 21726 8820 21732 8832
rect 20824 8792 21732 8820
rect 16301 8783 16359 8789
rect 21726 8780 21732 8792
rect 21784 8780 21790 8832
rect 22094 8780 22100 8832
rect 22152 8820 22158 8832
rect 22189 8823 22247 8829
rect 22189 8820 22201 8823
rect 22152 8792 22201 8820
rect 22152 8780 22158 8792
rect 22189 8789 22201 8792
rect 22235 8789 22247 8823
rect 22189 8783 22247 8789
rect 33686 8780 33692 8832
rect 33744 8820 33750 8832
rect 33962 8820 33968 8832
rect 33744 8792 33968 8820
rect 33744 8780 33750 8792
rect 33962 8780 33968 8792
rect 34020 8780 34026 8832
rect 37550 8820 37556 8832
rect 37511 8792 37556 8820
rect 37550 8780 37556 8792
rect 37608 8780 37614 8832
rect 37660 8820 37688 8860
rect 39040 8860 47584 8888
rect 39040 8820 39068 8860
rect 47578 8848 47584 8860
rect 47636 8848 47642 8900
rect 47688 8888 47716 8928
rect 62022 8916 62028 8928
rect 62080 8916 62086 8968
rect 62761 8959 62819 8965
rect 62761 8925 62773 8959
rect 62807 8925 62819 8959
rect 62868 8956 62896 8996
rect 63034 8984 63040 8996
rect 63092 8984 63098 9036
rect 73801 9027 73859 9033
rect 73801 9024 73813 9027
rect 63144 8996 73813 9024
rect 63144 8956 63172 8996
rect 73801 8993 73813 8996
rect 73847 8993 73859 9027
rect 87064 9024 87092 9052
rect 88797 9027 88855 9033
rect 88797 9024 88809 9027
rect 87064 8996 88809 9024
rect 73801 8987 73859 8993
rect 88797 8993 88809 8996
rect 88843 8993 88855 9027
rect 88978 9024 88984 9036
rect 88939 8996 88984 9024
rect 88797 8987 88855 8993
rect 88978 8984 88984 8996
rect 89036 8984 89042 9036
rect 89346 9024 89352 9036
rect 89307 8996 89352 9024
rect 89346 8984 89352 8996
rect 89404 8984 89410 9036
rect 89456 9033 89484 9064
rect 89686 9064 94136 9092
rect 89441 9027 89499 9033
rect 89441 8993 89453 9027
rect 89487 8993 89499 9027
rect 89441 8987 89499 8993
rect 62868 8928 63172 8956
rect 62761 8919 62819 8925
rect 55306 8888 55312 8900
rect 47688 8860 55312 8888
rect 55306 8848 55312 8860
rect 55364 8848 55370 8900
rect 55582 8848 55588 8900
rect 55640 8888 55646 8900
rect 56778 8888 56784 8900
rect 55640 8860 56784 8888
rect 55640 8848 55646 8860
rect 56778 8848 56784 8860
rect 56836 8848 56842 8900
rect 58066 8848 58072 8900
rect 58124 8888 58130 8900
rect 61654 8888 61660 8900
rect 58124 8860 61660 8888
rect 58124 8848 58130 8860
rect 61654 8848 61660 8860
rect 61712 8848 61718 8900
rect 61746 8848 61752 8900
rect 61804 8888 61810 8900
rect 62776 8888 62804 8919
rect 63218 8916 63224 8968
rect 63276 8956 63282 8968
rect 64141 8959 64199 8965
rect 64141 8956 64153 8959
rect 63276 8928 64153 8956
rect 63276 8916 63282 8928
rect 64141 8925 64153 8928
rect 64187 8925 64199 8959
rect 64141 8919 64199 8925
rect 65518 8916 65524 8968
rect 65576 8956 65582 8968
rect 73948 8959 74006 8965
rect 73948 8956 73960 8959
rect 65576 8928 73960 8956
rect 65576 8916 65582 8928
rect 73948 8925 73960 8928
rect 73994 8925 74006 8959
rect 74166 8956 74172 8968
rect 74127 8928 74172 8956
rect 73948 8919 74006 8925
rect 74166 8916 74172 8928
rect 74224 8916 74230 8968
rect 88426 8956 88432 8968
rect 88387 8928 88432 8956
rect 88426 8916 88432 8928
rect 88484 8916 88490 8968
rect 74077 8891 74135 8897
rect 74077 8888 74089 8891
rect 61804 8860 62804 8888
rect 64064 8860 74089 8888
rect 61804 8848 61810 8860
rect 37660 8792 39068 8820
rect 45002 8780 45008 8832
rect 45060 8820 45066 8832
rect 51810 8820 51816 8832
rect 45060 8792 51816 8820
rect 45060 8780 45066 8792
rect 51810 8780 51816 8792
rect 51868 8780 51874 8832
rect 52362 8780 52368 8832
rect 52420 8820 52426 8832
rect 64064 8820 64092 8860
rect 74077 8857 74089 8860
rect 74123 8857 74135 8891
rect 89686 8888 89714 9064
rect 94130 9052 94136 9064
rect 94188 9052 94194 9104
rect 95510 9092 95516 9104
rect 95471 9064 95516 9092
rect 95510 9052 95516 9064
rect 95568 9052 95574 9104
rect 95142 9024 95148 9036
rect 95103 8996 95148 9024
rect 95142 8984 95148 8996
rect 95200 8984 95206 9036
rect 74077 8851 74135 8857
rect 80026 8860 89714 8888
rect 52420 8792 64092 8820
rect 52420 8780 52426 8792
rect 64506 8780 64512 8832
rect 64564 8820 64570 8832
rect 80026 8820 80054 8860
rect 64564 8792 80054 8820
rect 64564 8780 64570 8792
rect 89714 8780 89720 8832
rect 89772 8820 89778 8832
rect 94866 8820 94872 8832
rect 89772 8792 94872 8820
rect 89772 8780 89778 8792
rect 94866 8780 94872 8792
rect 94924 8780 94930 8832
rect 1104 8730 98808 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 65686 8730
rect 65738 8678 65750 8730
rect 65802 8678 65814 8730
rect 65866 8678 65878 8730
rect 65930 8678 96406 8730
rect 96458 8678 96470 8730
rect 96522 8678 96534 8730
rect 96586 8678 96598 8730
rect 96650 8678 98808 8730
rect 1104 8656 98808 8678
rect 20438 8616 20444 8628
rect 20399 8588 20444 8616
rect 20438 8576 20444 8588
rect 20496 8576 20502 8628
rect 23658 8616 23664 8628
rect 23619 8588 23664 8616
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 33410 8576 33416 8628
rect 33468 8616 33474 8628
rect 39390 8616 39396 8628
rect 33468 8588 39396 8616
rect 33468 8576 33474 8588
rect 39390 8576 39396 8588
rect 39448 8576 39454 8628
rect 39485 8619 39543 8625
rect 39485 8585 39497 8619
rect 39531 8616 39543 8619
rect 39942 8616 39948 8628
rect 39531 8588 39948 8616
rect 39531 8585 39543 8588
rect 39485 8579 39543 8585
rect 39942 8576 39948 8588
rect 40000 8576 40006 8628
rect 41322 8576 41328 8628
rect 41380 8616 41386 8628
rect 46474 8616 46480 8628
rect 41380 8588 46480 8616
rect 41380 8576 41386 8588
rect 46474 8576 46480 8588
rect 46532 8576 46538 8628
rect 47670 8576 47676 8628
rect 47728 8616 47734 8628
rect 47728 8588 50936 8616
rect 47728 8576 47734 8588
rect 23124 8520 33548 8548
rect 19886 8440 19892 8492
rect 19944 8480 19950 8492
rect 20073 8483 20131 8489
rect 20073 8480 20085 8483
rect 19944 8452 20085 8480
rect 19944 8440 19950 8452
rect 20073 8449 20085 8452
rect 20119 8449 20131 8483
rect 20073 8443 20131 8449
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8480 20223 8483
rect 20254 8480 20260 8492
rect 20211 8452 20260 8480
rect 20211 8449 20223 8452
rect 20165 8443 20223 8449
rect 20254 8440 20260 8452
rect 20312 8440 20318 8492
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 19797 8415 19855 8421
rect 19797 8412 19809 8415
rect 19392 8384 19809 8412
rect 19392 8372 19398 8384
rect 19797 8381 19809 8384
rect 19843 8381 19855 8415
rect 19978 8412 19984 8424
rect 19939 8384 19984 8412
rect 19797 8375 19855 8381
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 20349 8415 20407 8421
rect 20349 8412 20361 8415
rect 20088 8384 20361 8412
rect 6638 8304 6644 8356
rect 6696 8344 6702 8356
rect 9214 8344 9220 8356
rect 6696 8316 9220 8344
rect 6696 8304 6702 8316
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 16206 8304 16212 8356
rect 16264 8344 16270 8356
rect 16482 8344 16488 8356
rect 16264 8316 16488 8344
rect 16264 8304 16270 8316
rect 16482 8304 16488 8316
rect 16540 8344 16546 8356
rect 20088 8344 20116 8384
rect 20349 8381 20361 8384
rect 20395 8381 20407 8415
rect 23014 8412 23020 8424
rect 22975 8384 23020 8412
rect 20349 8375 20407 8381
rect 23014 8372 23020 8384
rect 23072 8372 23078 8424
rect 23124 8421 23152 8520
rect 31846 8480 31852 8492
rect 23308 8452 31852 8480
rect 23308 8421 23336 8452
rect 31846 8440 31852 8452
rect 31904 8440 31910 8492
rect 33520 8480 33548 8520
rect 33704 8520 38654 8548
rect 33704 8480 33732 8520
rect 34330 8480 34336 8492
rect 33520 8452 33732 8480
rect 34291 8452 34336 8480
rect 34330 8440 34336 8452
rect 34388 8440 34394 8492
rect 34606 8440 34612 8492
rect 34664 8480 34670 8492
rect 38626 8480 38654 8520
rect 40402 8508 40408 8560
rect 40460 8548 40466 8560
rect 50798 8548 50804 8560
rect 40460 8520 50804 8548
rect 40460 8508 40466 8520
rect 50798 8508 50804 8520
rect 50856 8508 50862 8560
rect 50908 8548 50936 8588
rect 56594 8576 56600 8628
rect 56652 8616 56658 8628
rect 60734 8616 60740 8628
rect 56652 8588 60740 8616
rect 56652 8576 56658 8588
rect 60734 8576 60740 8588
rect 60792 8576 60798 8628
rect 60826 8576 60832 8628
rect 60884 8616 60890 8628
rect 67269 8619 67327 8625
rect 67269 8616 67281 8619
rect 60884 8588 67281 8616
rect 60884 8576 60890 8588
rect 67269 8585 67281 8588
rect 67315 8585 67327 8619
rect 67269 8579 67327 8585
rect 67358 8576 67364 8628
rect 67416 8616 67422 8628
rect 78950 8616 78956 8628
rect 67416 8588 78956 8616
rect 67416 8576 67422 8588
rect 78950 8576 78956 8588
rect 79008 8576 79014 8628
rect 94130 8616 94136 8628
rect 94091 8588 94136 8616
rect 94130 8576 94136 8588
rect 94188 8576 94194 8628
rect 94593 8619 94651 8625
rect 94593 8585 94605 8619
rect 94639 8616 94651 8619
rect 95145 8619 95203 8625
rect 95145 8616 95157 8619
rect 94639 8588 95157 8616
rect 94639 8585 94651 8588
rect 94593 8579 94651 8585
rect 95145 8585 95157 8588
rect 95191 8585 95203 8619
rect 95145 8579 95203 8585
rect 50908 8520 51212 8548
rect 47486 8480 47492 8492
rect 34664 8452 35572 8480
rect 38626 8452 47492 8480
rect 34664 8440 34670 8452
rect 23110 8415 23168 8421
rect 23110 8381 23122 8415
rect 23156 8381 23168 8415
rect 23110 8375 23168 8381
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8381 23351 8415
rect 23293 8375 23351 8381
rect 23523 8415 23581 8421
rect 23523 8381 23535 8415
rect 23569 8412 23581 8415
rect 33410 8412 33416 8424
rect 23569 8384 33416 8412
rect 23569 8381 23581 8384
rect 23523 8375 23581 8381
rect 33410 8372 33416 8384
rect 33468 8372 33474 8424
rect 33686 8412 33692 8424
rect 33647 8384 33692 8412
rect 33686 8372 33692 8384
rect 33744 8372 33750 8424
rect 35437 8415 35495 8421
rect 35437 8412 35449 8415
rect 33796 8384 35449 8412
rect 23382 8344 23388 8356
rect 16540 8316 20116 8344
rect 20364 8316 20576 8344
rect 23343 8316 23388 8344
rect 16540 8304 16546 8316
rect 3694 8236 3700 8288
rect 3752 8276 3758 8288
rect 20364 8276 20392 8316
rect 3752 8248 20392 8276
rect 20548 8276 20576 8316
rect 23382 8304 23388 8316
rect 23440 8304 23446 8356
rect 30282 8304 30288 8356
rect 30340 8344 30346 8356
rect 33796 8344 33824 8384
rect 35437 8381 35449 8384
rect 35483 8381 35495 8415
rect 35437 8375 35495 8381
rect 30340 8316 33824 8344
rect 30340 8304 30346 8316
rect 34422 8304 34428 8356
rect 34480 8344 34486 8356
rect 35253 8347 35311 8353
rect 35253 8344 35265 8347
rect 34480 8316 35265 8344
rect 34480 8304 34486 8316
rect 35253 8313 35265 8316
rect 35299 8313 35311 8347
rect 35544 8344 35572 8452
rect 35710 8412 35716 8424
rect 35671 8384 35716 8412
rect 35710 8372 35716 8384
rect 35768 8372 35774 8424
rect 38746 8372 38752 8424
rect 38804 8412 38810 8424
rect 38949 8421 38977 8452
rect 47486 8440 47492 8452
rect 47544 8440 47550 8492
rect 50522 8440 50528 8492
rect 50580 8480 50586 8492
rect 50580 8452 50844 8480
rect 50580 8440 50586 8452
rect 38841 8415 38899 8421
rect 38841 8412 38853 8415
rect 38804 8384 38853 8412
rect 38804 8372 38810 8384
rect 38841 8381 38853 8384
rect 38887 8381 38899 8415
rect 38841 8375 38899 8381
rect 38934 8415 38992 8421
rect 38934 8381 38946 8415
rect 38980 8381 38992 8415
rect 38934 8375 38992 8381
rect 39022 8372 39028 8424
rect 39080 8412 39086 8424
rect 39390 8421 39396 8424
rect 39209 8415 39267 8421
rect 39209 8412 39221 8415
rect 39080 8384 39221 8412
rect 39080 8372 39086 8384
rect 39209 8381 39221 8384
rect 39255 8381 39267 8415
rect 39347 8415 39396 8421
rect 39347 8412 39359 8415
rect 39303 8384 39359 8412
rect 39209 8375 39267 8381
rect 39347 8381 39359 8384
rect 39393 8381 39396 8415
rect 39347 8375 39396 8381
rect 39390 8372 39396 8375
rect 39448 8412 39454 8424
rect 41506 8412 41512 8424
rect 39448 8384 41512 8412
rect 39448 8372 39454 8384
rect 41506 8372 41512 8384
rect 41564 8372 41570 8424
rect 49234 8412 49240 8424
rect 49195 8384 49240 8412
rect 49234 8372 49240 8384
rect 49292 8372 49298 8424
rect 50430 8372 50436 8424
rect 50488 8412 50494 8424
rect 50697 8415 50755 8421
rect 50697 8412 50709 8415
rect 50488 8384 50709 8412
rect 50488 8372 50494 8384
rect 50697 8381 50709 8384
rect 50743 8381 50755 8415
rect 50816 8412 50844 8452
rect 51074 8440 51080 8492
rect 51132 8440 51138 8492
rect 51184 8480 51212 8520
rect 51534 8508 51540 8560
rect 51592 8548 51598 8560
rect 55582 8548 55588 8560
rect 51592 8520 55588 8548
rect 51592 8508 51598 8520
rect 55582 8508 55588 8520
rect 55640 8508 55646 8560
rect 56502 8508 56508 8560
rect 56560 8548 56566 8560
rect 61105 8551 61163 8557
rect 61105 8548 61117 8551
rect 56560 8520 61117 8548
rect 56560 8508 56566 8520
rect 61105 8517 61117 8520
rect 61151 8517 61163 8551
rect 68094 8548 68100 8560
rect 61105 8511 61163 8517
rect 61672 8520 68100 8548
rect 61672 8480 61700 8520
rect 68094 8508 68100 8520
rect 68152 8508 68158 8560
rect 68278 8508 68284 8560
rect 68336 8548 68342 8560
rect 94455 8551 94513 8557
rect 94455 8548 94467 8551
rect 68336 8520 94467 8548
rect 68336 8508 68342 8520
rect 94455 8517 94467 8520
rect 94501 8517 94513 8551
rect 94455 8511 94513 8517
rect 94608 8480 94636 8579
rect 94866 8548 94872 8560
rect 94700 8520 94872 8548
rect 94700 8489 94728 8520
rect 94866 8508 94872 8520
rect 94924 8508 94930 8560
rect 51184 8452 61700 8480
rect 61764 8452 67588 8480
rect 50985 8415 51043 8421
rect 50985 8412 50997 8415
rect 50816 8384 50997 8412
rect 50697 8375 50755 8381
rect 50985 8381 50997 8384
rect 51031 8381 51043 8415
rect 50985 8375 51043 8381
rect 35621 8347 35679 8353
rect 35621 8344 35633 8347
rect 35544 8316 35633 8344
rect 35253 8307 35311 8313
rect 35621 8313 35633 8316
rect 35667 8313 35679 8347
rect 35621 8307 35679 8313
rect 38654 8304 38660 8356
rect 38712 8344 38718 8356
rect 39117 8347 39175 8353
rect 39117 8344 39129 8347
rect 38712 8316 39129 8344
rect 38712 8304 38718 8316
rect 39117 8313 39129 8316
rect 39163 8313 39175 8347
rect 48498 8344 48504 8356
rect 39117 8307 39175 8313
rect 41386 8316 48504 8344
rect 25958 8276 25964 8288
rect 20548 8248 25964 8276
rect 3752 8236 3758 8248
rect 25958 8236 25964 8248
rect 26016 8236 26022 8288
rect 30926 8236 30932 8288
rect 30984 8276 30990 8288
rect 37550 8276 37556 8288
rect 30984 8248 37556 8276
rect 30984 8236 30990 8248
rect 37550 8236 37556 8248
rect 37608 8236 37614 8288
rect 37642 8236 37648 8288
rect 37700 8276 37706 8288
rect 41386 8276 41414 8316
rect 48498 8304 48504 8316
rect 48556 8304 48562 8356
rect 49326 8304 49332 8356
rect 49384 8344 49390 8356
rect 49970 8344 49976 8356
rect 49384 8316 49976 8344
rect 49384 8304 49390 8316
rect 49970 8304 49976 8316
rect 50028 8304 50034 8356
rect 50525 8347 50583 8353
rect 50525 8313 50537 8347
rect 50571 8344 50583 8347
rect 50798 8344 50804 8356
rect 50571 8316 50804 8344
rect 50571 8313 50583 8316
rect 50525 8307 50583 8313
rect 50798 8304 50804 8316
rect 50856 8304 50862 8356
rect 50893 8347 50951 8353
rect 50893 8313 50905 8347
rect 50939 8344 50951 8347
rect 51092 8344 51120 8440
rect 53834 8372 53840 8424
rect 53892 8412 53898 8424
rect 54297 8415 54355 8421
rect 54297 8412 54309 8415
rect 53892 8384 54309 8412
rect 53892 8372 53898 8384
rect 54297 8381 54309 8384
rect 54343 8381 54355 8415
rect 54297 8375 54355 8381
rect 56597 8415 56655 8421
rect 56597 8381 56609 8415
rect 56643 8412 56655 8415
rect 60826 8412 60832 8424
rect 56643 8384 60832 8412
rect 56643 8381 56655 8384
rect 56597 8375 56655 8381
rect 60826 8372 60832 8384
rect 60884 8372 60890 8424
rect 61105 8415 61163 8421
rect 61105 8381 61117 8415
rect 61151 8412 61163 8415
rect 61289 8415 61347 8421
rect 61289 8412 61301 8415
rect 61151 8384 61301 8412
rect 61151 8381 61163 8384
rect 61105 8375 61163 8381
rect 61289 8381 61301 8384
rect 61335 8412 61347 8415
rect 61654 8412 61660 8424
rect 61335 8384 61660 8412
rect 61335 8381 61347 8384
rect 61289 8375 61347 8381
rect 61654 8372 61660 8384
rect 61712 8372 61718 8424
rect 50939 8316 51120 8344
rect 50939 8313 50951 8316
rect 50893 8307 50951 8313
rect 51166 8304 51172 8356
rect 51224 8344 51230 8356
rect 61764 8344 61792 8452
rect 62206 8372 62212 8424
rect 62264 8412 62270 8424
rect 65518 8412 65524 8424
rect 62264 8384 65524 8412
rect 62264 8372 62270 8384
rect 65518 8372 65524 8384
rect 65576 8372 65582 8424
rect 65978 8412 65984 8424
rect 65939 8384 65984 8412
rect 65978 8372 65984 8384
rect 66036 8412 66042 8424
rect 66162 8412 66168 8424
rect 66036 8384 66168 8412
rect 66036 8372 66042 8384
rect 66162 8372 66168 8384
rect 66220 8372 66226 8424
rect 67450 8412 67456 8424
rect 67411 8384 67456 8412
rect 67450 8372 67456 8384
rect 67508 8372 67514 8424
rect 67560 8412 67588 8452
rect 67836 8452 77294 8480
rect 67836 8412 67864 8452
rect 67560 8384 67864 8412
rect 77266 8412 77294 8452
rect 80026 8452 94636 8480
rect 94685 8483 94743 8489
rect 80026 8412 80054 8452
rect 94685 8449 94697 8483
rect 94731 8449 94743 8483
rect 94685 8443 94743 8449
rect 94777 8483 94835 8489
rect 94777 8449 94789 8483
rect 94823 8449 94835 8483
rect 94777 8443 94835 8449
rect 94792 8412 94820 8443
rect 77266 8384 80054 8412
rect 93826 8384 94820 8412
rect 51224 8316 61792 8344
rect 51224 8304 51230 8316
rect 61838 8304 61844 8356
rect 61896 8344 61902 8356
rect 63862 8344 63868 8356
rect 61896 8316 63868 8344
rect 61896 8304 61902 8316
rect 63862 8304 63868 8316
rect 63920 8304 63926 8356
rect 65242 8304 65248 8356
rect 65300 8344 65306 8356
rect 66070 8344 66076 8356
rect 65300 8316 66076 8344
rect 65300 8304 65306 8316
rect 66070 8304 66076 8316
rect 66128 8344 66134 8356
rect 66349 8347 66407 8353
rect 66349 8344 66361 8347
rect 66128 8316 66361 8344
rect 66128 8304 66134 8316
rect 66349 8313 66361 8316
rect 66395 8313 66407 8347
rect 66349 8307 66407 8313
rect 67269 8347 67327 8353
rect 67269 8313 67281 8347
rect 67315 8344 67327 8347
rect 67821 8347 67879 8353
rect 67821 8344 67833 8347
rect 67315 8316 67833 8344
rect 67315 8313 67327 8316
rect 67269 8307 67327 8313
rect 67821 8313 67833 8316
rect 67867 8313 67879 8347
rect 67821 8307 67879 8313
rect 68094 8304 68100 8356
rect 68152 8344 68158 8356
rect 93826 8344 93854 8384
rect 68152 8316 93854 8344
rect 68152 8304 68158 8316
rect 94130 8304 94136 8356
rect 94188 8344 94194 8356
rect 94317 8347 94375 8353
rect 94317 8344 94329 8347
rect 94188 8316 94329 8344
rect 94188 8304 94194 8316
rect 94317 8313 94329 8316
rect 94363 8313 94375 8347
rect 94317 8307 94375 8313
rect 37700 8248 41414 8276
rect 37700 8236 37706 8248
rect 46198 8236 46204 8288
rect 46256 8276 46262 8288
rect 74074 8276 74080 8288
rect 46256 8248 74080 8276
rect 46256 8236 46262 8248
rect 74074 8236 74080 8248
rect 74132 8236 74138 8288
rect 1104 8186 98808 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 50326 8186
rect 50378 8134 50390 8186
rect 50442 8134 50454 8186
rect 50506 8134 50518 8186
rect 50570 8134 81046 8186
rect 81098 8134 81110 8186
rect 81162 8134 81174 8186
rect 81226 8134 81238 8186
rect 81290 8134 98808 8186
rect 1104 8112 98808 8134
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 33318 8072 33324 8084
rect 10928 8044 33180 8072
rect 33279 8044 33324 8072
rect 10928 8032 10934 8044
rect 9490 8004 9496 8016
rect 1780 7976 9496 8004
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1486 7936 1492 7948
rect 1443 7908 1492 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1486 7896 1492 7908
rect 1544 7896 1550 7948
rect 1780 7945 1808 7976
rect 9490 7964 9496 7976
rect 9548 7964 9554 8016
rect 27338 8004 27344 8016
rect 10980 7976 27344 8004
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7905 1823 7939
rect 2038 7936 2044 7948
rect 1999 7908 2044 7936
rect 1765 7899 1823 7905
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2866 7936 2872 7948
rect 2179 7908 2872 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 10410 7936 10416 7948
rect 10371 7908 10416 7936
rect 10410 7896 10416 7908
rect 10468 7896 10474 7948
rect 10980 7945 11008 7976
rect 27338 7964 27344 7976
rect 27396 7964 27402 8016
rect 33152 8004 33180 8044
rect 33318 8032 33324 8044
rect 33376 8032 33382 8084
rect 33686 8032 33692 8084
rect 33744 8072 33750 8084
rect 37642 8072 37648 8084
rect 33744 8044 37648 8072
rect 33744 8032 33750 8044
rect 37642 8032 37648 8044
rect 37700 8032 37706 8084
rect 40218 8032 40224 8084
rect 40276 8072 40282 8084
rect 46198 8072 46204 8084
rect 40276 8044 46204 8072
rect 40276 8032 40282 8044
rect 46198 8032 46204 8044
rect 46256 8032 46262 8084
rect 46290 8032 46296 8084
rect 46348 8072 46354 8084
rect 46348 8044 46428 8072
rect 46348 8032 46354 8044
rect 38838 8004 38844 8016
rect 33152 7976 38844 8004
rect 38838 7964 38844 7976
rect 38896 7964 38902 8016
rect 40034 8004 40040 8016
rect 39132 7976 40040 8004
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7905 11023 7939
rect 10965 7899 11023 7905
rect 1854 7868 1860 7880
rect 1815 7840 1860 7868
rect 1854 7828 1860 7840
rect 1912 7828 1918 7880
rect 2682 7868 2688 7880
rect 2643 7840 2688 7868
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 10042 7868 10048 7880
rect 10003 7840 10048 7868
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7868 10563 7871
rect 10594 7868 10600 7880
rect 10551 7840 10600 7868
rect 10551 7837 10563 7840
rect 10505 7831 10563 7837
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 10796 7868 10824 7899
rect 25774 7896 25780 7948
rect 25832 7936 25838 7948
rect 31846 7936 31852 7948
rect 25832 7908 31852 7936
rect 25832 7896 25838 7908
rect 31846 7896 31852 7908
rect 31904 7896 31910 7948
rect 31941 7939 31999 7945
rect 31941 7905 31953 7939
rect 31987 7936 31999 7939
rect 32030 7936 32036 7948
rect 31987 7908 32036 7936
rect 31987 7905 31999 7908
rect 31941 7899 31999 7905
rect 32030 7896 32036 7908
rect 32088 7896 32094 7948
rect 32214 7936 32220 7948
rect 32175 7908 32220 7936
rect 32214 7896 32220 7908
rect 32272 7896 32278 7948
rect 37274 7936 37280 7948
rect 37235 7908 37280 7936
rect 37274 7896 37280 7908
rect 37332 7896 37338 7948
rect 37645 7939 37703 7945
rect 37645 7905 37657 7939
rect 37691 7905 37703 7939
rect 38010 7936 38016 7948
rect 37971 7908 38016 7936
rect 37645 7899 37703 7905
rect 32674 7868 32680 7880
rect 10796 7840 32680 7868
rect 9677 7803 9735 7809
rect 9677 7769 9689 7803
rect 9723 7800 9735 7803
rect 10796 7800 10824 7840
rect 32674 7828 32680 7840
rect 32732 7868 32738 7880
rect 33042 7868 33048 7880
rect 32732 7840 33048 7868
rect 32732 7828 32738 7840
rect 33042 7828 33048 7840
rect 33100 7828 33106 7880
rect 37550 7868 37556 7880
rect 37511 7840 37556 7868
rect 37550 7828 37556 7840
rect 37608 7828 37614 7880
rect 9723 7772 10824 7800
rect 37660 7800 37688 7899
rect 38010 7896 38016 7908
rect 38068 7896 38074 7948
rect 39132 7945 39160 7976
rect 40034 7964 40040 7976
rect 40092 7964 40098 8016
rect 39117 7939 39175 7945
rect 39117 7905 39129 7939
rect 39163 7905 39175 7939
rect 39117 7899 39175 7905
rect 39206 7896 39212 7948
rect 39264 7936 39270 7948
rect 39301 7939 39359 7945
rect 39301 7936 39313 7939
rect 39264 7908 39313 7936
rect 39264 7896 39270 7908
rect 39301 7905 39313 7908
rect 39347 7905 39359 7939
rect 39301 7899 39359 7905
rect 39393 7939 39451 7945
rect 39393 7905 39405 7939
rect 39439 7905 39451 7939
rect 39393 7899 39451 7905
rect 38102 7868 38108 7880
rect 38063 7840 38108 7868
rect 38102 7828 38108 7840
rect 38160 7828 38166 7880
rect 38562 7868 38568 7880
rect 38396 7840 38568 7868
rect 38396 7800 38424 7840
rect 38562 7828 38568 7840
rect 38620 7828 38626 7880
rect 38654 7828 38660 7880
rect 38712 7868 38718 7880
rect 39408 7868 39436 7899
rect 39482 7896 39488 7948
rect 39540 7945 39546 7948
rect 39540 7939 39595 7945
rect 39540 7905 39549 7939
rect 39583 7936 39595 7939
rect 46198 7936 46204 7948
rect 39583 7908 46204 7936
rect 39583 7905 39595 7908
rect 39540 7899 39595 7905
rect 39540 7896 39546 7899
rect 46198 7896 46204 7908
rect 46256 7896 46262 7948
rect 46400 7936 46428 8044
rect 49142 8032 49148 8084
rect 49200 8072 49206 8084
rect 87506 8072 87512 8084
rect 49200 8044 87512 8072
rect 49200 8032 49206 8044
rect 87506 8032 87512 8044
rect 87564 8032 87570 8084
rect 47854 7964 47860 8016
rect 47912 8004 47918 8016
rect 90174 8004 90180 8016
rect 47912 7976 90180 8004
rect 47912 7964 47918 7976
rect 90174 7964 90180 7976
rect 90232 7964 90238 8016
rect 81710 7936 81716 7948
rect 46400 7908 81716 7936
rect 81710 7896 81716 7908
rect 81768 7936 81774 7948
rect 81894 7936 81900 7948
rect 81768 7908 81900 7936
rect 81768 7896 81774 7908
rect 81894 7896 81900 7908
rect 81952 7896 81958 7948
rect 83274 7896 83280 7948
rect 83332 7936 83338 7948
rect 94501 7939 94559 7945
rect 94501 7936 94513 7939
rect 83332 7908 94513 7936
rect 83332 7896 83338 7908
rect 94501 7905 94513 7908
rect 94547 7905 94559 7939
rect 94501 7899 94559 7905
rect 38712 7840 39436 7868
rect 39686 7871 39744 7877
rect 38712 7828 38718 7840
rect 39686 7837 39698 7871
rect 39732 7868 39744 7871
rect 46106 7868 46112 7880
rect 39732 7840 46112 7868
rect 39732 7837 39744 7840
rect 39686 7831 39744 7837
rect 46106 7828 46112 7840
rect 46164 7828 46170 7880
rect 46474 7828 46480 7880
rect 46532 7868 46538 7880
rect 67726 7868 67732 7880
rect 46532 7840 67732 7868
rect 46532 7828 46538 7840
rect 67726 7828 67732 7840
rect 67784 7828 67790 7880
rect 73062 7828 73068 7880
rect 73120 7868 73126 7880
rect 94777 7871 94835 7877
rect 94777 7868 94789 7871
rect 73120 7840 94789 7868
rect 73120 7828 73126 7840
rect 94777 7837 94789 7840
rect 94823 7837 94835 7871
rect 94777 7831 94835 7837
rect 37660 7772 38424 7800
rect 38473 7803 38531 7809
rect 9723 7769 9735 7772
rect 9677 7763 9735 7769
rect 38473 7769 38485 7803
rect 38519 7800 38531 7803
rect 91278 7800 91284 7812
rect 38519 7772 91284 7800
rect 38519 7769 38531 7772
rect 38473 7763 38531 7769
rect 91278 7760 91284 7772
rect 91336 7760 91342 7812
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 45370 7732 45376 7744
rect 10100 7704 45376 7732
rect 10100 7692 10106 7704
rect 45370 7692 45376 7704
rect 45428 7692 45434 7744
rect 45554 7692 45560 7744
rect 45612 7732 45618 7744
rect 46474 7732 46480 7744
rect 45612 7704 46480 7732
rect 45612 7692 45618 7704
rect 46474 7692 46480 7704
rect 46532 7692 46538 7744
rect 46566 7692 46572 7744
rect 46624 7732 46630 7744
rect 49694 7732 49700 7744
rect 46624 7704 49700 7732
rect 46624 7692 46630 7704
rect 49694 7692 49700 7704
rect 49752 7692 49758 7744
rect 50154 7692 50160 7744
rect 50212 7732 50218 7744
rect 50706 7732 50712 7744
rect 50212 7704 50712 7732
rect 50212 7692 50218 7704
rect 50706 7692 50712 7704
rect 50764 7692 50770 7744
rect 54662 7692 54668 7744
rect 54720 7732 54726 7744
rect 56226 7732 56232 7744
rect 54720 7704 56232 7732
rect 54720 7692 54726 7704
rect 56226 7692 56232 7704
rect 56284 7692 56290 7744
rect 56870 7692 56876 7744
rect 56928 7732 56934 7744
rect 63954 7732 63960 7744
rect 56928 7704 63960 7732
rect 56928 7692 56934 7704
rect 63954 7692 63960 7704
rect 64012 7692 64018 7744
rect 66990 7692 66996 7744
rect 67048 7732 67054 7744
rect 67266 7732 67272 7744
rect 67048 7704 67272 7732
rect 67048 7692 67054 7704
rect 67266 7692 67272 7704
rect 67324 7692 67330 7744
rect 77386 7692 77392 7744
rect 77444 7732 77450 7744
rect 77754 7732 77760 7744
rect 77444 7704 77760 7732
rect 77444 7692 77450 7704
rect 77754 7692 77760 7704
rect 77812 7692 77818 7744
rect 77846 7692 77852 7744
rect 77904 7732 77910 7744
rect 83366 7732 83372 7744
rect 77904 7704 83372 7732
rect 77904 7692 77910 7704
rect 83366 7692 83372 7704
rect 83424 7692 83430 7744
rect 1104 7642 98808 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 65686 7642
rect 65738 7590 65750 7642
rect 65802 7590 65814 7642
rect 65866 7590 65878 7642
rect 65930 7590 96406 7642
rect 96458 7590 96470 7642
rect 96522 7590 96534 7642
rect 96586 7590 96598 7642
rect 96650 7590 98808 7642
rect 1104 7568 98808 7590
rect 1854 7488 1860 7540
rect 1912 7528 1918 7540
rect 20898 7528 20904 7540
rect 1912 7500 20904 7528
rect 1912 7488 1918 7500
rect 20898 7488 20904 7500
rect 20956 7528 20962 7540
rect 23382 7528 23388 7540
rect 20956 7500 23388 7528
rect 20956 7488 20962 7500
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 25041 7531 25099 7537
rect 25041 7497 25053 7531
rect 25087 7528 25099 7531
rect 26786 7528 26792 7540
rect 25087 7500 26792 7528
rect 25087 7497 25099 7500
rect 25041 7491 25099 7497
rect 26786 7488 26792 7500
rect 26844 7488 26850 7540
rect 31018 7488 31024 7540
rect 31076 7528 31082 7540
rect 31076 7500 53972 7528
rect 31076 7488 31082 7500
rect 11882 7460 11888 7472
rect 11843 7432 11888 7460
rect 11882 7420 11888 7432
rect 11940 7460 11946 7472
rect 12253 7463 12311 7469
rect 12253 7460 12265 7463
rect 11940 7432 12265 7460
rect 11940 7420 11946 7432
rect 12253 7429 12265 7432
rect 12299 7429 12311 7463
rect 12253 7423 12311 7429
rect 16942 7420 16948 7472
rect 17000 7460 17006 7472
rect 17770 7460 17776 7472
rect 17000 7432 17776 7460
rect 17000 7420 17006 7432
rect 17770 7420 17776 7432
rect 17828 7420 17834 7472
rect 24949 7463 25007 7469
rect 24949 7429 24961 7463
rect 24995 7460 25007 7463
rect 25774 7460 25780 7472
rect 24995 7432 25780 7460
rect 24995 7429 25007 7432
rect 24949 7423 25007 7429
rect 25774 7420 25780 7432
rect 25832 7420 25838 7472
rect 27157 7463 27215 7469
rect 27157 7429 27169 7463
rect 27203 7460 27215 7463
rect 32582 7460 32588 7472
rect 27203 7432 32588 7460
rect 27203 7429 27215 7432
rect 27157 7423 27215 7429
rect 32582 7420 32588 7432
rect 32640 7420 32646 7472
rect 34698 7460 34704 7472
rect 33244 7432 34704 7460
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 9585 7395 9643 7401
rect 2924 7364 9260 7392
rect 2924 7352 2930 7364
rect 1486 7284 1492 7336
rect 1544 7324 1550 7336
rect 9122 7324 9128 7336
rect 1544 7296 9128 7324
rect 1544 7284 1550 7296
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9232 7256 9260 7364
rect 9585 7361 9597 7395
rect 9631 7392 9643 7395
rect 19334 7392 19340 7404
rect 9631 7364 19340 7392
rect 9631 7361 9643 7364
rect 9585 7355 9643 7361
rect 19334 7352 19340 7364
rect 19392 7352 19398 7404
rect 22922 7352 22928 7404
rect 22980 7392 22986 7404
rect 25409 7395 25467 7401
rect 25409 7392 25421 7395
rect 22980 7364 25421 7392
rect 22980 7352 22986 7364
rect 25409 7361 25421 7364
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 25501 7395 25559 7401
rect 25501 7361 25513 7395
rect 25547 7392 25559 7395
rect 33244 7392 33272 7432
rect 34698 7420 34704 7432
rect 34756 7420 34762 7472
rect 37274 7420 37280 7472
rect 37332 7460 37338 7472
rect 45278 7460 45284 7472
rect 37332 7432 45284 7460
rect 37332 7420 37338 7432
rect 45278 7420 45284 7432
rect 45336 7420 45342 7472
rect 45462 7420 45468 7472
rect 45520 7460 45526 7472
rect 49602 7460 49608 7472
rect 45520 7432 49608 7460
rect 45520 7420 45526 7432
rect 49602 7420 49608 7432
rect 49660 7420 49666 7472
rect 49694 7420 49700 7472
rect 49752 7460 49758 7472
rect 53944 7460 53972 7500
rect 54018 7488 54024 7540
rect 54076 7528 54082 7540
rect 54386 7528 54392 7540
rect 54076 7500 54392 7528
rect 54076 7488 54082 7500
rect 54386 7488 54392 7500
rect 54444 7488 54450 7540
rect 60182 7488 60188 7540
rect 60240 7528 60246 7540
rect 65334 7528 65340 7540
rect 60240 7500 65340 7528
rect 60240 7488 60246 7500
rect 65334 7488 65340 7500
rect 65392 7488 65398 7540
rect 69566 7528 69572 7540
rect 69527 7500 69572 7528
rect 69566 7488 69572 7500
rect 69624 7528 69630 7540
rect 69937 7531 69995 7537
rect 69937 7528 69949 7531
rect 69624 7500 69949 7528
rect 69624 7488 69630 7500
rect 69937 7497 69949 7500
rect 69983 7497 69995 7531
rect 78674 7528 78680 7540
rect 69937 7491 69995 7497
rect 70366 7500 78680 7528
rect 57698 7460 57704 7472
rect 49752 7432 53880 7460
rect 53944 7432 57704 7460
rect 49752 7420 49758 7432
rect 25547 7364 33272 7392
rect 25547 7361 25559 7364
rect 25501 7355 25559 7361
rect 9490 7324 9496 7336
rect 9451 7296 9496 7324
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 9861 7327 9919 7333
rect 9861 7293 9873 7327
rect 9907 7293 9919 7327
rect 10042 7324 10048 7336
rect 10003 7296 10048 7324
rect 9861 7287 9919 7293
rect 9876 7256 9904 7287
rect 10042 7284 10048 7296
rect 10100 7284 10106 7336
rect 20622 7284 20628 7336
rect 20680 7324 20686 7336
rect 24854 7324 24860 7336
rect 20680 7296 24860 7324
rect 20680 7284 20686 7296
rect 24854 7284 24860 7296
rect 24912 7284 24918 7336
rect 25225 7327 25283 7333
rect 25225 7293 25237 7327
rect 25271 7324 25283 7327
rect 25314 7324 25320 7336
rect 25271 7296 25320 7324
rect 25271 7293 25283 7296
rect 25225 7287 25283 7293
rect 25314 7284 25320 7296
rect 25372 7284 25378 7336
rect 9232 7228 9904 7256
rect 10413 7259 10471 7265
rect 10413 7225 10425 7259
rect 10459 7256 10471 7259
rect 24118 7256 24124 7268
rect 10459 7228 24124 7256
rect 10459 7225 10471 7228
rect 10413 7219 10471 7225
rect 24118 7216 24124 7228
rect 24176 7216 24182 7268
rect 25424 7256 25452 7355
rect 34238 7352 34244 7404
rect 34296 7392 34302 7404
rect 39022 7392 39028 7404
rect 34296 7364 39028 7392
rect 34296 7352 34302 7364
rect 39022 7352 39028 7364
rect 39080 7352 39086 7404
rect 39298 7352 39304 7404
rect 39356 7392 39362 7404
rect 39850 7392 39856 7404
rect 39356 7364 39856 7392
rect 39356 7352 39362 7364
rect 39850 7352 39856 7364
rect 39908 7352 39914 7404
rect 40034 7352 40040 7404
rect 40092 7392 40098 7404
rect 40954 7392 40960 7404
rect 40092 7364 40960 7392
rect 40092 7352 40098 7364
rect 40954 7352 40960 7364
rect 41012 7392 41018 7404
rect 53650 7392 53656 7404
rect 41012 7364 53656 7392
rect 41012 7352 41018 7364
rect 53650 7352 53656 7364
rect 53708 7352 53714 7404
rect 25593 7327 25651 7333
rect 25593 7293 25605 7327
rect 25639 7324 25651 7327
rect 25682 7324 25688 7336
rect 25639 7296 25688 7324
rect 25639 7293 25651 7296
rect 25593 7287 25651 7293
rect 25682 7284 25688 7296
rect 25740 7284 25746 7336
rect 25774 7284 25780 7336
rect 25832 7324 25838 7336
rect 25958 7324 25964 7336
rect 25832 7296 25877 7324
rect 25919 7296 25964 7324
rect 25832 7284 25838 7296
rect 25958 7284 25964 7296
rect 26016 7284 26022 7336
rect 26602 7284 26608 7336
rect 26660 7324 26666 7336
rect 26660 7296 31754 7324
rect 26660 7284 26666 7296
rect 27157 7259 27215 7265
rect 27157 7256 27169 7259
rect 25424 7228 27169 7256
rect 27157 7225 27169 7228
rect 27203 7225 27215 7259
rect 31726 7256 31754 7296
rect 31846 7284 31852 7336
rect 31904 7324 31910 7336
rect 38286 7324 38292 7336
rect 31904 7296 38292 7324
rect 31904 7284 31910 7296
rect 38286 7284 38292 7296
rect 38344 7324 38350 7336
rect 38470 7324 38476 7336
rect 38344 7296 38476 7324
rect 38344 7284 38350 7296
rect 38470 7284 38476 7296
rect 38528 7284 38534 7336
rect 38565 7327 38623 7333
rect 38565 7293 38577 7327
rect 38611 7324 38623 7327
rect 42702 7324 42708 7336
rect 38611 7296 42708 7324
rect 38611 7293 38623 7296
rect 38565 7287 38623 7293
rect 42702 7284 42708 7296
rect 42760 7284 42766 7336
rect 46566 7324 46572 7336
rect 46124 7296 46572 7324
rect 38654 7256 38660 7268
rect 31726 7228 38660 7256
rect 27157 7219 27215 7225
rect 38654 7216 38660 7228
rect 38712 7216 38718 7268
rect 38746 7216 38752 7268
rect 38804 7256 38810 7268
rect 46124 7256 46152 7296
rect 46566 7284 46572 7296
rect 46624 7284 46630 7336
rect 49050 7284 49056 7336
rect 49108 7324 49114 7336
rect 49226 7327 49284 7333
rect 49226 7324 49238 7327
rect 49108 7296 49238 7324
rect 49108 7284 49114 7296
rect 49226 7293 49238 7296
rect 49272 7293 49284 7327
rect 49418 7324 49424 7336
rect 49379 7296 49424 7324
rect 49226 7287 49284 7293
rect 49418 7284 49424 7296
rect 49476 7284 49482 7336
rect 49602 7284 49608 7336
rect 49660 7324 49666 7336
rect 50062 7333 50068 7336
rect 49881 7327 49939 7333
rect 49660 7296 49705 7324
rect 49660 7284 49666 7296
rect 49881 7293 49893 7327
rect 49927 7293 49939 7327
rect 49881 7287 49939 7293
rect 50019 7327 50068 7333
rect 50019 7293 50031 7327
rect 50065 7293 50068 7327
rect 50019 7287 50068 7293
rect 48866 7256 48872 7268
rect 38804 7228 46152 7256
rect 46216 7228 48872 7256
rect 38804 7216 38810 7228
rect 18046 7148 18052 7200
rect 18104 7188 18110 7200
rect 20162 7188 20168 7200
rect 18104 7160 20168 7188
rect 18104 7148 18110 7160
rect 20162 7148 20168 7160
rect 20220 7148 20226 7200
rect 25958 7148 25964 7200
rect 26016 7188 26022 7200
rect 46216 7188 46244 7228
rect 48866 7216 48872 7228
rect 48924 7216 48930 7268
rect 26016 7160 46244 7188
rect 26016 7148 26022 7160
rect 46290 7148 46296 7200
rect 46348 7188 46354 7200
rect 48958 7188 48964 7200
rect 46348 7160 48964 7188
rect 46348 7148 46354 7160
rect 48958 7148 48964 7160
rect 49016 7148 49022 7200
rect 49694 7148 49700 7200
rect 49752 7188 49758 7200
rect 49896 7188 49924 7287
rect 50062 7284 50068 7287
rect 50120 7284 50126 7336
rect 50525 7327 50583 7333
rect 50525 7293 50537 7327
rect 50571 7324 50583 7327
rect 53852 7324 53880 7432
rect 57698 7420 57704 7432
rect 57756 7420 57762 7472
rect 58894 7420 58900 7472
rect 58952 7460 58958 7472
rect 62942 7460 62948 7472
rect 58952 7432 62948 7460
rect 58952 7420 58958 7432
rect 62942 7420 62948 7432
rect 63000 7420 63006 7472
rect 64782 7420 64788 7472
rect 64840 7460 64846 7472
rect 64966 7460 64972 7472
rect 64840 7432 64972 7460
rect 64840 7420 64846 7432
rect 64966 7420 64972 7432
rect 65024 7420 65030 7472
rect 61562 7352 61568 7404
rect 61620 7392 61626 7404
rect 69474 7392 69480 7404
rect 61620 7364 69480 7392
rect 61620 7352 61626 7364
rect 69474 7352 69480 7364
rect 69532 7352 69538 7404
rect 61838 7324 61844 7336
rect 50571 7296 51074 7324
rect 53852 7296 61844 7324
rect 50571 7293 50583 7296
rect 50525 7287 50583 7293
rect 51046 7256 51074 7296
rect 61838 7284 61844 7296
rect 61896 7324 61902 7336
rect 70366 7324 70394 7500
rect 78674 7488 78680 7500
rect 78732 7488 78738 7540
rect 71222 7420 71228 7472
rect 71280 7460 71286 7472
rect 77846 7460 77852 7472
rect 71280 7432 77852 7460
rect 71280 7420 71286 7432
rect 77846 7420 77852 7432
rect 77904 7420 77910 7472
rect 82446 7420 82452 7472
rect 82504 7460 82510 7472
rect 87230 7460 87236 7472
rect 82504 7432 87236 7460
rect 82504 7420 82510 7432
rect 87230 7420 87236 7432
rect 87288 7420 87294 7472
rect 87046 7392 87052 7404
rect 87007 7364 87052 7392
rect 87046 7352 87052 7364
rect 87104 7352 87110 7404
rect 61896 7296 70394 7324
rect 61896 7284 61902 7296
rect 84194 7284 84200 7336
rect 84252 7324 84258 7336
rect 86865 7327 86923 7333
rect 86865 7324 86877 7327
rect 84252 7296 86877 7324
rect 84252 7284 84258 7296
rect 86865 7293 86877 7296
rect 86911 7293 86923 7327
rect 86865 7287 86923 7293
rect 97718 7284 97724 7336
rect 97776 7324 97782 7336
rect 97905 7327 97963 7333
rect 97905 7324 97917 7327
rect 97776 7296 97917 7324
rect 97776 7284 97782 7296
rect 97905 7293 97917 7296
rect 97951 7293 97963 7327
rect 97905 7287 97963 7293
rect 86678 7256 86684 7268
rect 51046 7228 86684 7256
rect 86678 7216 86684 7228
rect 86736 7216 86742 7268
rect 49752 7160 49924 7188
rect 49752 7148 49758 7160
rect 50154 7148 50160 7200
rect 50212 7188 50218 7200
rect 59906 7188 59912 7200
rect 50212 7160 59912 7188
rect 50212 7148 50218 7160
rect 59906 7148 59912 7160
rect 59964 7148 59970 7200
rect 77938 7148 77944 7200
rect 77996 7188 78002 7200
rect 83918 7188 83924 7200
rect 77996 7160 83924 7188
rect 77996 7148 78002 7160
rect 83918 7148 83924 7160
rect 83976 7148 83982 7200
rect 1104 7098 98808 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 50326 7098
rect 50378 7046 50390 7098
rect 50442 7046 50454 7098
rect 50506 7046 50518 7098
rect 50570 7046 81046 7098
rect 81098 7046 81110 7098
rect 81162 7046 81174 7098
rect 81226 7046 81238 7098
rect 81290 7046 98808 7098
rect 1104 7024 98808 7046
rect 3142 6944 3148 6996
rect 3200 6984 3206 6996
rect 3200 6956 6914 6984
rect 3200 6944 3206 6956
rect 6886 6916 6914 6956
rect 19334 6944 19340 6996
rect 19392 6984 19398 6996
rect 20438 6984 20444 6996
rect 19392 6956 20444 6984
rect 19392 6944 19398 6956
rect 20438 6944 20444 6956
rect 20496 6984 20502 6996
rect 34238 6984 34244 6996
rect 20496 6956 34244 6984
rect 20496 6944 20502 6956
rect 34238 6944 34244 6956
rect 34296 6944 34302 6996
rect 39206 6984 39212 6996
rect 34348 6956 39212 6984
rect 34348 6916 34376 6956
rect 39206 6944 39212 6956
rect 39264 6944 39270 6996
rect 46014 6984 46020 6996
rect 41386 6956 46020 6984
rect 5184 6888 5856 6916
rect 6886 6888 34376 6916
rect 4893 6851 4951 6857
rect 4893 6817 4905 6851
rect 4939 6848 4951 6851
rect 5184 6848 5212 6888
rect 4939 6820 5212 6848
rect 5261 6851 5319 6857
rect 4939 6817 4951 6820
rect 4893 6811 4951 6817
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5626 6848 5632 6860
rect 5307 6820 5396 6848
rect 5587 6820 5632 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 5368 6792 5396 6820
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5828 6848 5856 6888
rect 34422 6876 34428 6928
rect 34480 6916 34486 6928
rect 41386 6916 41414 6956
rect 46014 6944 46020 6956
rect 46072 6944 46078 6996
rect 46106 6944 46112 6996
rect 46164 6984 46170 6996
rect 68186 6984 68192 6996
rect 46164 6956 68192 6984
rect 46164 6944 46170 6956
rect 68186 6944 68192 6956
rect 68244 6944 68250 6996
rect 34480 6888 41414 6916
rect 34480 6876 34486 6888
rect 42150 6876 42156 6928
rect 42208 6916 42214 6928
rect 45094 6916 45100 6928
rect 42208 6888 45100 6916
rect 42208 6876 42214 6888
rect 45094 6876 45100 6888
rect 45152 6876 45158 6928
rect 45370 6876 45376 6928
rect 45428 6916 45434 6928
rect 49326 6916 49332 6928
rect 45428 6888 49332 6916
rect 45428 6876 45434 6888
rect 49326 6876 49332 6888
rect 49384 6876 49390 6928
rect 49694 6876 49700 6928
rect 49752 6916 49758 6928
rect 54754 6916 54760 6928
rect 49752 6888 54760 6916
rect 49752 6876 49758 6888
rect 54754 6876 54760 6888
rect 54812 6876 54818 6928
rect 72142 6876 72148 6928
rect 72200 6916 72206 6928
rect 72200 6888 72924 6916
rect 72200 6876 72206 6888
rect 10962 6848 10968 6860
rect 5828 6820 10968 6848
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 19426 6808 19432 6860
rect 19484 6848 19490 6860
rect 43346 6848 43352 6860
rect 19484 6820 41414 6848
rect 43307 6820 43352 6848
rect 19484 6808 19490 6820
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5000 6712 5028 6743
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 6454 6780 6460 6792
rect 5491 6752 6460 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 33870 6780 33876 6792
rect 6564 6752 33876 6780
rect 6564 6712 6592 6752
rect 33870 6740 33876 6752
rect 33928 6740 33934 6792
rect 35434 6740 35440 6792
rect 35492 6780 35498 6792
rect 36906 6780 36912 6792
rect 35492 6752 36912 6780
rect 35492 6740 35498 6752
rect 36906 6740 36912 6752
rect 36964 6740 36970 6792
rect 41386 6780 41414 6820
rect 43346 6808 43352 6820
rect 43404 6808 43410 6860
rect 48590 6808 48596 6860
rect 48648 6848 48654 6860
rect 48648 6820 50108 6848
rect 48648 6808 48654 6820
rect 49970 6780 49976 6792
rect 41386 6752 49976 6780
rect 49970 6740 49976 6752
rect 50028 6740 50034 6792
rect 50080 6780 50108 6820
rect 50706 6808 50712 6860
rect 50764 6848 50770 6860
rect 62209 6851 62267 6857
rect 62209 6848 62221 6851
rect 50764 6820 62221 6848
rect 50764 6808 50770 6820
rect 62209 6817 62221 6820
rect 62255 6817 62267 6851
rect 63586 6848 63592 6860
rect 63547 6820 63592 6848
rect 62209 6811 62267 6817
rect 63586 6808 63592 6820
rect 63644 6808 63650 6860
rect 71958 6808 71964 6860
rect 72016 6848 72022 6860
rect 72421 6851 72479 6857
rect 72421 6848 72433 6851
rect 72016 6820 72433 6848
rect 72016 6808 72022 6820
rect 72421 6817 72433 6820
rect 72467 6817 72479 6851
rect 72602 6848 72608 6860
rect 72563 6820 72608 6848
rect 72421 6811 72479 6817
rect 72602 6808 72608 6820
rect 72660 6808 72666 6860
rect 72896 6857 72924 6888
rect 72789 6851 72847 6857
rect 72789 6817 72801 6851
rect 72835 6817 72847 6851
rect 72789 6811 72847 6817
rect 72881 6851 72939 6857
rect 72881 6817 72893 6851
rect 72927 6817 72939 6851
rect 72881 6811 72939 6817
rect 55674 6780 55680 6792
rect 50080 6752 55680 6780
rect 55674 6740 55680 6752
rect 55732 6740 55738 6792
rect 61746 6740 61752 6792
rect 61804 6780 61810 6792
rect 61933 6783 61991 6789
rect 61933 6780 61945 6783
rect 61804 6752 61945 6780
rect 61804 6740 61810 6752
rect 61933 6749 61945 6752
rect 61979 6749 61991 6783
rect 61933 6743 61991 6749
rect 68462 6740 68468 6792
rect 68520 6780 68526 6792
rect 72804 6780 72832 6811
rect 78398 6808 78404 6860
rect 78456 6848 78462 6860
rect 91462 6848 91468 6860
rect 78456 6820 91468 6848
rect 78456 6808 78462 6820
rect 91462 6808 91468 6820
rect 91520 6808 91526 6860
rect 97537 6851 97595 6857
rect 97537 6817 97549 6851
rect 97583 6848 97595 6851
rect 98270 6848 98276 6860
rect 97583 6820 98276 6848
rect 97583 6817 97595 6820
rect 97537 6811 97595 6817
rect 98270 6808 98276 6820
rect 98328 6808 98334 6860
rect 68520 6752 72832 6780
rect 68520 6740 68526 6752
rect 80514 6740 80520 6792
rect 80572 6780 80578 6792
rect 95878 6780 95884 6792
rect 80572 6752 95884 6780
rect 80572 6740 80578 6752
rect 95878 6740 95884 6752
rect 95936 6740 95942 6792
rect 5000 6684 6592 6712
rect 7466 6672 7472 6724
rect 7524 6712 7530 6724
rect 56594 6712 56600 6724
rect 7524 6684 56600 6712
rect 7524 6672 7530 6684
rect 56594 6672 56600 6684
rect 56652 6672 56658 6724
rect 83182 6712 83188 6724
rect 63236 6684 83188 6712
rect 3513 6647 3571 6653
rect 3513 6613 3525 6647
rect 3559 6644 3571 6647
rect 3697 6647 3755 6653
rect 3697 6644 3709 6647
rect 3559 6616 3709 6644
rect 3559 6613 3571 6616
rect 3513 6607 3571 6613
rect 3697 6613 3709 6616
rect 3743 6644 3755 6647
rect 3973 6647 4031 6653
rect 3973 6644 3985 6647
rect 3743 6616 3985 6644
rect 3743 6613 3755 6616
rect 3697 6607 3755 6613
rect 3973 6613 3985 6616
rect 4019 6644 4031 6647
rect 4157 6647 4215 6653
rect 4157 6644 4169 6647
rect 4019 6616 4169 6644
rect 4019 6613 4031 6616
rect 3973 6607 4031 6613
rect 4157 6613 4169 6616
rect 4203 6644 4215 6647
rect 4433 6647 4491 6653
rect 4433 6644 4445 6647
rect 4203 6616 4445 6644
rect 4203 6613 4215 6616
rect 4157 6607 4215 6613
rect 4433 6613 4445 6616
rect 4479 6644 4491 6647
rect 5813 6647 5871 6653
rect 5813 6644 5825 6647
rect 4479 6616 5825 6644
rect 4479 6613 4491 6616
rect 4433 6607 4491 6613
rect 5813 6613 5825 6616
rect 5859 6644 5871 6647
rect 5997 6647 6055 6653
rect 5997 6644 6009 6647
rect 5859 6616 6009 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 5997 6613 6009 6616
rect 6043 6644 6055 6647
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 6043 6616 6193 6644
rect 6043 6613 6055 6616
rect 5997 6607 6055 6613
rect 6181 6613 6193 6616
rect 6227 6644 6239 6647
rect 6365 6647 6423 6653
rect 6365 6644 6377 6647
rect 6227 6616 6377 6644
rect 6227 6613 6239 6616
rect 6181 6607 6239 6613
rect 6365 6613 6377 6616
rect 6411 6644 6423 6647
rect 6454 6644 6460 6656
rect 6411 6616 6460 6644
rect 6411 6613 6423 6616
rect 6365 6607 6423 6613
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 6546 6604 6552 6656
rect 6604 6644 6610 6656
rect 6604 6616 6649 6644
rect 6604 6604 6610 6616
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 21910 6644 21916 6656
rect 7800 6616 21916 6644
rect 7800 6604 7806 6616
rect 21910 6604 21916 6616
rect 21968 6604 21974 6656
rect 22002 6604 22008 6656
rect 22060 6644 22066 6656
rect 28350 6644 28356 6656
rect 22060 6616 28356 6644
rect 22060 6604 22066 6616
rect 28350 6604 28356 6616
rect 28408 6644 28414 6656
rect 44818 6644 44824 6656
rect 28408 6616 44824 6644
rect 28408 6604 28414 6616
rect 44818 6604 44824 6616
rect 44876 6644 44882 6656
rect 45462 6644 45468 6656
rect 44876 6616 45468 6644
rect 44876 6604 44882 6616
rect 45462 6604 45468 6616
rect 45520 6604 45526 6656
rect 50798 6604 50804 6656
rect 50856 6644 50862 6656
rect 63236 6644 63264 6684
rect 83182 6672 83188 6684
rect 83240 6672 83246 6724
rect 50856 6616 63264 6644
rect 50856 6604 50862 6616
rect 65978 6604 65984 6656
rect 66036 6644 66042 6656
rect 72602 6644 72608 6656
rect 66036 6616 72608 6644
rect 66036 6604 66042 6616
rect 72602 6604 72608 6616
rect 72660 6604 72666 6656
rect 81342 6604 81348 6656
rect 81400 6644 81406 6656
rect 87598 6644 87604 6656
rect 81400 6616 87604 6644
rect 81400 6604 81406 6616
rect 87598 6604 87604 6616
rect 87656 6604 87662 6656
rect 1104 6554 98808 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 65686 6554
rect 65738 6502 65750 6554
rect 65802 6502 65814 6554
rect 65866 6502 65878 6554
rect 65930 6502 96406 6554
rect 96458 6502 96470 6554
rect 96522 6502 96534 6554
rect 96586 6502 96598 6554
rect 96650 6502 98808 6554
rect 1104 6480 98808 6502
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 72878 6440 72884 6452
rect 8444 6412 72884 6440
rect 8444 6400 8450 6412
rect 72878 6400 72884 6412
rect 72936 6400 72942 6452
rect 78306 6400 78312 6452
rect 78364 6440 78370 6452
rect 82081 6443 82139 6449
rect 82081 6440 82093 6443
rect 78364 6412 82093 6440
rect 78364 6400 78370 6412
rect 82081 6409 82093 6412
rect 82127 6409 82139 6443
rect 82081 6403 82139 6409
rect 93486 6400 93492 6452
rect 93544 6440 93550 6452
rect 96065 6443 96123 6449
rect 96065 6440 96077 6443
rect 93544 6412 96077 6440
rect 93544 6400 93550 6412
rect 96065 6409 96077 6412
rect 96111 6440 96123 6443
rect 96249 6443 96307 6449
rect 96249 6440 96261 6443
rect 96111 6412 96261 6440
rect 96111 6409 96123 6412
rect 96065 6403 96123 6409
rect 96249 6409 96261 6412
rect 96295 6409 96307 6443
rect 96249 6403 96307 6409
rect 7190 6332 7196 6384
rect 7248 6372 7254 6384
rect 8202 6372 8208 6384
rect 7248 6344 8208 6372
rect 7248 6332 7254 6344
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 9122 6332 9128 6384
rect 9180 6372 9186 6384
rect 15194 6372 15200 6384
rect 9180 6344 15200 6372
rect 9180 6332 9186 6344
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 15304 6344 15700 6372
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 11514 6304 11520 6316
rect 5408 6276 11520 6304
rect 5408 6264 5414 6276
rect 11514 6264 11520 6276
rect 11572 6264 11578 6316
rect 15304 6304 15332 6344
rect 15470 6304 15476 6316
rect 11624 6276 15332 6304
rect 15431 6276 15476 6304
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6236 3387 6239
rect 3510 6236 3516 6248
rect 3375 6208 3516 6236
rect 3375 6205 3387 6208
rect 3329 6199 3387 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 4341 6239 4399 6245
rect 4341 6236 4353 6239
rect 4028 6208 4353 6236
rect 4028 6196 4034 6208
rect 4341 6205 4353 6208
rect 4387 6205 4399 6239
rect 4341 6199 4399 6205
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 10226 6236 10232 6248
rect 6604 6208 10232 6236
rect 6604 6196 6610 6208
rect 10226 6196 10232 6208
rect 10284 6236 10290 6248
rect 11624 6236 11652 6276
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 15672 6304 15700 6344
rect 15746 6332 15752 6384
rect 15804 6372 15810 6384
rect 15841 6375 15899 6381
rect 15841 6372 15853 6375
rect 15804 6344 15853 6372
rect 15804 6332 15810 6344
rect 15841 6341 15853 6344
rect 15887 6341 15899 6375
rect 21082 6372 21088 6384
rect 21043 6344 21088 6372
rect 15841 6335 15899 6341
rect 21082 6332 21088 6344
rect 21140 6332 21146 6384
rect 21223 6375 21281 6381
rect 21223 6341 21235 6375
rect 21269 6372 21281 6375
rect 21818 6372 21824 6384
rect 21269 6344 21824 6372
rect 21269 6341 21281 6344
rect 21223 6335 21281 6341
rect 21818 6332 21824 6344
rect 21876 6332 21882 6384
rect 21910 6332 21916 6384
rect 21968 6372 21974 6384
rect 48406 6372 48412 6384
rect 21968 6344 48412 6372
rect 21968 6332 21974 6344
rect 48406 6332 48412 6344
rect 48464 6332 48470 6384
rect 51442 6372 51448 6384
rect 51403 6344 51448 6372
rect 51442 6332 51448 6344
rect 51500 6332 51506 6384
rect 53024 6344 57974 6372
rect 53024 6304 53052 6344
rect 15672 6276 53052 6304
rect 57946 6304 57974 6344
rect 62022 6332 62028 6384
rect 62080 6372 62086 6384
rect 94406 6372 94412 6384
rect 62080 6344 94412 6372
rect 62080 6332 62086 6344
rect 94406 6332 94412 6344
rect 94464 6332 94470 6384
rect 81342 6304 81348 6316
rect 57946 6276 81348 6304
rect 81342 6264 81348 6276
rect 81400 6264 81406 6316
rect 84194 6304 84200 6316
rect 81544 6276 84200 6304
rect 10284 6208 11652 6236
rect 10284 6196 10290 6208
rect 14182 6196 14188 6248
rect 14240 6236 14246 6248
rect 15105 6239 15163 6245
rect 15105 6236 15117 6239
rect 14240 6208 15117 6236
rect 14240 6196 14246 6208
rect 15105 6205 15117 6208
rect 15151 6205 15163 6239
rect 15286 6236 15292 6248
rect 15247 6208 15292 6236
rect 15105 6199 15163 6205
rect 15286 6196 15292 6208
rect 15344 6196 15350 6248
rect 15378 6196 15384 6248
rect 15436 6236 15442 6248
rect 15657 6239 15715 6245
rect 15436 6208 15481 6236
rect 15436 6196 15442 6208
rect 15657 6205 15669 6239
rect 15703 6236 15715 6239
rect 20346 6236 20352 6248
rect 15703 6208 20352 6236
rect 15703 6205 15715 6208
rect 15657 6199 15715 6205
rect 20346 6196 20352 6208
rect 20404 6196 20410 6248
rect 21022 6239 21080 6245
rect 21022 6236 21034 6239
rect 20916 6208 21034 6236
rect 7926 6128 7932 6180
rect 7984 6168 7990 6180
rect 11882 6168 11888 6180
rect 7984 6140 11888 6168
rect 7984 6128 7990 6140
rect 11882 6128 11888 6140
rect 11940 6128 11946 6180
rect 13538 6128 13544 6180
rect 13596 6168 13602 6180
rect 15013 6171 15071 6177
rect 15013 6168 15025 6171
rect 13596 6140 15025 6168
rect 13596 6128 13602 6140
rect 15013 6137 15025 6140
rect 15059 6168 15071 6171
rect 15304 6168 15332 6196
rect 15059 6140 15332 6168
rect 15059 6137 15071 6140
rect 15013 6131 15071 6137
rect 15470 6128 15476 6180
rect 15528 6168 15534 6180
rect 18414 6168 18420 6180
rect 15528 6140 18420 6168
rect 15528 6128 15534 6140
rect 18414 6128 18420 6140
rect 18472 6128 18478 6180
rect 20916 6168 20944 6208
rect 21022 6205 21034 6208
rect 21068 6205 21080 6239
rect 21022 6199 21080 6205
rect 21818 6196 21824 6248
rect 21876 6236 21882 6248
rect 28994 6236 29000 6248
rect 21876 6208 29000 6236
rect 21876 6196 21882 6208
rect 28994 6196 29000 6208
rect 29052 6236 29058 6248
rect 29270 6236 29276 6248
rect 29052 6208 29276 6236
rect 29052 6196 29058 6208
rect 29270 6196 29276 6208
rect 29328 6196 29334 6248
rect 33137 6239 33195 6245
rect 33137 6205 33149 6239
rect 33183 6236 33195 6239
rect 33183 6208 34376 6236
rect 33183 6205 33195 6208
rect 33137 6199 33195 6205
rect 21358 6168 21364 6180
rect 20548 6140 20944 6168
rect 21319 6140 21364 6168
rect 7650 6060 7656 6112
rect 7708 6100 7714 6112
rect 11606 6100 11612 6112
rect 7708 6072 11612 6100
rect 7708 6060 7714 6072
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 15102 6060 15108 6112
rect 15160 6100 15166 6112
rect 17310 6100 17316 6112
rect 15160 6072 17316 6100
rect 15160 6060 15166 6072
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 20254 6060 20260 6112
rect 20312 6100 20318 6112
rect 20548 6109 20576 6140
rect 21358 6128 21364 6140
rect 21416 6128 21422 6180
rect 21634 6128 21640 6180
rect 21692 6168 21698 6180
rect 33689 6171 33747 6177
rect 33689 6168 33701 6171
rect 21692 6140 33701 6168
rect 21692 6128 21698 6140
rect 33689 6137 33701 6140
rect 33735 6168 33747 6171
rect 33870 6168 33876 6180
rect 33735 6140 33876 6168
rect 33735 6137 33747 6140
rect 33689 6131 33747 6137
rect 33870 6128 33876 6140
rect 33928 6128 33934 6180
rect 34348 6168 34376 6208
rect 34422 6196 34428 6248
rect 34480 6236 34486 6248
rect 34480 6208 34525 6236
rect 34480 6196 34486 6208
rect 42794 6196 42800 6248
rect 42852 6236 42858 6248
rect 43806 6236 43812 6248
rect 42852 6208 43812 6236
rect 42852 6196 42858 6208
rect 43806 6196 43812 6208
rect 43864 6196 43870 6248
rect 51261 6239 51319 6245
rect 51261 6205 51273 6239
rect 51307 6236 51319 6239
rect 52730 6236 52736 6248
rect 51307 6208 52736 6236
rect 51307 6205 51319 6208
rect 51261 6199 51319 6205
rect 52730 6196 52736 6208
rect 52788 6196 52794 6248
rect 53002 6239 53060 6245
rect 53002 6205 53014 6239
rect 53048 6205 53060 6239
rect 53002 6199 53060 6205
rect 51994 6168 52000 6180
rect 34348 6140 52000 6168
rect 51994 6128 52000 6140
rect 52052 6128 52058 6180
rect 20533 6103 20591 6109
rect 20533 6100 20545 6103
rect 20312 6072 20545 6100
rect 20312 6060 20318 6072
rect 20533 6069 20545 6072
rect 20579 6069 20591 6103
rect 20714 6100 20720 6112
rect 20675 6072 20720 6100
rect 20533 6063 20591 6069
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 20806 6060 20812 6112
rect 20864 6100 20870 6112
rect 42794 6100 42800 6112
rect 20864 6072 42800 6100
rect 20864 6060 20870 6072
rect 42794 6060 42800 6072
rect 42852 6060 42858 6112
rect 43346 6060 43352 6112
rect 43404 6100 43410 6112
rect 51902 6100 51908 6112
rect 43404 6072 51908 6100
rect 43404 6060 43410 6072
rect 51902 6060 51908 6072
rect 51960 6060 51966 6112
rect 53024 6100 53052 6199
rect 53190 6196 53196 6248
rect 53248 6236 53254 6248
rect 69474 6236 69480 6248
rect 53248 6208 69480 6236
rect 53248 6196 53254 6208
rect 69474 6196 69480 6208
rect 69532 6196 69538 6248
rect 81544 6245 81572 6276
rect 84194 6264 84200 6276
rect 84252 6264 84258 6316
rect 86586 6304 86592 6316
rect 86547 6276 86592 6304
rect 86586 6264 86592 6276
rect 86644 6264 86650 6316
rect 97810 6304 97816 6316
rect 93826 6276 97816 6304
rect 81529 6239 81587 6245
rect 81529 6236 81541 6239
rect 71608 6208 81541 6236
rect 53650 6128 53656 6180
rect 53708 6168 53714 6180
rect 71608 6168 71636 6208
rect 81529 6205 81541 6208
rect 81575 6205 81587 6239
rect 81894 6236 81900 6248
rect 81855 6208 81900 6236
rect 81529 6199 81587 6205
rect 81894 6196 81900 6208
rect 81952 6196 81958 6248
rect 84838 6236 84844 6248
rect 82004 6208 84844 6236
rect 53708 6140 71636 6168
rect 53708 6128 53714 6140
rect 81434 6128 81440 6180
rect 81492 6168 81498 6180
rect 81713 6171 81771 6177
rect 81713 6168 81725 6171
rect 81492 6140 81725 6168
rect 81492 6128 81498 6140
rect 81713 6137 81725 6140
rect 81759 6137 81771 6171
rect 81713 6131 81771 6137
rect 81805 6171 81863 6177
rect 81805 6137 81817 6171
rect 81851 6168 81863 6171
rect 82004 6168 82032 6208
rect 84838 6196 84844 6208
rect 84896 6196 84902 6248
rect 85942 6236 85948 6248
rect 85903 6208 85948 6236
rect 85942 6196 85948 6208
rect 86000 6196 86006 6248
rect 81851 6140 82032 6168
rect 81851 6137 81863 6140
rect 81805 6131 81863 6137
rect 61746 6100 61752 6112
rect 53024 6072 61752 6100
rect 61746 6060 61752 6072
rect 61804 6060 61810 6112
rect 69474 6060 69480 6112
rect 69532 6100 69538 6112
rect 93826 6100 93854 6276
rect 97810 6264 97816 6276
rect 97868 6264 97874 6316
rect 96982 6236 96988 6248
rect 96943 6208 96988 6236
rect 96982 6196 96988 6208
rect 97040 6196 97046 6248
rect 97626 6236 97632 6248
rect 97587 6208 97632 6236
rect 97626 6196 97632 6208
rect 97684 6196 97690 6248
rect 69532 6072 93854 6100
rect 69532 6060 69538 6072
rect 1104 6010 98808 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 50326 6010
rect 50378 5958 50390 6010
rect 50442 5958 50454 6010
rect 50506 5958 50518 6010
rect 50570 5958 81046 6010
rect 81098 5958 81110 6010
rect 81162 5958 81174 6010
rect 81226 5958 81238 6010
rect 81290 5958 98808 6010
rect 1104 5936 98808 5958
rect 8297 5899 8355 5905
rect 4448 5868 8064 5896
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 2409 5763 2467 5769
rect 2409 5760 2421 5763
rect 1912 5732 2421 5760
rect 1912 5720 1918 5732
rect 2409 5729 2421 5732
rect 2455 5729 2467 5763
rect 2409 5723 2467 5729
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 4448 5769 4476 5868
rect 7377 5831 7435 5837
rect 7377 5797 7389 5831
rect 7423 5828 7435 5831
rect 8036 5828 8064 5868
rect 8297 5865 8309 5899
rect 8343 5896 8355 5899
rect 20806 5896 20812 5908
rect 8343 5868 20812 5896
rect 8343 5865 8355 5868
rect 8297 5859 8355 5865
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 23382 5856 23388 5908
rect 23440 5896 23446 5908
rect 71590 5896 71596 5908
rect 23440 5868 71596 5896
rect 23440 5856 23446 5868
rect 71590 5856 71596 5868
rect 71648 5856 71654 5908
rect 73890 5896 73896 5908
rect 73851 5868 73896 5896
rect 73890 5856 73896 5868
rect 73948 5856 73954 5908
rect 91830 5856 91836 5908
rect 91888 5896 91894 5908
rect 95878 5896 95884 5908
rect 91888 5868 95556 5896
rect 95839 5868 95884 5896
rect 91888 5856 91894 5868
rect 11698 5828 11704 5840
rect 7423 5800 7879 5828
rect 8036 5800 11704 5828
rect 7423 5797 7435 5800
rect 7377 5791 7435 5797
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 2832 5732 3065 5760
rect 2832 5720 2838 5732
rect 3053 5729 3065 5732
rect 3099 5729 3111 5763
rect 3053 5723 3111 5729
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7009 5763 7067 5769
rect 7009 5760 7021 5763
rect 6972 5732 7021 5760
rect 6972 5720 6978 5732
rect 7009 5729 7021 5732
rect 7055 5729 7067 5763
rect 7650 5760 7656 5772
rect 7009 5723 7067 5729
rect 7116 5732 7656 5760
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 7116 5692 7144 5732
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7851 5769 7879 5800
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 11882 5788 11888 5840
rect 11940 5828 11946 5840
rect 17218 5828 17224 5840
rect 11940 5800 17224 5828
rect 11940 5788 11946 5800
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 17310 5788 17316 5840
rect 17368 5828 17374 5840
rect 22002 5828 22008 5840
rect 17368 5800 22008 5828
rect 17368 5788 17374 5800
rect 22002 5788 22008 5800
rect 22060 5788 22066 5840
rect 29730 5788 29736 5840
rect 29788 5828 29794 5840
rect 29788 5800 36584 5828
rect 29788 5788 29794 5800
rect 7836 5763 7894 5769
rect 7836 5729 7848 5763
rect 7882 5729 7894 5763
rect 7836 5723 7894 5729
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5760 8263 5763
rect 8573 5763 8631 5769
rect 8573 5760 8585 5763
rect 8251 5732 8585 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 8573 5729 8585 5732
rect 8619 5760 8631 5763
rect 15102 5760 15108 5772
rect 8619 5732 15108 5760
rect 8619 5729 8631 5732
rect 8573 5723 8631 5729
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 21634 5760 21640 5772
rect 15252 5732 21640 5760
rect 15252 5720 15258 5732
rect 21634 5720 21640 5732
rect 21692 5720 21698 5772
rect 26510 5760 26516 5772
rect 22480 5732 26372 5760
rect 26471 5732 26516 5760
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 5684 5664 7144 5692
rect 7668 5664 7941 5692
rect 5684 5652 5690 5664
rect 7668 5636 7696 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 7650 5584 7656 5636
rect 7708 5584 7714 5636
rect 8036 5624 8064 5655
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 22480 5692 22508 5732
rect 8812 5664 22508 5692
rect 8812 5652 8818 5664
rect 22830 5652 22836 5704
rect 22888 5692 22894 5704
rect 26234 5692 26240 5704
rect 22888 5664 24900 5692
rect 26195 5664 26240 5692
rect 22888 5652 22894 5664
rect 8202 5624 8208 5636
rect 8036 5596 8208 5624
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 11698 5584 11704 5636
rect 11756 5624 11762 5636
rect 23934 5624 23940 5636
rect 11756 5596 23940 5624
rect 11756 5584 11762 5596
rect 23934 5584 23940 5596
rect 23992 5584 23998 5636
rect 5074 5556 5080 5568
rect 5035 5528 5080 5556
rect 5074 5516 5080 5528
rect 5132 5516 5138 5568
rect 7377 5559 7435 5565
rect 7377 5525 7389 5559
rect 7423 5556 7435 5559
rect 7561 5559 7619 5565
rect 7561 5556 7573 5559
rect 7423 5528 7573 5556
rect 7423 5525 7435 5528
rect 7377 5519 7435 5525
rect 7561 5525 7573 5528
rect 7607 5556 7619 5559
rect 8386 5556 8392 5568
rect 7607 5528 8392 5556
rect 7607 5525 7619 5528
rect 7561 5519 7619 5525
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 15470 5556 15476 5568
rect 8536 5528 15476 5556
rect 8536 5516 8542 5528
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 17218 5516 17224 5568
rect 17276 5556 17282 5568
rect 24762 5556 24768 5568
rect 17276 5528 24768 5556
rect 17276 5516 17282 5528
rect 24762 5516 24768 5528
rect 24820 5516 24826 5568
rect 24872 5556 24900 5664
rect 26234 5652 26240 5664
rect 26292 5652 26298 5704
rect 26344 5692 26372 5732
rect 26510 5720 26516 5732
rect 26568 5720 26574 5772
rect 32398 5720 32404 5772
rect 32456 5760 32462 5772
rect 35986 5760 35992 5772
rect 32456 5732 35992 5760
rect 32456 5720 32462 5732
rect 35986 5720 35992 5732
rect 36044 5720 36050 5772
rect 36556 5760 36584 5800
rect 36630 5788 36636 5840
rect 36688 5828 36694 5840
rect 53466 5828 53472 5840
rect 36688 5800 53472 5828
rect 36688 5788 36694 5800
rect 53466 5788 53472 5800
rect 53524 5788 53530 5840
rect 58526 5788 58532 5840
rect 58584 5828 58590 5840
rect 58584 5800 80054 5828
rect 58584 5788 58590 5800
rect 36556 5732 41414 5760
rect 34790 5692 34796 5704
rect 26344 5664 34796 5692
rect 34790 5652 34796 5664
rect 34848 5652 34854 5704
rect 37642 5584 37648 5636
rect 37700 5624 37706 5636
rect 40678 5624 40684 5636
rect 37700 5596 40684 5624
rect 37700 5584 37706 5596
rect 40678 5584 40684 5596
rect 40736 5584 40742 5636
rect 41386 5624 41414 5732
rect 44910 5720 44916 5772
rect 44968 5760 44974 5772
rect 58986 5760 58992 5772
rect 44968 5732 58992 5760
rect 44968 5720 44974 5732
rect 58986 5720 58992 5732
rect 59044 5720 59050 5772
rect 74074 5760 74080 5772
rect 74035 5732 74080 5760
rect 74074 5720 74080 5732
rect 74132 5720 74138 5772
rect 80026 5760 80054 5800
rect 95237 5763 95295 5769
rect 95237 5760 95249 5763
rect 80026 5732 95249 5760
rect 95237 5729 95249 5732
rect 95283 5729 95295 5763
rect 95237 5723 95295 5729
rect 95326 5720 95332 5772
rect 95384 5760 95390 5772
rect 95528 5769 95556 5868
rect 95878 5856 95884 5868
rect 95936 5856 95942 5908
rect 95420 5763 95478 5769
rect 95420 5760 95432 5763
rect 95384 5732 95432 5760
rect 95384 5720 95390 5732
rect 95420 5729 95432 5732
rect 95466 5729 95478 5763
rect 95420 5723 95478 5729
rect 95513 5763 95571 5769
rect 95513 5729 95525 5763
rect 95559 5729 95571 5763
rect 95513 5723 95571 5729
rect 95789 5763 95847 5769
rect 95789 5729 95801 5763
rect 95835 5729 95847 5763
rect 95789 5723 95847 5729
rect 46750 5652 46756 5704
rect 46808 5692 46814 5704
rect 59446 5692 59452 5704
rect 46808 5664 59452 5692
rect 46808 5652 46814 5664
rect 59446 5652 59452 5664
rect 59504 5652 59510 5704
rect 83734 5692 83740 5704
rect 60706 5664 83740 5692
rect 60706 5624 60734 5664
rect 83734 5652 83740 5664
rect 83792 5652 83798 5704
rect 91462 5652 91468 5704
rect 91520 5692 91526 5704
rect 95605 5695 95663 5701
rect 95605 5692 95617 5695
rect 91520 5664 95617 5692
rect 91520 5652 91526 5664
rect 95605 5661 95617 5664
rect 95651 5661 95663 5695
rect 95605 5655 95663 5661
rect 67634 5624 67640 5636
rect 41386 5596 60734 5624
rect 61396 5596 67640 5624
rect 27617 5559 27675 5565
rect 27617 5556 27629 5559
rect 24872 5528 27629 5556
rect 27617 5525 27629 5528
rect 27663 5525 27675 5559
rect 27617 5519 27675 5525
rect 31110 5516 31116 5568
rect 31168 5556 31174 5568
rect 34054 5556 34060 5568
rect 31168 5528 34060 5556
rect 31168 5516 31174 5528
rect 34054 5516 34060 5528
rect 34112 5516 34118 5568
rect 36538 5516 36544 5568
rect 36596 5556 36602 5568
rect 46198 5556 46204 5568
rect 36596 5528 46204 5556
rect 36596 5516 36602 5528
rect 46198 5516 46204 5528
rect 46256 5516 46262 5568
rect 52822 5516 52828 5568
rect 52880 5556 52886 5568
rect 61396 5556 61424 5596
rect 67634 5584 67640 5596
rect 67692 5584 67698 5636
rect 69934 5584 69940 5636
rect 69992 5624 69998 5636
rect 69992 5596 80054 5624
rect 69992 5584 69998 5596
rect 52880 5528 61424 5556
rect 52880 5516 52886 5528
rect 61470 5516 61476 5568
rect 61528 5556 61534 5568
rect 62758 5556 62764 5568
rect 61528 5528 62764 5556
rect 61528 5516 61534 5528
rect 62758 5516 62764 5528
rect 62816 5516 62822 5568
rect 73982 5516 73988 5568
rect 74040 5556 74046 5568
rect 76558 5556 76564 5568
rect 74040 5528 76564 5556
rect 74040 5516 74046 5528
rect 76558 5516 76564 5528
rect 76616 5516 76622 5568
rect 80026 5556 80054 5596
rect 89346 5584 89352 5636
rect 89404 5624 89410 5636
rect 95804 5624 95832 5723
rect 96246 5720 96252 5772
rect 96304 5760 96310 5772
rect 96433 5763 96491 5769
rect 96433 5760 96445 5763
rect 96304 5732 96445 5760
rect 96304 5720 96310 5732
rect 96433 5729 96445 5732
rect 96479 5729 96491 5763
rect 96433 5723 96491 5729
rect 97537 5763 97595 5769
rect 97537 5729 97549 5763
rect 97583 5760 97595 5763
rect 99006 5760 99012 5772
rect 97583 5732 99012 5760
rect 97583 5729 97595 5732
rect 97537 5723 97595 5729
rect 99006 5720 99012 5732
rect 99064 5720 99070 5772
rect 89404 5596 95832 5624
rect 89404 5584 89410 5596
rect 95053 5559 95111 5565
rect 95053 5556 95065 5559
rect 80026 5528 95065 5556
rect 95053 5525 95065 5528
rect 95099 5556 95111 5559
rect 95326 5556 95332 5568
rect 95099 5528 95332 5556
rect 95099 5525 95111 5528
rect 95053 5519 95111 5525
rect 95326 5516 95332 5528
rect 95384 5516 95390 5568
rect 1104 5466 98808 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 65686 5466
rect 65738 5414 65750 5466
rect 65802 5414 65814 5466
rect 65866 5414 65878 5466
rect 65930 5414 96406 5466
rect 96458 5414 96470 5466
rect 96522 5414 96534 5466
rect 96586 5414 96598 5466
rect 96650 5414 98808 5466
rect 1104 5392 98808 5414
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 7558 5352 7564 5364
rect 6503 5324 7564 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 16022 5312 16028 5364
rect 16080 5352 16086 5364
rect 24302 5352 24308 5364
rect 16080 5324 24164 5352
rect 24263 5324 24308 5352
rect 16080 5312 16086 5324
rect 6273 5287 6331 5293
rect 6273 5253 6285 5287
rect 6319 5284 6331 5287
rect 22922 5284 22928 5296
rect 6319 5256 8524 5284
rect 6319 5253 6331 5256
rect 6273 5247 6331 5253
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5216 2467 5219
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 2455 5188 2697 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 2685 5185 2697 5188
rect 2731 5216 2743 5219
rect 2869 5219 2927 5225
rect 2869 5216 2881 5219
rect 2731 5188 2881 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 2869 5185 2881 5188
rect 2915 5216 2927 5219
rect 2915 5188 8432 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5148 3387 5151
rect 5258 5148 5264 5160
rect 3375 5120 5264 5148
rect 3375 5117 3387 5120
rect 3329 5111 3387 5117
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 6457 5151 6515 5157
rect 6457 5148 6469 5151
rect 5675 5120 6469 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 6457 5117 6469 5120
rect 6503 5117 6515 5151
rect 6457 5111 6515 5117
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6788 5120 6837 5148
rect 6788 5108 6794 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 8294 5148 8300 5160
rect 8067 5120 8300 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 1857 5083 1915 5089
rect 1857 5049 1869 5083
rect 1903 5080 1915 5083
rect 2038 5080 2044 5092
rect 1903 5052 2044 5080
rect 1903 5049 1915 5052
rect 1857 5043 1915 5049
rect 2038 5040 2044 5052
rect 2096 5040 2102 5092
rect 4341 5083 4399 5089
rect 4341 5049 4353 5083
rect 4387 5080 4399 5083
rect 6273 5083 6331 5089
rect 6273 5080 6285 5083
rect 4387 5052 6285 5080
rect 4387 5049 4399 5052
rect 4341 5043 4399 5049
rect 6273 5049 6285 5052
rect 6319 5049 6331 5083
rect 6273 5043 6331 5049
rect 7009 5083 7067 5089
rect 7009 5049 7021 5083
rect 7055 5080 7067 5083
rect 7055 5052 7089 5080
rect 7055 5049 7067 5052
rect 7009 5043 7067 5049
rect 474 4972 480 5024
rect 532 5012 538 5024
rect 1949 5015 2007 5021
rect 1949 5012 1961 5015
rect 532 4984 1961 5012
rect 532 4972 538 4984
rect 1949 4981 1961 4984
rect 1995 4981 2007 5015
rect 3418 5012 3424 5024
rect 3379 4984 3424 5012
rect 1949 4975 2007 4981
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 4433 5015 4491 5021
rect 4433 4981 4445 5015
rect 4479 5012 4491 5015
rect 4890 5012 4896 5024
rect 4479 4984 4896 5012
rect 4479 4981 4491 4984
rect 4433 4975 4491 4981
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5684 4984 5733 5012
rect 5684 4972 5690 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 5721 4975 5779 4981
rect 6733 5015 6791 5021
rect 6733 4981 6745 5015
rect 6779 5012 6791 5015
rect 7024 5012 7052 5043
rect 8202 5012 8208 5024
rect 6779 4984 8208 5012
rect 6779 4981 6791 4984
rect 6733 4975 6791 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 8404 5012 8432 5188
rect 8496 5080 8524 5256
rect 8588 5256 22928 5284
rect 8588 5225 8616 5256
rect 22922 5244 22928 5256
rect 22980 5244 22986 5296
rect 24136 5284 24164 5324
rect 24302 5312 24308 5324
rect 24360 5312 24366 5364
rect 24964 5324 55904 5352
rect 24964 5284 24992 5324
rect 24136 5256 24992 5284
rect 29270 5244 29276 5296
rect 29328 5284 29334 5296
rect 34333 5287 34391 5293
rect 29328 5256 34100 5284
rect 29328 5244 29334 5256
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 12529 5219 12587 5225
rect 12529 5185 12541 5219
rect 12575 5216 12587 5219
rect 23198 5216 23204 5228
rect 12575 5188 23060 5216
rect 23159 5188 23204 5216
rect 12575 5185 12587 5188
rect 12529 5179 12587 5185
rect 9122 5148 9128 5160
rect 9083 5120 9128 5148
rect 9122 5108 9128 5120
rect 9180 5108 9186 5160
rect 21726 5108 21732 5160
rect 21784 5148 21790 5160
rect 22925 5151 22983 5157
rect 22925 5148 22937 5151
rect 21784 5120 22937 5148
rect 21784 5108 21790 5120
rect 22925 5117 22937 5120
rect 22971 5117 22983 5151
rect 23032 5148 23060 5188
rect 23198 5176 23204 5188
rect 23256 5176 23262 5228
rect 31386 5216 31392 5228
rect 23308 5188 31392 5216
rect 23308 5148 23336 5188
rect 31386 5176 31392 5188
rect 31444 5176 31450 5228
rect 25038 5148 25044 5160
rect 23032 5120 23336 5148
rect 24999 5120 25044 5148
rect 22925 5111 22983 5117
rect 25038 5108 25044 5120
rect 25096 5108 25102 5160
rect 25682 5148 25688 5160
rect 25643 5120 25688 5148
rect 25682 5108 25688 5120
rect 25740 5108 25746 5160
rect 26326 5148 26332 5160
rect 26287 5120 26332 5148
rect 26326 5108 26332 5120
rect 26384 5108 26390 5160
rect 27798 5148 27804 5160
rect 27759 5120 27804 5148
rect 27798 5108 27804 5120
rect 27856 5108 27862 5160
rect 33502 5108 33508 5160
rect 33560 5148 33566 5160
rect 33781 5151 33839 5157
rect 33781 5148 33793 5151
rect 33560 5120 33793 5148
rect 33560 5108 33566 5120
rect 33781 5117 33793 5120
rect 33827 5117 33839 5151
rect 33781 5111 33839 5117
rect 18598 5080 18604 5092
rect 8496 5052 18604 5080
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 31662 5040 31668 5092
rect 31720 5080 31726 5092
rect 34072 5089 34100 5256
rect 34333 5253 34345 5287
rect 34379 5253 34391 5287
rect 34333 5247 34391 5253
rect 34348 5216 34376 5247
rect 34606 5244 34612 5296
rect 34664 5284 34670 5296
rect 38010 5284 38016 5296
rect 34664 5256 38016 5284
rect 34664 5244 34670 5256
rect 38010 5244 38016 5256
rect 38068 5244 38074 5296
rect 38473 5287 38531 5293
rect 38473 5253 38485 5287
rect 38519 5284 38531 5287
rect 38519 5256 46244 5284
rect 38519 5253 38531 5256
rect 38473 5247 38531 5253
rect 43438 5216 43444 5228
rect 34348 5188 43444 5216
rect 43438 5176 43444 5188
rect 43496 5176 43502 5228
rect 45002 5216 45008 5228
rect 44928 5188 45008 5216
rect 34146 5108 34152 5160
rect 34204 5148 34210 5160
rect 36357 5151 36415 5157
rect 34204 5120 34249 5148
rect 34204 5108 34210 5120
rect 36357 5117 36369 5151
rect 36403 5148 36415 5151
rect 36630 5148 36636 5160
rect 36403 5120 36636 5148
rect 36403 5117 36415 5120
rect 36357 5111 36415 5117
rect 36630 5108 36636 5120
rect 36688 5108 36694 5160
rect 36814 5148 36820 5160
rect 36775 5120 36820 5148
rect 36814 5108 36820 5120
rect 36872 5108 36878 5160
rect 36909 5151 36967 5157
rect 36909 5117 36921 5151
rect 36955 5148 36967 5151
rect 37182 5148 37188 5160
rect 36955 5120 37188 5148
rect 36955 5117 36967 5120
rect 36909 5111 36967 5117
rect 37182 5108 37188 5120
rect 37240 5108 37246 5160
rect 38746 5148 38752 5160
rect 38707 5120 38752 5148
rect 38746 5108 38752 5120
rect 38804 5108 38810 5160
rect 39206 5148 39212 5160
rect 39167 5120 39212 5148
rect 39206 5108 39212 5120
rect 39264 5108 39270 5160
rect 44928 5157 44956 5188
rect 45002 5176 45008 5188
rect 45060 5176 45066 5228
rect 45278 5216 45284 5228
rect 45239 5188 45284 5216
rect 45278 5176 45284 5188
rect 45336 5176 45342 5228
rect 46216 5216 46244 5256
rect 46290 5244 46296 5296
rect 46348 5284 46354 5296
rect 55766 5284 55772 5296
rect 46348 5256 55772 5284
rect 46348 5244 46354 5256
rect 55766 5244 55772 5256
rect 55824 5244 55830 5296
rect 55876 5284 55904 5324
rect 55950 5312 55956 5364
rect 56008 5352 56014 5364
rect 65245 5355 65303 5361
rect 65245 5352 65257 5355
rect 56008 5324 65257 5352
rect 56008 5312 56014 5324
rect 65245 5321 65257 5324
rect 65291 5321 65303 5355
rect 65245 5315 65303 5321
rect 66162 5312 66168 5364
rect 66220 5352 66226 5364
rect 73982 5352 73988 5364
rect 66220 5324 73988 5352
rect 66220 5312 66226 5324
rect 73982 5312 73988 5324
rect 74040 5312 74046 5364
rect 74074 5312 74080 5364
rect 74132 5352 74138 5364
rect 79689 5355 79747 5361
rect 79689 5352 79701 5355
rect 74132 5324 79701 5352
rect 74132 5312 74138 5324
rect 79689 5321 79701 5324
rect 79735 5321 79747 5355
rect 79689 5315 79747 5321
rect 82170 5312 82176 5364
rect 82228 5352 82234 5364
rect 90818 5352 90824 5364
rect 82228 5324 90824 5352
rect 82228 5312 82234 5324
rect 90818 5312 90824 5324
rect 90876 5312 90882 5364
rect 55876 5256 56180 5284
rect 51994 5216 52000 5228
rect 46216 5188 52000 5216
rect 51994 5176 52000 5188
rect 52052 5176 52058 5228
rect 52178 5176 52184 5228
rect 52236 5216 52242 5228
rect 55858 5216 55864 5228
rect 52236 5188 55864 5216
rect 52236 5176 52242 5188
rect 55858 5176 55864 5188
rect 55916 5176 55922 5228
rect 44913 5151 44971 5157
rect 44913 5117 44925 5151
rect 44959 5117 44971 5151
rect 54570 5148 54576 5160
rect 44913 5111 44971 5117
rect 45112 5120 54576 5148
rect 33965 5083 34023 5089
rect 33965 5080 33977 5083
rect 31720 5052 33977 5080
rect 31720 5040 31726 5052
rect 33965 5049 33977 5052
rect 34011 5049 34023 5083
rect 33965 5043 34023 5049
rect 34057 5083 34115 5089
rect 34057 5049 34069 5083
rect 34103 5049 34115 5083
rect 34057 5043 34115 5049
rect 34256 5052 41414 5080
rect 34256 5012 34284 5052
rect 36446 5012 36452 5024
rect 8404 4984 34284 5012
rect 36407 4984 36452 5012
rect 36446 4972 36452 4984
rect 36504 4972 36510 5024
rect 36814 4972 36820 5024
rect 36872 5012 36878 5024
rect 38473 5015 38531 5021
rect 38473 5012 38485 5015
rect 36872 4984 38485 5012
rect 36872 4972 36878 4984
rect 38473 4981 38485 4984
rect 38519 4981 38531 5015
rect 41386 5012 41414 5052
rect 44082 5040 44088 5092
rect 44140 5080 44146 5092
rect 45112 5080 45140 5120
rect 54570 5108 54576 5120
rect 54628 5108 54634 5160
rect 56152 5148 56180 5256
rect 57882 5244 57888 5296
rect 57940 5284 57946 5296
rect 64966 5284 64972 5296
rect 57940 5256 64972 5284
rect 57940 5244 57946 5256
rect 64966 5244 64972 5256
rect 65024 5244 65030 5296
rect 65150 5244 65156 5296
rect 65208 5284 65214 5296
rect 65518 5284 65524 5296
rect 65208 5256 65524 5284
rect 65208 5244 65214 5256
rect 65518 5244 65524 5256
rect 65576 5244 65582 5296
rect 67082 5244 67088 5296
rect 67140 5284 67146 5296
rect 68094 5284 68100 5296
rect 67140 5256 68100 5284
rect 67140 5244 67146 5256
rect 68094 5244 68100 5256
rect 68152 5244 68158 5296
rect 68554 5244 68560 5296
rect 68612 5284 68618 5296
rect 68612 5256 84884 5284
rect 68612 5244 68618 5256
rect 56226 5176 56232 5228
rect 56284 5216 56290 5228
rect 59078 5216 59084 5228
rect 56284 5188 59084 5216
rect 56284 5176 56290 5188
rect 59078 5176 59084 5188
rect 59136 5176 59142 5228
rect 65334 5176 65340 5228
rect 65392 5216 65398 5228
rect 71038 5216 71044 5228
rect 65392 5188 71044 5216
rect 65392 5176 65398 5188
rect 71038 5176 71044 5188
rect 71096 5176 71102 5228
rect 82170 5216 82176 5228
rect 71148 5188 82176 5216
rect 58894 5148 58900 5160
rect 56152 5120 58900 5148
rect 58894 5108 58900 5120
rect 58952 5108 58958 5160
rect 64598 5108 64604 5160
rect 64656 5148 64662 5160
rect 64693 5151 64751 5157
rect 64693 5148 64705 5151
rect 64656 5120 64705 5148
rect 64656 5108 64662 5120
rect 64693 5117 64705 5120
rect 64739 5117 64751 5151
rect 64874 5148 64880 5160
rect 64835 5120 64880 5148
rect 64693 5111 64751 5117
rect 64874 5108 64880 5120
rect 64932 5108 64938 5160
rect 65058 5148 65064 5160
rect 65019 5120 65064 5148
rect 65058 5108 65064 5120
rect 65116 5108 65122 5160
rect 65150 5108 65156 5160
rect 65208 5148 65214 5160
rect 71148 5148 71176 5188
rect 82170 5176 82176 5188
rect 82228 5176 82234 5228
rect 82630 5176 82636 5228
rect 82688 5216 82694 5228
rect 82725 5219 82783 5225
rect 82725 5216 82737 5219
rect 82688 5188 82737 5216
rect 82688 5176 82694 5188
rect 82725 5185 82737 5188
rect 82771 5185 82783 5219
rect 84856 5216 84884 5256
rect 91373 5219 91431 5225
rect 91373 5216 91385 5219
rect 84856 5188 91385 5216
rect 82725 5179 82783 5185
rect 91373 5185 91385 5188
rect 91419 5185 91431 5219
rect 91373 5179 91431 5185
rect 76926 5148 76932 5160
rect 65208 5120 71176 5148
rect 76887 5120 76932 5148
rect 65208 5108 65214 5120
rect 76926 5108 76932 5120
rect 76984 5108 76990 5160
rect 77478 5108 77484 5160
rect 77536 5148 77542 5160
rect 77573 5151 77631 5157
rect 77573 5148 77585 5151
rect 77536 5120 77585 5148
rect 77536 5108 77542 5120
rect 77573 5117 77585 5120
rect 77619 5117 77631 5151
rect 77573 5111 77631 5117
rect 79689 5151 79747 5157
rect 79689 5117 79701 5151
rect 79735 5148 79747 5151
rect 82081 5151 82139 5157
rect 82081 5148 82093 5151
rect 79735 5120 82093 5148
rect 79735 5117 79747 5120
rect 79689 5111 79747 5117
rect 82081 5117 82093 5120
rect 82127 5148 82139 5151
rect 82449 5151 82507 5157
rect 82449 5148 82461 5151
rect 82127 5120 82461 5148
rect 82127 5117 82139 5120
rect 82081 5111 82139 5117
rect 82449 5117 82461 5120
rect 82495 5117 82507 5151
rect 82449 5111 82507 5117
rect 85853 5151 85911 5157
rect 85853 5117 85865 5151
rect 85899 5148 85911 5151
rect 87322 5148 87328 5160
rect 85899 5120 87328 5148
rect 85899 5117 85911 5120
rect 85853 5111 85911 5117
rect 87322 5108 87328 5120
rect 87380 5108 87386 5160
rect 87598 5148 87604 5160
rect 87559 5120 87604 5148
rect 87598 5108 87604 5120
rect 87656 5108 87662 5160
rect 88061 5151 88119 5157
rect 88061 5117 88073 5151
rect 88107 5117 88119 5151
rect 88061 5111 88119 5117
rect 59262 5080 59268 5092
rect 44140 5052 45140 5080
rect 51736 5052 59268 5080
rect 44140 5040 44146 5052
rect 51736 5012 51764 5052
rect 59262 5040 59268 5052
rect 59320 5040 59326 5092
rect 64782 5040 64788 5092
rect 64840 5080 64846 5092
rect 64969 5083 65027 5089
rect 64969 5080 64981 5083
rect 64840 5052 64981 5080
rect 64840 5040 64846 5052
rect 64969 5049 64981 5052
rect 65015 5049 65027 5083
rect 64969 5043 65027 5049
rect 65076 5052 80054 5080
rect 41386 4984 51764 5012
rect 38473 4975 38531 4981
rect 51994 4972 52000 5024
rect 52052 5012 52058 5024
rect 65076 5012 65104 5052
rect 52052 4984 65104 5012
rect 52052 4972 52058 4984
rect 65518 4972 65524 5024
rect 65576 5012 65582 5024
rect 68830 5012 68836 5024
rect 65576 4984 68836 5012
rect 65576 4972 65582 4984
rect 68830 4972 68836 4984
rect 68888 4972 68894 5024
rect 80026 5012 80054 5052
rect 82170 5040 82176 5092
rect 82228 5080 82234 5092
rect 82265 5083 82323 5089
rect 82265 5080 82277 5083
rect 82228 5052 82277 5080
rect 82228 5040 82234 5052
rect 82265 5049 82277 5052
rect 82311 5049 82323 5083
rect 85945 5083 86003 5089
rect 85945 5080 85957 5083
rect 82265 5043 82323 5049
rect 82372 5052 85957 5080
rect 82372 5012 82400 5052
rect 85945 5049 85957 5052
rect 85991 5049 86003 5083
rect 85945 5043 86003 5049
rect 80026 4984 82400 5012
rect 87230 4972 87236 5024
rect 87288 5012 87294 5024
rect 88076 5012 88104 5111
rect 88518 5108 88524 5160
rect 88576 5148 88582 5160
rect 88705 5151 88763 5157
rect 88705 5148 88717 5151
rect 88576 5120 88717 5148
rect 88576 5108 88582 5120
rect 88705 5117 88717 5120
rect 88751 5117 88763 5151
rect 90726 5148 90732 5160
rect 90687 5120 90732 5148
rect 88705 5111 88763 5117
rect 90726 5108 90732 5120
rect 90784 5108 90790 5160
rect 90818 5108 90824 5160
rect 90876 5148 90882 5160
rect 90913 5151 90971 5157
rect 90913 5148 90925 5151
rect 90876 5120 90925 5148
rect 90876 5108 90882 5120
rect 90913 5117 90925 5120
rect 90959 5117 90971 5151
rect 90913 5111 90971 5117
rect 91097 5151 91155 5157
rect 91097 5117 91109 5151
rect 91143 5117 91155 5151
rect 91462 5148 91468 5160
rect 91423 5120 91468 5148
rect 91097 5111 91155 5117
rect 91112 5080 91140 5111
rect 91462 5108 91468 5120
rect 91520 5108 91526 5160
rect 92934 5148 92940 5160
rect 92895 5120 92940 5148
rect 92934 5108 92940 5120
rect 92992 5108 92998 5160
rect 94225 5151 94283 5157
rect 94225 5117 94237 5151
rect 94271 5117 94283 5151
rect 94225 5111 94283 5117
rect 94869 5151 94927 5157
rect 94869 5117 94881 5151
rect 94915 5148 94927 5151
rect 95694 5148 95700 5160
rect 94915 5120 95700 5148
rect 94915 5117 94927 5120
rect 94869 5111 94927 5117
rect 91830 5080 91836 5092
rect 91112 5052 91836 5080
rect 91830 5040 91836 5052
rect 91888 5040 91894 5092
rect 87288 4984 88104 5012
rect 87288 4972 87294 4984
rect 89806 4972 89812 5024
rect 89864 5012 89870 5024
rect 90085 5015 90143 5021
rect 90085 5012 90097 5015
rect 89864 4984 90097 5012
rect 89864 4972 89870 4984
rect 90085 4981 90097 4984
rect 90131 5012 90143 5015
rect 90361 5015 90419 5021
rect 90361 5012 90373 5015
rect 90131 4984 90373 5012
rect 90131 4981 90143 4984
rect 90085 4975 90143 4981
rect 90361 4981 90373 4984
rect 90407 5012 90419 5015
rect 90545 5015 90603 5021
rect 90545 5012 90557 5015
rect 90407 4984 90557 5012
rect 90407 4981 90419 4984
rect 90361 4975 90419 4981
rect 90545 4981 90557 4984
rect 90591 5012 90603 5015
rect 91925 5015 91983 5021
rect 91925 5012 91937 5015
rect 90591 4984 91937 5012
rect 90591 4981 90603 4984
rect 90545 4975 90603 4981
rect 91925 4981 91937 4984
rect 91971 5012 91983 5015
rect 92201 5015 92259 5021
rect 92201 5012 92213 5015
rect 91971 4984 92213 5012
rect 91971 4981 91983 4984
rect 91925 4975 91983 4981
rect 92201 4981 92213 4984
rect 92247 5012 92259 5015
rect 92385 5015 92443 5021
rect 92385 5012 92397 5015
rect 92247 4984 92397 5012
rect 92247 4981 92259 4984
rect 92201 4975 92259 4981
rect 92385 4981 92397 4984
rect 92431 5012 92443 5015
rect 92569 5015 92627 5021
rect 92569 5012 92581 5015
rect 92431 4984 92581 5012
rect 92431 4981 92443 4984
rect 92385 4975 92443 4981
rect 92569 4981 92581 4984
rect 92615 5012 92627 5015
rect 92753 5015 92811 5021
rect 92753 5012 92765 5015
rect 92615 4984 92765 5012
rect 92615 4981 92627 4984
rect 92569 4975 92627 4981
rect 92753 4981 92765 4984
rect 92799 4981 92811 5015
rect 94240 5012 94268 5111
rect 95694 5108 95700 5120
rect 95752 5108 95758 5160
rect 95973 5151 96031 5157
rect 95973 5117 95985 5151
rect 96019 5117 96031 5151
rect 95973 5111 96031 5117
rect 97169 5151 97227 5157
rect 97169 5117 97181 5151
rect 97215 5117 97227 5151
rect 97810 5148 97816 5160
rect 97771 5120 97816 5148
rect 97169 5111 97227 5117
rect 95234 5040 95240 5092
rect 95292 5080 95298 5092
rect 95988 5080 96016 5111
rect 95292 5052 96016 5080
rect 97184 5080 97212 5111
rect 97810 5108 97816 5120
rect 97868 5108 97874 5160
rect 98454 5080 98460 5092
rect 97184 5052 98460 5080
rect 95292 5040 95298 5052
rect 98454 5040 98460 5052
rect 98512 5040 98518 5092
rect 96154 5012 96160 5024
rect 94240 4984 96160 5012
rect 92753 4975 92811 4981
rect 96154 4972 96160 4984
rect 96212 4972 96218 5024
rect 1104 4922 98808 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 50326 4922
rect 50378 4870 50390 4922
rect 50442 4870 50454 4922
rect 50506 4870 50518 4922
rect 50570 4870 81046 4922
rect 81098 4870 81110 4922
rect 81162 4870 81174 4922
rect 81226 4870 81238 4922
rect 81290 4870 98808 4922
rect 1104 4848 98808 4870
rect 1946 4808 1952 4820
rect 1907 4780 1952 4808
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2498 4808 2504 4820
rect 2459 4780 2504 4808
rect 2498 4768 2504 4780
rect 2556 4808 2562 4820
rect 6825 4811 6883 4817
rect 2556 4780 2912 4808
rect 2556 4768 2562 4780
rect 2884 4749 2912 4780
rect 6825 4777 6837 4811
rect 6871 4808 6883 4811
rect 7009 4811 7067 4817
rect 7009 4808 7021 4811
rect 6871 4780 7021 4808
rect 6871 4777 6883 4780
rect 6825 4771 6883 4777
rect 7009 4777 7021 4780
rect 7055 4808 7067 4811
rect 7561 4811 7619 4817
rect 7561 4808 7573 4811
rect 7055 4780 7573 4808
rect 7055 4777 7067 4780
rect 7009 4771 7067 4777
rect 7561 4777 7573 4780
rect 7607 4808 7619 4811
rect 8938 4808 8944 4820
rect 7607 4780 8944 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4709 2927 4743
rect 6638 4740 6644 4752
rect 6599 4712 6644 4740
rect 2869 4703 2927 4709
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 842 4632 848 4684
rect 900 4672 906 4684
rect 1857 4675 1915 4681
rect 1857 4672 1869 4675
rect 900 4644 1869 4672
rect 900 4632 906 4644
rect 1857 4641 1869 4644
rect 1903 4641 1915 4675
rect 1857 4635 1915 4641
rect 3973 4675 4031 4681
rect 3973 4641 3985 4675
rect 4019 4672 4031 4675
rect 4157 4675 4215 4681
rect 4157 4672 4169 4675
rect 4019 4644 4169 4672
rect 4019 4641 4031 4644
rect 3973 4635 4031 4641
rect 4157 4641 4169 4644
rect 4203 4672 4215 4675
rect 4341 4675 4399 4681
rect 4341 4672 4353 4675
rect 4203 4644 4353 4672
rect 4203 4641 4215 4644
rect 4157 4635 4215 4641
rect 4341 4641 4353 4644
rect 4387 4672 4399 4675
rect 4525 4675 4583 4681
rect 4525 4672 4537 4675
rect 4387 4644 4537 4672
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 4525 4641 4537 4644
rect 4571 4672 4583 4675
rect 4709 4675 4767 4681
rect 4709 4672 4721 4675
rect 4571 4644 4721 4672
rect 4571 4641 4583 4644
rect 4525 4635 4583 4641
rect 4709 4641 4721 4644
rect 4755 4672 4767 4675
rect 4893 4675 4951 4681
rect 4893 4672 4905 4675
rect 4755 4644 4905 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 4893 4641 4905 4644
rect 4939 4672 4951 4675
rect 5261 4675 5319 4681
rect 5261 4672 5273 4675
rect 4939 4644 5273 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 5261 4641 5273 4644
rect 5307 4672 5319 4675
rect 6840 4672 6868 4771
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 25130 4768 25136 4820
rect 25188 4808 25194 4820
rect 32861 4811 32919 4817
rect 25188 4780 31754 4808
rect 25188 4768 25194 4780
rect 7282 4740 7288 4752
rect 7243 4712 7288 4740
rect 7282 4700 7288 4712
rect 7340 4740 7346 4752
rect 7653 4743 7711 4749
rect 7653 4740 7665 4743
rect 7340 4712 7665 4740
rect 7340 4700 7346 4712
rect 7653 4709 7665 4712
rect 7699 4709 7711 4743
rect 7653 4703 7711 4709
rect 7929 4743 7987 4749
rect 7929 4709 7941 4743
rect 7975 4740 7987 4743
rect 8110 4740 8116 4752
rect 7975 4712 8116 4740
rect 7975 4709 7987 4712
rect 7929 4703 7987 4709
rect 8110 4700 8116 4712
rect 8168 4700 8174 4752
rect 20070 4700 20076 4752
rect 20128 4740 20134 4752
rect 24946 4740 24952 4752
rect 20128 4712 24952 4740
rect 20128 4700 20134 4712
rect 24946 4700 24952 4712
rect 25004 4700 25010 4752
rect 25314 4700 25320 4752
rect 25372 4740 25378 4752
rect 25958 4740 25964 4752
rect 25372 4712 25964 4740
rect 25372 4700 25378 4712
rect 25958 4700 25964 4712
rect 26016 4740 26022 4752
rect 26973 4743 27031 4749
rect 26016 4712 26372 4740
rect 26016 4700 26022 4712
rect 5307 4644 6868 4672
rect 5307 4641 5319 4644
rect 5261 4635 5319 4641
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 9493 4675 9551 4681
rect 9493 4672 9505 4675
rect 8904 4644 9505 4672
rect 8904 4632 8910 4644
rect 9493 4641 9505 4644
rect 9539 4641 9551 4675
rect 10594 4672 10600 4684
rect 10555 4644 10600 4672
rect 9493 4635 9551 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 11238 4672 11244 4684
rect 11199 4644 11244 4672
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 11882 4672 11888 4684
rect 11843 4644 11888 4672
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 12492 4644 12541 4672
rect 12492 4632 12498 4644
rect 12529 4641 12541 4644
rect 12575 4641 12587 4675
rect 12529 4635 12587 4641
rect 14274 4632 14280 4684
rect 14332 4672 14338 4684
rect 14737 4675 14795 4681
rect 14737 4672 14749 4675
rect 14332 4644 14749 4672
rect 14332 4632 14338 4644
rect 14737 4641 14749 4644
rect 14783 4641 14795 4675
rect 14737 4635 14795 4641
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15381 4675 15439 4681
rect 15381 4672 15393 4675
rect 15252 4644 15393 4672
rect 15252 4632 15258 4644
rect 15381 4641 15393 4644
rect 15427 4641 15439 4675
rect 16114 4672 16120 4684
rect 16075 4644 16120 4672
rect 15381 4635 15439 4641
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 17310 4672 17316 4684
rect 17271 4644 17316 4672
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 17954 4672 17960 4684
rect 17915 4644 17960 4672
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 18598 4672 18604 4684
rect 18559 4644 18604 4672
rect 18598 4632 18604 4644
rect 18656 4632 18662 4684
rect 19886 4632 19892 4684
rect 19944 4672 19950 4684
rect 19981 4675 20039 4681
rect 19981 4672 19993 4675
rect 19944 4644 19993 4672
rect 19944 4632 19950 4644
rect 19981 4641 19993 4644
rect 20027 4641 20039 4675
rect 20990 4672 20996 4684
rect 20951 4644 20996 4672
rect 19981 4635 20039 4641
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 21726 4632 21732 4684
rect 21784 4672 21790 4684
rect 22005 4675 22063 4681
rect 22005 4672 22017 4675
rect 21784 4644 22017 4672
rect 21784 4632 21790 4644
rect 22005 4641 22017 4644
rect 22051 4641 22063 4675
rect 22646 4672 22652 4684
rect 22607 4644 22652 4672
rect 22005 4635 22063 4641
rect 22646 4632 22652 4644
rect 22704 4632 22710 4684
rect 23198 4632 23204 4684
rect 23256 4672 23262 4684
rect 23293 4675 23351 4681
rect 23293 4672 23305 4675
rect 23256 4644 23305 4672
rect 23256 4632 23262 4644
rect 23293 4641 23305 4644
rect 23339 4641 23351 4675
rect 23293 4635 23351 4641
rect 25685 4675 25743 4681
rect 25685 4641 25697 4675
rect 25731 4672 25743 4675
rect 25866 4672 25872 4684
rect 25731 4644 25872 4672
rect 25731 4641 25743 4644
rect 25685 4635 25743 4641
rect 25866 4632 25872 4644
rect 25924 4632 25930 4684
rect 26050 4672 26056 4684
rect 26011 4644 26056 4672
rect 26050 4632 26056 4644
rect 26108 4632 26114 4684
rect 26344 4681 26372 4712
rect 26973 4709 26985 4743
rect 27019 4740 27031 4743
rect 27430 4740 27436 4752
rect 27019 4712 27436 4740
rect 27019 4709 27031 4712
rect 26973 4703 27031 4709
rect 27430 4700 27436 4712
rect 27488 4700 27494 4752
rect 31726 4740 31754 4780
rect 32861 4777 32873 4811
rect 32907 4808 32919 4811
rect 32950 4808 32956 4820
rect 32907 4780 32956 4808
rect 32907 4777 32919 4780
rect 32861 4771 32919 4777
rect 32950 4768 32956 4780
rect 33008 4768 33014 4820
rect 33318 4768 33324 4820
rect 33376 4808 33382 4820
rect 37366 4808 37372 4820
rect 33376 4780 37372 4808
rect 33376 4768 33382 4780
rect 37366 4768 37372 4780
rect 37424 4768 37430 4820
rect 52914 4768 52920 4820
rect 52972 4808 52978 4820
rect 53285 4811 53343 4817
rect 53285 4808 53297 4811
rect 52972 4780 53297 4808
rect 52972 4768 52978 4780
rect 53285 4777 53297 4780
rect 53331 4808 53343 4811
rect 53929 4811 53987 4817
rect 53929 4808 53941 4811
rect 53331 4780 53941 4808
rect 53331 4777 53343 4780
rect 53285 4771 53343 4777
rect 53929 4777 53941 4780
rect 53975 4808 53987 4811
rect 54113 4811 54171 4817
rect 54113 4808 54125 4811
rect 53975 4780 54125 4808
rect 53975 4777 53987 4780
rect 53929 4771 53987 4777
rect 54113 4777 54125 4780
rect 54159 4777 54171 4811
rect 54113 4771 54171 4777
rect 54205 4811 54263 4817
rect 54205 4777 54217 4811
rect 54251 4808 54263 4811
rect 54251 4780 78352 4808
rect 54251 4777 54263 4780
rect 54205 4771 54263 4777
rect 36538 4740 36544 4752
rect 31726 4712 36544 4740
rect 36538 4700 36544 4712
rect 36596 4700 36602 4752
rect 39025 4743 39083 4749
rect 39025 4709 39037 4743
rect 39071 4740 39083 4743
rect 39942 4740 39948 4752
rect 39071 4712 39948 4740
rect 39071 4709 39083 4712
rect 39025 4703 39083 4709
rect 39942 4700 39948 4712
rect 40000 4700 40006 4752
rect 50982 4700 50988 4752
rect 51040 4740 51046 4752
rect 51040 4712 54432 4740
rect 51040 4700 51046 4712
rect 26329 4675 26387 4681
rect 26329 4641 26341 4675
rect 26375 4641 26387 4675
rect 26329 4635 26387 4641
rect 26421 4675 26479 4681
rect 26421 4641 26433 4675
rect 26467 4672 26479 4675
rect 26878 4672 26884 4684
rect 26467 4644 26884 4672
rect 26467 4641 26479 4644
rect 26421 4635 26479 4641
rect 26878 4632 26884 4644
rect 26936 4632 26942 4684
rect 27062 4632 27068 4684
rect 27120 4672 27126 4684
rect 27525 4675 27583 4681
rect 27525 4672 27537 4675
rect 27120 4644 27537 4672
rect 27120 4632 27126 4644
rect 27525 4641 27537 4644
rect 27571 4641 27583 4675
rect 29086 4672 29092 4684
rect 29047 4644 29092 4672
rect 27525 4635 27583 4641
rect 29086 4632 29092 4644
rect 29144 4632 29150 4684
rect 32950 4632 32956 4684
rect 33008 4672 33014 4684
rect 33137 4675 33195 4681
rect 33137 4672 33149 4675
rect 33008 4644 33149 4672
rect 33008 4632 33014 4644
rect 33137 4641 33149 4644
rect 33183 4641 33195 4675
rect 34238 4672 34244 4684
rect 34199 4644 34244 4672
rect 33137 4635 33195 4641
rect 34238 4632 34244 4644
rect 34296 4632 34302 4684
rect 36078 4672 36084 4684
rect 36039 4644 36084 4672
rect 36078 4632 36084 4644
rect 36136 4632 36142 4684
rect 36630 4632 36636 4684
rect 36688 4672 36694 4684
rect 36725 4675 36783 4681
rect 36725 4672 36737 4675
rect 36688 4644 36737 4672
rect 36688 4632 36694 4644
rect 36725 4641 36737 4644
rect 36771 4641 36783 4675
rect 36725 4635 36783 4641
rect 37277 4675 37335 4681
rect 37277 4641 37289 4675
rect 37323 4672 37335 4675
rect 37642 4672 37648 4684
rect 37323 4644 37648 4672
rect 37323 4641 37335 4644
rect 37277 4635 37335 4641
rect 37642 4632 37648 4644
rect 37700 4632 37706 4684
rect 39482 4672 39488 4684
rect 39443 4644 39488 4672
rect 39482 4632 39488 4644
rect 39540 4632 39546 4684
rect 40310 4632 40316 4684
rect 40368 4672 40374 4684
rect 40957 4675 41015 4681
rect 40957 4672 40969 4675
rect 40368 4644 40969 4672
rect 40368 4632 40374 4644
rect 40957 4641 40969 4644
rect 41003 4641 41015 4675
rect 40957 4635 41015 4641
rect 41506 4632 41512 4684
rect 41564 4672 41570 4684
rect 41601 4675 41659 4681
rect 41601 4672 41613 4675
rect 41564 4644 41613 4672
rect 41564 4632 41570 4644
rect 41601 4641 41613 4644
rect 41647 4641 41659 4675
rect 43990 4672 43996 4684
rect 43951 4644 43996 4672
rect 41601 4635 41659 4641
rect 43990 4632 43996 4644
rect 44048 4632 44054 4684
rect 44542 4632 44548 4684
rect 44600 4672 44606 4684
rect 44637 4675 44695 4681
rect 44637 4672 44649 4675
rect 44600 4644 44649 4672
rect 44600 4632 44606 4644
rect 44637 4641 44649 4644
rect 44683 4641 44695 4675
rect 44637 4635 44695 4641
rect 45830 4632 45836 4684
rect 45888 4672 45894 4684
rect 46201 4675 46259 4681
rect 46201 4672 46213 4675
rect 45888 4644 46213 4672
rect 45888 4632 45894 4644
rect 46201 4641 46213 4644
rect 46247 4641 46259 4675
rect 47026 4672 47032 4684
rect 46987 4644 47032 4672
rect 46201 4635 46259 4641
rect 47026 4632 47032 4644
rect 47084 4632 47090 4684
rect 47578 4632 47584 4684
rect 47636 4672 47642 4684
rect 47673 4675 47731 4681
rect 47673 4672 47685 4675
rect 47636 4644 47685 4672
rect 47636 4632 47642 4644
rect 47673 4641 47685 4644
rect 47719 4641 47731 4675
rect 47673 4635 47731 4641
rect 49234 4632 49240 4684
rect 49292 4672 49298 4684
rect 52362 4672 52368 4684
rect 49292 4644 52368 4672
rect 49292 4632 49298 4644
rect 52362 4632 52368 4644
rect 52420 4632 52426 4684
rect 52546 4672 52552 4684
rect 52507 4644 52552 4672
rect 52546 4632 52552 4644
rect 52604 4632 52610 4684
rect 53466 4672 53472 4684
rect 53427 4644 53472 4672
rect 53466 4632 53472 4644
rect 53524 4632 53530 4684
rect 53650 4672 53656 4684
rect 53611 4644 53656 4672
rect 53650 4632 53656 4644
rect 53708 4632 53714 4684
rect 53837 4675 53895 4681
rect 53837 4641 53849 4675
rect 53883 4672 53895 4675
rect 54113 4675 54171 4681
rect 54113 4672 54125 4675
rect 53883 4644 54125 4672
rect 53883 4641 53895 4644
rect 53837 4635 53895 4641
rect 54113 4641 54125 4644
rect 54159 4641 54171 4675
rect 54294 4672 54300 4684
rect 54255 4644 54300 4672
rect 54113 4635 54171 4641
rect 54294 4632 54300 4644
rect 54352 4632 54358 4684
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4604 5043 4607
rect 6178 4604 6184 4616
rect 5031 4576 6184 4604
rect 5031 4573 5043 4576
rect 4985 4567 5043 4573
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 21174 4604 21180 4616
rect 8352 4576 21180 4604
rect 8352 4564 8358 4576
rect 21174 4564 21180 4576
rect 21232 4564 21238 4616
rect 26145 4607 26203 4613
rect 26145 4573 26157 4607
rect 26191 4573 26203 4607
rect 36446 4604 36452 4616
rect 26145 4567 26203 4573
rect 26712 4576 36452 4604
rect 1670 4496 1676 4548
rect 1728 4536 1734 4548
rect 2685 4539 2743 4545
rect 2685 4536 2697 4539
rect 1728 4508 2697 4536
rect 1728 4496 1734 4508
rect 2685 4505 2697 4508
rect 2731 4505 2743 4539
rect 7098 4536 7104 4548
rect 7059 4508 7104 4536
rect 2685 4499 2743 4505
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 7374 4496 7380 4548
rect 7432 4536 7438 4548
rect 8113 4539 8171 4545
rect 8113 4536 8125 4539
rect 7432 4508 8125 4536
rect 7432 4496 7438 4508
rect 8113 4505 8125 4508
rect 8159 4505 8171 4539
rect 8113 4499 8171 4505
rect 19978 4496 19984 4548
rect 20036 4536 20042 4548
rect 22830 4536 22836 4548
rect 20036 4508 22836 4536
rect 20036 4496 20042 4508
rect 22830 4496 22836 4508
rect 22888 4496 22894 4548
rect 26160 4536 26188 4567
rect 26712 4536 26740 4576
rect 36446 4564 36452 4576
rect 36504 4564 36510 4616
rect 37369 4607 37427 4613
rect 37369 4573 37381 4607
rect 37415 4604 37427 4607
rect 37734 4604 37740 4616
rect 37415 4576 37740 4604
rect 37415 4573 37427 4576
rect 37369 4567 37427 4573
rect 37734 4564 37740 4576
rect 37792 4564 37798 4616
rect 49510 4564 49516 4616
rect 49568 4604 49574 4616
rect 54404 4604 54432 4712
rect 55122 4700 55128 4752
rect 55180 4740 55186 4752
rect 62022 4740 62028 4752
rect 55180 4712 62028 4740
rect 55180 4700 55186 4712
rect 62022 4700 62028 4712
rect 62080 4700 62086 4752
rect 62390 4740 62396 4752
rect 62132 4712 62396 4740
rect 55306 4632 55312 4684
rect 55364 4672 55370 4684
rect 57330 4672 57336 4684
rect 55364 4644 57336 4672
rect 55364 4632 55370 4644
rect 57330 4632 57336 4644
rect 57388 4632 57394 4684
rect 61838 4632 61844 4684
rect 61896 4672 61902 4684
rect 62132 4681 62160 4712
rect 62390 4700 62396 4712
rect 62448 4700 62454 4752
rect 65613 4743 65671 4749
rect 65613 4709 65625 4743
rect 65659 4740 65671 4743
rect 66162 4740 66168 4752
rect 65659 4712 66168 4740
rect 65659 4709 65671 4712
rect 65613 4703 65671 4709
rect 66162 4700 66168 4712
rect 66220 4700 66226 4752
rect 71038 4700 71044 4752
rect 71096 4740 71102 4752
rect 78214 4740 78220 4752
rect 71096 4712 78076 4740
rect 78175 4712 78220 4740
rect 71096 4700 71102 4712
rect 61933 4675 61991 4681
rect 61933 4672 61945 4675
rect 61896 4644 61945 4672
rect 61896 4632 61902 4644
rect 61933 4641 61945 4644
rect 61979 4641 61991 4675
rect 61933 4635 61991 4641
rect 62116 4675 62174 4681
rect 62116 4641 62128 4675
rect 62162 4641 62174 4675
rect 62298 4672 62304 4684
rect 62259 4644 62304 4672
rect 62116 4635 62174 4641
rect 62298 4632 62304 4644
rect 62356 4632 62362 4684
rect 62485 4675 62543 4681
rect 62485 4641 62497 4675
rect 62531 4672 62543 4675
rect 62574 4672 62580 4684
rect 62531 4644 62580 4672
rect 62531 4641 62543 4644
rect 62485 4635 62543 4641
rect 62574 4632 62580 4644
rect 62632 4632 62638 4684
rect 64230 4672 64236 4684
rect 64191 4644 64236 4672
rect 64230 4632 64236 4644
rect 64288 4632 64294 4684
rect 64322 4632 64328 4684
rect 64380 4672 64386 4684
rect 65426 4672 65432 4684
rect 64380 4644 65432 4672
rect 64380 4632 64386 4644
rect 65426 4632 65432 4644
rect 65484 4632 65490 4684
rect 65978 4632 65984 4684
rect 66036 4672 66042 4684
rect 66073 4675 66131 4681
rect 66073 4672 66085 4675
rect 66036 4644 66085 4672
rect 66036 4632 66042 4644
rect 66073 4641 66085 4644
rect 66119 4641 66131 4675
rect 68370 4672 68376 4684
rect 68331 4644 68376 4672
rect 66073 4635 66131 4641
rect 68370 4632 68376 4644
rect 68428 4632 68434 4684
rect 70762 4672 70768 4684
rect 70723 4644 70768 4672
rect 70762 4632 70768 4644
rect 70820 4632 70826 4684
rect 73798 4672 73804 4684
rect 73759 4644 73804 4672
rect 73798 4632 73804 4644
rect 73856 4632 73862 4684
rect 76282 4672 76288 4684
rect 76243 4644 76288 4672
rect 76282 4632 76288 4644
rect 76340 4632 76346 4684
rect 77938 4672 77944 4684
rect 77899 4644 77944 4672
rect 77938 4632 77944 4644
rect 77996 4632 78002 4684
rect 78048 4672 78076 4712
rect 78214 4700 78220 4712
rect 78272 4700 78278 4752
rect 78324 4740 78352 4780
rect 78398 4768 78404 4820
rect 78456 4808 78462 4820
rect 97534 4808 97540 4820
rect 78456 4780 97540 4808
rect 78456 4768 78462 4780
rect 97534 4768 97540 4780
rect 97592 4768 97598 4820
rect 78324 4712 84148 4740
rect 78125 4675 78183 4681
rect 78125 4672 78137 4675
rect 78048 4644 78137 4672
rect 78125 4641 78137 4644
rect 78171 4641 78183 4675
rect 78674 4672 78680 4684
rect 78635 4644 78680 4672
rect 78125 4635 78183 4641
rect 78674 4632 78680 4644
rect 78732 4632 78738 4684
rect 78766 4632 78772 4684
rect 78824 4672 78830 4684
rect 79321 4675 79379 4681
rect 79321 4672 79333 4675
rect 78824 4644 79333 4672
rect 78824 4632 78830 4644
rect 79321 4641 79333 4644
rect 79367 4641 79379 4675
rect 79321 4635 79379 4641
rect 79410 4632 79416 4684
rect 79468 4672 79474 4684
rect 79965 4675 80023 4681
rect 79965 4672 79977 4675
rect 79468 4644 79977 4672
rect 79468 4632 79474 4644
rect 79965 4641 79977 4644
rect 80011 4641 80023 4675
rect 79965 4635 80023 4641
rect 80054 4632 80060 4684
rect 80112 4672 80118 4684
rect 80609 4675 80667 4681
rect 80609 4672 80621 4675
rect 80112 4644 80621 4672
rect 80112 4632 80118 4644
rect 80609 4641 80621 4644
rect 80655 4641 80667 4675
rect 80609 4635 80667 4641
rect 81253 4675 81311 4681
rect 81253 4641 81265 4675
rect 81299 4641 81311 4675
rect 82906 4672 82912 4684
rect 82867 4644 82912 4672
rect 81253 4635 81311 4641
rect 61010 4604 61016 4616
rect 49568 4576 54340 4604
rect 54404 4576 61016 4604
rect 49568 4564 49574 4576
rect 52086 4536 52092 4548
rect 26160 4508 26740 4536
rect 26896 4508 37320 4536
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 26896 4468 26924 4508
rect 28626 4468 28632 4480
rect 8260 4440 26924 4468
rect 28587 4440 28632 4468
rect 8260 4428 8266 4440
rect 28626 4428 28632 4440
rect 28684 4428 28690 4480
rect 33042 4428 33048 4480
rect 33100 4468 33106 4480
rect 36814 4468 36820 4480
rect 33100 4440 36820 4468
rect 33100 4428 33106 4440
rect 36814 4428 36820 4440
rect 36872 4428 36878 4480
rect 37292 4468 37320 4508
rect 38304 4508 52092 4536
rect 38304 4468 38332 4508
rect 52086 4496 52092 4508
rect 52144 4496 52150 4548
rect 54205 4539 54263 4545
rect 54205 4536 54217 4539
rect 53392 4508 54217 4536
rect 37292 4440 38332 4468
rect 42150 4428 42156 4480
rect 42208 4468 42214 4480
rect 42797 4471 42855 4477
rect 42797 4468 42809 4471
rect 42208 4440 42809 4468
rect 42208 4428 42214 4440
rect 42797 4437 42809 4440
rect 42843 4437 42855 4471
rect 42797 4431 42855 4437
rect 46382 4428 46388 4480
rect 46440 4468 46446 4480
rect 53392 4468 53420 4508
rect 54205 4505 54217 4508
rect 54251 4505 54263 4539
rect 54312 4536 54340 4576
rect 61010 4564 61016 4576
rect 61068 4564 61074 4616
rect 62209 4607 62267 4613
rect 62209 4604 62221 4607
rect 62132 4576 62221 4604
rect 62132 4548 62160 4576
rect 62209 4573 62221 4576
rect 62255 4573 62267 4607
rect 62209 4567 62267 4573
rect 63497 4607 63555 4613
rect 63497 4573 63509 4607
rect 63543 4604 63555 4607
rect 63862 4604 63868 4616
rect 63543 4576 63868 4604
rect 63543 4573 63555 4576
rect 63497 4567 63555 4573
rect 63862 4564 63868 4576
rect 63920 4564 63926 4616
rect 63957 4607 64015 4613
rect 63957 4573 63969 4607
rect 64003 4573 64015 4607
rect 63957 4567 64015 4573
rect 58250 4536 58256 4548
rect 54312 4508 58256 4536
rect 54205 4499 54263 4505
rect 58250 4496 58256 4508
rect 58308 4496 58314 4548
rect 62114 4496 62120 4548
rect 62172 4496 62178 4548
rect 62850 4496 62856 4548
rect 62908 4536 62914 4548
rect 63972 4536 64000 4567
rect 64414 4564 64420 4616
rect 64472 4604 64478 4616
rect 64472 4576 77892 4604
rect 64472 4564 64478 4576
rect 62908 4508 64000 4536
rect 62908 4496 62914 4508
rect 64966 4496 64972 4548
rect 65024 4536 65030 4548
rect 77757 4539 77815 4545
rect 77757 4536 77769 4539
rect 65024 4508 77769 4536
rect 65024 4496 65030 4508
rect 77757 4505 77769 4508
rect 77803 4505 77815 4539
rect 77864 4536 77892 4576
rect 78950 4564 78956 4616
rect 79008 4604 79014 4616
rect 79008 4576 80468 4604
rect 79008 4564 79014 4576
rect 78398 4536 78404 4548
rect 77864 4508 78404 4536
rect 77757 4499 77815 4505
rect 78398 4496 78404 4508
rect 78456 4496 78462 4548
rect 80440 4536 80468 4576
rect 80514 4564 80520 4616
rect 80572 4604 80578 4616
rect 81268 4604 81296 4635
rect 82906 4632 82912 4644
rect 82964 4632 82970 4684
rect 83550 4672 83556 4684
rect 83511 4644 83556 4672
rect 83550 4632 83556 4644
rect 83608 4632 83614 4684
rect 80572 4576 81296 4604
rect 84120 4604 84148 4712
rect 84286 4700 84292 4752
rect 84344 4740 84350 4752
rect 85482 4740 85488 4752
rect 84344 4712 85488 4740
rect 84344 4700 84350 4712
rect 85482 4700 85488 4712
rect 85540 4740 85546 4752
rect 87598 4740 87604 4752
rect 85540 4712 87604 4740
rect 85540 4700 85546 4712
rect 87598 4700 87604 4712
rect 87656 4700 87662 4752
rect 85390 4672 85396 4684
rect 85351 4644 85396 4672
rect 85390 4632 85396 4644
rect 85448 4632 85454 4684
rect 86034 4672 86040 4684
rect 85995 4644 86040 4672
rect 86034 4632 86040 4644
rect 86092 4632 86098 4684
rect 86954 4632 86960 4684
rect 87012 4672 87018 4684
rect 88153 4675 88211 4681
rect 88153 4672 88165 4675
rect 87012 4644 88165 4672
rect 87012 4632 87018 4644
rect 88153 4641 88165 4644
rect 88199 4641 88211 4675
rect 88794 4672 88800 4684
rect 88755 4644 88800 4672
rect 88153 4635 88211 4641
rect 88794 4632 88800 4644
rect 88852 4632 88858 4684
rect 89070 4632 89076 4684
rect 89128 4672 89134 4684
rect 89441 4675 89499 4681
rect 89441 4672 89453 4675
rect 89128 4644 89453 4672
rect 89128 4632 89134 4644
rect 89441 4641 89453 4644
rect 89487 4641 89499 4675
rect 89441 4635 89499 4641
rect 89714 4632 89720 4684
rect 89772 4672 89778 4684
rect 90085 4675 90143 4681
rect 90085 4672 90097 4675
rect 89772 4644 90097 4672
rect 89772 4632 89778 4644
rect 90085 4641 90097 4644
rect 90131 4641 90143 4675
rect 90085 4635 90143 4641
rect 90266 4632 90272 4684
rect 90324 4672 90330 4684
rect 90729 4675 90787 4681
rect 90729 4672 90741 4675
rect 90324 4644 90741 4672
rect 90324 4632 90330 4644
rect 90729 4641 90741 4644
rect 90775 4641 90787 4675
rect 90729 4635 90787 4641
rect 91094 4632 91100 4684
rect 91152 4672 91158 4684
rect 91373 4675 91431 4681
rect 91373 4672 91385 4675
rect 91152 4644 91385 4672
rect 91152 4632 91158 4644
rect 91373 4641 91385 4644
rect 91419 4641 91431 4675
rect 91373 4635 91431 4641
rect 91646 4632 91652 4684
rect 91704 4672 91710 4684
rect 92017 4675 92075 4681
rect 92017 4672 92029 4675
rect 91704 4644 92029 4672
rect 91704 4632 91710 4644
rect 92017 4641 92029 4644
rect 92063 4641 92075 4675
rect 92017 4635 92075 4641
rect 92750 4632 92756 4684
rect 92808 4672 92814 4684
rect 93397 4675 93455 4681
rect 93397 4672 93409 4675
rect 92808 4644 93409 4672
rect 92808 4632 92814 4644
rect 93397 4641 93409 4644
rect 93443 4641 93455 4675
rect 93397 4635 93455 4641
rect 93854 4632 93860 4684
rect 93912 4672 93918 4684
rect 94041 4675 94099 4681
rect 94041 4672 94053 4675
rect 93912 4644 94053 4672
rect 93912 4632 93918 4644
rect 94041 4641 94053 4644
rect 94087 4641 94099 4675
rect 94041 4635 94099 4641
rect 94222 4632 94228 4684
rect 94280 4672 94286 4684
rect 94685 4675 94743 4681
rect 94685 4672 94697 4675
rect 94280 4644 94697 4672
rect 94280 4632 94286 4644
rect 94685 4641 94697 4644
rect 94731 4641 94743 4675
rect 95326 4672 95332 4684
rect 95287 4644 95332 4672
rect 94685 4635 94743 4641
rect 95326 4632 95332 4644
rect 95384 4632 95390 4684
rect 95970 4672 95976 4684
rect 95931 4644 95976 4672
rect 95970 4632 95976 4644
rect 96028 4632 96034 4684
rect 96617 4675 96675 4681
rect 96617 4641 96629 4675
rect 96663 4672 96675 4675
rect 96706 4672 96712 4684
rect 96663 4644 96712 4672
rect 96663 4641 96675 4644
rect 96617 4635 96675 4641
rect 96706 4632 96712 4644
rect 96764 4632 96770 4684
rect 97258 4672 97264 4684
rect 97219 4644 97264 4672
rect 97258 4632 97264 4644
rect 97316 4632 97322 4684
rect 88334 4604 88340 4616
rect 84120 4576 88340 4604
rect 80572 4564 80578 4576
rect 88334 4564 88340 4576
rect 88392 4564 88398 4616
rect 90726 4536 90732 4548
rect 80440 4508 90732 4536
rect 90726 4496 90732 4508
rect 90784 4496 90790 4548
rect 46440 4440 53420 4468
rect 46440 4428 46446 4440
rect 53466 4428 53472 4480
rect 53524 4468 53530 4480
rect 62022 4468 62028 4480
rect 53524 4440 62028 4468
rect 53524 4428 53530 4440
rect 62022 4428 62028 4440
rect 62080 4428 62086 4480
rect 62298 4428 62304 4480
rect 62356 4468 62362 4480
rect 62577 4471 62635 4477
rect 62577 4468 62589 4471
rect 62356 4440 62589 4468
rect 62356 4428 62362 4440
rect 62577 4437 62589 4440
rect 62623 4437 62635 4471
rect 62577 4431 62635 4437
rect 67634 4428 67640 4480
rect 67692 4468 67698 4480
rect 74166 4468 74172 4480
rect 67692 4440 74172 4468
rect 67692 4428 67698 4440
rect 74166 4428 74172 4440
rect 74224 4428 74230 4480
rect 87049 4471 87107 4477
rect 87049 4437 87061 4471
rect 87095 4468 87107 4471
rect 89346 4468 89352 4480
rect 87095 4440 89352 4468
rect 87095 4437 87107 4440
rect 87049 4431 87107 4437
rect 89346 4428 89352 4440
rect 89404 4428 89410 4480
rect 1104 4378 98808 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 65686 4378
rect 65738 4326 65750 4378
rect 65802 4326 65814 4378
rect 65866 4326 65878 4378
rect 65930 4326 96406 4378
rect 96458 4326 96470 4378
rect 96522 4326 96534 4378
rect 96586 4326 96598 4378
rect 96650 4326 98808 4378
rect 1104 4304 98808 4326
rect 15304 4236 16252 4264
rect 3789 4199 3847 4205
rect 3789 4165 3801 4199
rect 3835 4165 3847 4199
rect 3789 4159 3847 4165
rect 2958 4128 2964 4140
rect 2919 4100 2964 4128
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3804 4128 3832 4159
rect 5258 4128 5264 4140
rect 3804 4100 5264 4128
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 7098 4128 7104 4140
rect 6236 4100 7104 4128
rect 6236 4088 6242 4100
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 15304 4128 15332 4236
rect 8588 4100 15332 4128
rect 15396 4168 16160 4196
rect 1210 4020 1216 4072
rect 1268 4060 1274 4072
rect 2685 4063 2743 4069
rect 2685 4060 2697 4063
rect 1268 4032 2697 4060
rect 1268 4020 1274 4032
rect 2685 4029 2697 4032
rect 2731 4029 2743 4063
rect 2685 4023 2743 4029
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 3200 4032 3617 4060
rect 3200 4020 3206 4032
rect 3605 4029 3617 4032
rect 3651 4029 3663 4063
rect 4706 4060 4712 4072
rect 4667 4032 4712 4060
rect 3605 4023 3663 4029
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 5442 4060 5448 4072
rect 4908 4032 5448 4060
rect 658 3952 664 4004
rect 716 3992 722 4004
rect 1857 3995 1915 4001
rect 1857 3992 1869 3995
rect 716 3964 1869 3992
rect 716 3952 722 3964
rect 1857 3961 1869 3964
rect 1903 3961 1915 3995
rect 2222 3992 2228 4004
rect 2183 3964 2228 3992
rect 1857 3955 1915 3961
rect 2222 3952 2228 3964
rect 2280 3952 2286 4004
rect 3326 3952 3332 4004
rect 3384 3992 3390 4004
rect 4341 3995 4399 4001
rect 3384 3964 3924 3992
rect 3384 3952 3390 3964
rect 3896 3924 3924 3964
rect 4341 3961 4353 3995
rect 4387 3992 4399 3995
rect 4908 3992 4936 4032
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 6546 4020 6552 4072
rect 6604 4060 6610 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6604 4032 6837 4060
rect 6604 4020 6610 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 7742 4060 7748 4072
rect 7703 4032 7748 4060
rect 6825 4023 6883 4029
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 4387 3964 4936 3992
rect 4985 3995 5043 4001
rect 4387 3961 4399 3964
rect 4341 3955 4399 3961
rect 4985 3961 4997 3995
rect 5031 3992 5043 3995
rect 5258 3992 5264 4004
rect 5031 3964 5264 3992
rect 5031 3961 5043 3964
rect 4985 3955 5043 3961
rect 5258 3952 5264 3964
rect 5316 3952 5322 4004
rect 5721 3995 5779 4001
rect 5721 3961 5733 3995
rect 5767 3992 5779 3995
rect 8588 3992 8616 4100
rect 9398 4060 9404 4072
rect 9359 4032 9404 4060
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 9548 4032 10057 4060
rect 9548 4020 9554 4032
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 10689 4063 10747 4069
rect 10689 4060 10701 4063
rect 10192 4032 10701 4060
rect 10192 4020 10198 4032
rect 10689 4029 10701 4032
rect 10735 4029 10747 4063
rect 10689 4023 10747 4029
rect 11422 4020 11428 4072
rect 11480 4060 11486 4072
rect 12345 4063 12403 4069
rect 12345 4060 12357 4063
rect 11480 4032 12357 4060
rect 11480 4020 11486 4032
rect 12345 4029 12357 4032
rect 12391 4029 12403 4063
rect 12345 4023 12403 4029
rect 12897 4063 12955 4069
rect 12897 4029 12909 4063
rect 12943 4060 12955 4063
rect 13170 4060 13176 4072
rect 12943 4032 13176 4060
rect 12943 4029 12955 4032
rect 12897 4023 12955 4029
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 5767 3964 8616 3992
rect 8665 3995 8723 4001
rect 5767 3961 5779 3964
rect 5721 3955 5779 3961
rect 8665 3961 8677 3995
rect 8711 3992 8723 3995
rect 8711 3964 13032 3992
rect 8711 3961 8723 3964
rect 8665 3955 8723 3961
rect 4433 3927 4491 3933
rect 4433 3924 4445 3927
rect 3896 3896 4445 3924
rect 4433 3893 4445 3896
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 5813 3927 5871 3933
rect 5813 3924 5825 3927
rect 5132 3896 5825 3924
rect 5132 3884 5138 3896
rect 5813 3893 5825 3896
rect 5859 3893 5871 3927
rect 7006 3924 7012 3936
rect 6967 3896 7012 3924
rect 5813 3887 5871 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 7834 3884 7840 3936
rect 7892 3924 7898 3936
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 7892 3896 7941 3924
rect 7892 3884 7898 3896
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 7929 3887 7987 3893
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 8628 3896 8769 3924
rect 8628 3884 8634 3896
rect 8757 3893 8769 3896
rect 8803 3893 8815 3927
rect 8757 3887 8815 3893
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 8996 3896 9505 3924
rect 8996 3884 9002 3896
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 12437 3927 12495 3933
rect 12437 3924 12449 3927
rect 12308 3896 12449 3924
rect 12308 3884 12314 3896
rect 12437 3893 12449 3896
rect 12483 3893 12495 3927
rect 13004 3924 13032 3964
rect 13078 3952 13084 4004
rect 13136 3992 13142 4004
rect 13648 3992 13676 4023
rect 13722 4020 13728 4072
rect 13780 4060 13786 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 13780 4032 14289 4060
rect 13780 4020 13786 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 15396 4060 15424 4168
rect 14277 4023 14335 4029
rect 15212 4032 15424 4060
rect 13136 3964 13676 3992
rect 13136 3952 13142 3964
rect 15212 3924 15240 4032
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 16025 4063 16083 4069
rect 16025 4060 16037 4063
rect 15528 4032 16037 4060
rect 15528 4020 15534 4032
rect 16025 4029 16037 4032
rect 16071 4029 16083 4063
rect 16025 4023 16083 4029
rect 15381 3995 15439 4001
rect 15381 3961 15393 3995
rect 15427 3992 15439 3995
rect 16132 3992 16160 4168
rect 16224 4128 16252 4236
rect 33502 4224 33508 4276
rect 33560 4264 33566 4276
rect 46290 4264 46296 4276
rect 33560 4236 46296 4264
rect 33560 4224 33566 4236
rect 46290 4224 46296 4236
rect 46348 4224 46354 4276
rect 47946 4224 47952 4276
rect 48004 4264 48010 4276
rect 48004 4236 91876 4264
rect 48004 4224 48010 4236
rect 19981 4199 20039 4205
rect 19981 4165 19993 4199
rect 20027 4196 20039 4199
rect 21910 4196 21916 4208
rect 20027 4168 21916 4196
rect 20027 4165 20039 4168
rect 19981 4159 20039 4165
rect 21910 4156 21916 4168
rect 21968 4156 21974 4208
rect 33134 4156 33140 4208
rect 33192 4196 33198 4208
rect 33192 4168 42656 4196
rect 33192 4156 33198 4168
rect 34977 4131 35035 4137
rect 16224 4100 31754 4128
rect 16758 4020 16764 4072
rect 16816 4060 16822 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16816 4032 17325 4060
rect 16816 4020 16822 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 18322 4020 18328 4072
rect 18380 4060 18386 4072
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 18380 4032 18429 4060
rect 18380 4020 18386 4032
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 19242 4020 19248 4072
rect 19300 4060 19306 4072
rect 20441 4063 20499 4069
rect 20441 4060 20453 4063
rect 19300 4032 20453 4060
rect 19300 4020 19306 4032
rect 20441 4029 20453 4032
rect 20487 4029 20499 4063
rect 20441 4023 20499 4029
rect 21085 4063 21143 4069
rect 21085 4029 21097 4063
rect 21131 4029 21143 4063
rect 23014 4060 23020 4072
rect 22975 4032 23020 4060
rect 21085 4023 21143 4029
rect 18782 3992 18788 4004
rect 15427 3964 16068 3992
rect 16132 3964 18788 3992
rect 15427 3961 15439 3964
rect 15381 3955 15439 3961
rect 16040 3936 16068 3964
rect 18782 3952 18788 3964
rect 18840 3952 18846 4004
rect 19150 3992 19156 4004
rect 19111 3964 19156 3992
rect 19150 3952 19156 3964
rect 19208 3952 19214 4004
rect 20346 3952 20352 4004
rect 20404 3992 20410 4004
rect 21100 3992 21128 4023
rect 23014 4020 23020 4032
rect 23072 4020 23078 4072
rect 23474 4060 23480 4072
rect 23435 4032 23480 4060
rect 23474 4020 23480 4032
rect 23532 4020 23538 4072
rect 23842 4020 23848 4072
rect 23900 4060 23906 4072
rect 24397 4063 24455 4069
rect 24397 4060 24409 4063
rect 23900 4032 24409 4060
rect 23900 4020 23906 4032
rect 24397 4029 24409 4032
rect 24443 4029 24455 4063
rect 24397 4023 24455 4029
rect 24486 4020 24492 4072
rect 24544 4060 24550 4072
rect 25041 4063 25099 4069
rect 25041 4060 25053 4063
rect 24544 4032 25053 4060
rect 24544 4020 24550 4032
rect 25041 4029 25053 4032
rect 25087 4029 25099 4063
rect 25041 4023 25099 4029
rect 25593 4063 25651 4069
rect 25593 4029 25605 4063
rect 25639 4060 25651 4063
rect 25869 4063 25927 4069
rect 25869 4060 25881 4063
rect 25639 4032 25881 4060
rect 25639 4029 25651 4032
rect 25593 4023 25651 4029
rect 25869 4029 25881 4032
rect 25915 4060 25927 4063
rect 25958 4060 25964 4072
rect 25915 4032 25964 4060
rect 25915 4029 25927 4032
rect 25869 4023 25927 4029
rect 25958 4020 25964 4032
rect 26016 4020 26022 4072
rect 26329 4063 26387 4069
rect 26329 4029 26341 4063
rect 26375 4029 26387 4063
rect 26329 4023 26387 4029
rect 25314 3992 25320 4004
rect 20404 3964 21128 3992
rect 22066 3964 25320 3992
rect 20404 3952 20410 3964
rect 13004 3896 15240 3924
rect 12437 3887 12495 3893
rect 15286 3884 15292 3936
rect 15344 3924 15350 3936
rect 15473 3927 15531 3933
rect 15473 3924 15485 3927
rect 15344 3896 15485 3924
rect 15344 3884 15350 3896
rect 15473 3893 15485 3896
rect 15519 3893 15531 3927
rect 15473 3887 15531 3893
rect 16022 3884 16028 3936
rect 16080 3884 16086 3936
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 18509 3927 18567 3933
rect 18509 3924 18521 3927
rect 18380 3896 18521 3924
rect 18380 3884 18386 3896
rect 18509 3893 18521 3896
rect 18555 3893 18567 3927
rect 18509 3887 18567 3893
rect 18966 3884 18972 3936
rect 19024 3924 19030 3936
rect 19245 3927 19303 3933
rect 19245 3924 19257 3927
rect 19024 3896 19257 3924
rect 19024 3884 19030 3896
rect 19245 3893 19257 3896
rect 19291 3893 19303 3927
rect 19245 3887 19303 3893
rect 19334 3884 19340 3936
rect 19392 3924 19398 3936
rect 22066 3924 22094 3964
rect 25314 3952 25320 3964
rect 25372 3952 25378 4004
rect 25774 3952 25780 4004
rect 25832 3992 25838 4004
rect 26344 3992 26372 4023
rect 26510 4020 26516 4072
rect 26568 4060 26574 4072
rect 27801 4063 27859 4069
rect 27801 4060 27813 4063
rect 26568 4032 27813 4060
rect 26568 4020 26574 4032
rect 27801 4029 27813 4032
rect 27847 4029 27859 4063
rect 27801 4023 27859 4029
rect 28074 4020 28080 4072
rect 28132 4060 28138 4072
rect 28445 4063 28503 4069
rect 28445 4060 28457 4063
rect 28132 4032 28457 4060
rect 28132 4020 28138 4032
rect 28445 4029 28457 4032
rect 28491 4029 28503 4063
rect 28445 4023 28503 4029
rect 28718 4020 28724 4072
rect 28776 4060 28782 4072
rect 29089 4063 29147 4069
rect 29089 4060 29101 4063
rect 28776 4032 29101 4060
rect 28776 4020 28782 4032
rect 29089 4029 29101 4032
rect 29135 4029 29147 4063
rect 29089 4023 29147 4029
rect 29362 4020 29368 4072
rect 29420 4060 29426 4072
rect 29733 4063 29791 4069
rect 29733 4060 29745 4063
rect 29420 4032 29745 4060
rect 29420 4020 29426 4032
rect 29733 4029 29745 4032
rect 29779 4029 29791 4063
rect 31202 4060 31208 4072
rect 31163 4032 31208 4060
rect 29733 4023 29791 4029
rect 31202 4020 31208 4032
rect 31260 4020 31266 4072
rect 25832 3964 26372 3992
rect 25832 3952 25838 3964
rect 26418 3952 26424 4004
rect 26476 3992 26482 4004
rect 29914 3992 29920 4004
rect 26476 3964 29920 3992
rect 26476 3952 26482 3964
rect 29914 3952 29920 3964
rect 29972 3952 29978 4004
rect 19392 3896 22094 3924
rect 19392 3884 19398 3896
rect 23382 3884 23388 3936
rect 23440 3924 23446 3936
rect 23477 3927 23535 3933
rect 23477 3924 23489 3927
rect 23440 3896 23489 3924
rect 23440 3884 23446 3896
rect 23477 3893 23489 3896
rect 23523 3893 23535 3927
rect 23477 3887 23535 3893
rect 26878 3884 26884 3936
rect 26936 3924 26942 3936
rect 27798 3924 27804 3936
rect 26936 3896 27804 3924
rect 26936 3884 26942 3896
rect 27798 3884 27804 3896
rect 27856 3884 27862 3936
rect 31726 3924 31754 4100
rect 34977 4097 34989 4131
rect 35023 4128 35035 4131
rect 35618 4128 35624 4140
rect 35023 4100 35624 4128
rect 35023 4097 35035 4100
rect 34977 4091 35035 4097
rect 35618 4088 35624 4100
rect 35676 4088 35682 4140
rect 37274 4088 37280 4140
rect 37332 4128 37338 4140
rect 37332 4100 39344 4128
rect 37332 4088 37338 4100
rect 32950 4020 32956 4072
rect 33008 4060 33014 4072
rect 33045 4063 33103 4069
rect 33045 4060 33057 4063
rect 33008 4032 33057 4060
rect 33008 4020 33014 4032
rect 33045 4029 33057 4032
rect 33091 4029 33103 4063
rect 33045 4023 33103 4029
rect 33594 4020 33600 4072
rect 33652 4060 33658 4072
rect 33689 4063 33747 4069
rect 33689 4060 33701 4063
rect 33652 4032 33701 4060
rect 33652 4020 33658 4032
rect 33689 4029 33701 4032
rect 33735 4029 33747 4063
rect 33689 4023 33747 4029
rect 34330 4020 34336 4072
rect 34388 4060 34394 4072
rect 34425 4063 34483 4069
rect 34425 4060 34437 4063
rect 34388 4032 34437 4060
rect 34388 4020 34394 4032
rect 34425 4029 34437 4032
rect 34471 4029 34483 4063
rect 34425 4023 34483 4029
rect 34790 4020 34796 4072
rect 34848 4060 34854 4072
rect 35529 4063 35587 4069
rect 35529 4060 35541 4063
rect 34848 4032 35541 4060
rect 34848 4020 34854 4032
rect 35529 4029 35541 4032
rect 35575 4029 35587 4063
rect 35529 4023 35587 4029
rect 35710 4020 35716 4072
rect 35768 4060 35774 4072
rect 36173 4063 36231 4069
rect 36173 4060 36185 4063
rect 35768 4032 36185 4060
rect 35768 4020 35774 4032
rect 36173 4029 36185 4032
rect 36219 4029 36231 4063
rect 36814 4060 36820 4072
rect 36775 4032 36820 4060
rect 36173 4023 36231 4029
rect 36814 4020 36820 4032
rect 36872 4020 36878 4072
rect 38654 4060 38660 4072
rect 38615 4032 38660 4060
rect 38654 4020 38660 4032
rect 38712 4020 38718 4072
rect 39316 4069 39344 4100
rect 39390 4088 39396 4140
rect 39448 4128 39454 4140
rect 39448 4100 40632 4128
rect 39448 4088 39454 4100
rect 39301 4063 39359 4069
rect 39301 4029 39313 4063
rect 39347 4029 39359 4063
rect 39942 4060 39948 4072
rect 39903 4032 39948 4060
rect 39301 4023 39359 4029
rect 39942 4020 39948 4032
rect 40000 4020 40006 4072
rect 40604 4069 40632 4100
rect 40589 4063 40647 4069
rect 40589 4029 40601 4063
rect 40635 4029 40647 4063
rect 41233 4063 41291 4069
rect 41233 4060 41245 4063
rect 40589 4023 40647 4029
rect 40696 4032 41245 4060
rect 38562 3952 38568 4004
rect 38620 3992 38626 4004
rect 39206 3992 39212 4004
rect 38620 3964 39212 3992
rect 38620 3952 38626 3964
rect 39206 3952 39212 3964
rect 39264 3952 39270 4004
rect 39666 3952 39672 4004
rect 39724 3992 39730 4004
rect 40696 3992 40724 4032
rect 41233 4029 41245 4032
rect 41279 4029 41291 4063
rect 41877 4063 41935 4069
rect 41877 4060 41889 4063
rect 41233 4023 41291 4029
rect 41386 4032 41889 4060
rect 39724 3964 40724 3992
rect 39724 3952 39730 3964
rect 40954 3952 40960 4004
rect 41012 3992 41018 4004
rect 41386 3992 41414 4032
rect 41877 4029 41889 4032
rect 41923 4029 41935 4063
rect 41877 4023 41935 4029
rect 41012 3964 41414 3992
rect 41012 3952 41018 3964
rect 36354 3924 36360 3936
rect 31726 3896 36360 3924
rect 36354 3884 36360 3896
rect 36412 3884 36418 3936
rect 36538 3884 36544 3936
rect 36596 3924 36602 3936
rect 42334 3924 42340 3936
rect 36596 3896 42340 3924
rect 36596 3884 36602 3896
rect 42334 3884 42340 3896
rect 42392 3884 42398 3936
rect 42628 3924 42656 4168
rect 42702 4156 42708 4208
rect 42760 4156 42766 4208
rect 48498 4156 48504 4208
rect 48556 4196 48562 4208
rect 86865 4199 86923 4205
rect 86865 4196 86877 4199
rect 48556 4168 86877 4196
rect 48556 4156 48562 4168
rect 86865 4165 86877 4168
rect 86911 4165 86923 4199
rect 86865 4159 86923 4165
rect 42720 4128 42748 4156
rect 55766 4128 55772 4140
rect 42720 4100 55772 4128
rect 55766 4088 55772 4100
rect 55824 4088 55830 4140
rect 60918 4128 60924 4140
rect 58544 4100 60924 4128
rect 42702 4020 42708 4072
rect 42760 4060 42766 4072
rect 43533 4063 43591 4069
rect 43533 4060 43545 4063
rect 42760 4032 43545 4060
rect 42760 4020 42766 4032
rect 43533 4029 43545 4032
rect 43579 4029 43591 4063
rect 43533 4023 43591 4029
rect 44177 4063 44235 4069
rect 44177 4029 44189 4063
rect 44223 4029 44235 4063
rect 45370 4060 45376 4072
rect 45331 4032 45376 4060
rect 44177 4023 44235 4029
rect 43346 3952 43352 4004
rect 43404 3992 43410 4004
rect 44192 3992 44220 4023
rect 45370 4020 45376 4032
rect 45428 4020 45434 4072
rect 46014 4060 46020 4072
rect 45975 4032 46020 4060
rect 46014 4020 46020 4032
rect 46072 4020 46078 4072
rect 46661 4063 46719 4069
rect 46661 4060 46673 4063
rect 46124 4032 46673 4060
rect 43404 3964 44220 3992
rect 43404 3952 43410 3964
rect 45186 3952 45192 4004
rect 45244 3992 45250 4004
rect 46124 3992 46152 4032
rect 46661 4029 46673 4032
rect 46707 4029 46719 4063
rect 46661 4023 46719 4029
rect 47305 4063 47363 4069
rect 47305 4029 47317 4063
rect 47351 4029 47363 4063
rect 47305 4023 47363 4029
rect 45244 3964 46152 3992
rect 45244 3952 45250 3964
rect 46382 3952 46388 4004
rect 46440 3992 46446 4004
rect 47320 3992 47348 4023
rect 48222 4020 48228 4072
rect 48280 4060 48286 4072
rect 48777 4063 48835 4069
rect 48777 4060 48789 4063
rect 48280 4032 48789 4060
rect 48280 4020 48286 4032
rect 48777 4029 48789 4032
rect 48823 4029 48835 4063
rect 48777 4023 48835 4029
rect 48866 4020 48872 4072
rect 48924 4060 48930 4072
rect 49421 4063 49479 4069
rect 49421 4060 49433 4063
rect 48924 4032 49433 4060
rect 48924 4020 48930 4032
rect 49421 4029 49433 4032
rect 49467 4029 49479 4063
rect 49421 4023 49479 4029
rect 49510 4020 49516 4072
rect 49568 4060 49574 4072
rect 50065 4063 50123 4069
rect 50065 4060 50077 4063
rect 49568 4032 50077 4060
rect 49568 4020 49574 4032
rect 50065 4029 50077 4032
rect 50111 4029 50123 4063
rect 50065 4023 50123 4029
rect 50154 4020 50160 4072
rect 50212 4060 50218 4072
rect 50709 4063 50767 4069
rect 50709 4060 50721 4063
rect 50212 4032 50721 4060
rect 50212 4020 50218 4032
rect 50709 4029 50721 4032
rect 50755 4029 50767 4063
rect 50709 4023 50767 4029
rect 50798 4020 50804 4072
rect 50856 4060 50862 4072
rect 51353 4063 51411 4069
rect 51353 4060 51365 4063
rect 50856 4032 51365 4060
rect 50856 4020 50862 4032
rect 51353 4029 51365 4032
rect 51399 4029 51411 4063
rect 51997 4063 52055 4069
rect 51997 4060 52009 4063
rect 51353 4023 51411 4029
rect 51460 4032 52009 4060
rect 46440 3964 47348 3992
rect 46440 3952 46446 3964
rect 51258 3952 51264 4004
rect 51316 3992 51322 4004
rect 51460 3992 51488 4032
rect 51997 4029 52009 4032
rect 52043 4029 52055 4063
rect 51997 4023 52055 4029
rect 52638 4020 52644 4072
rect 52696 4060 52702 4072
rect 52696 4032 52741 4060
rect 52696 4020 52702 4032
rect 53098 4020 53104 4072
rect 53156 4060 53162 4072
rect 54021 4063 54079 4069
rect 54021 4060 54033 4063
rect 53156 4032 54033 4060
rect 53156 4020 53162 4032
rect 54021 4029 54033 4032
rect 54067 4029 54079 4063
rect 54021 4023 54079 4029
rect 54665 4063 54723 4069
rect 54665 4029 54677 4063
rect 54711 4029 54723 4063
rect 54665 4023 54723 4029
rect 51316 3964 51488 3992
rect 51316 3952 51322 3964
rect 53650 3952 53656 4004
rect 53708 3992 53714 4004
rect 54680 3992 54708 4023
rect 54938 4020 54944 4072
rect 54996 4060 55002 4072
rect 55309 4063 55367 4069
rect 55309 4060 55321 4063
rect 54996 4032 55321 4060
rect 54996 4020 55002 4032
rect 55309 4029 55321 4032
rect 55355 4029 55367 4063
rect 55309 4023 55367 4029
rect 55582 4020 55588 4072
rect 55640 4060 55646 4072
rect 55953 4063 56011 4069
rect 55953 4060 55965 4063
rect 55640 4032 55965 4060
rect 55640 4020 55646 4032
rect 55953 4029 55965 4032
rect 55999 4029 56011 4063
rect 55953 4023 56011 4029
rect 56226 4020 56232 4072
rect 56284 4060 56290 4072
rect 56597 4063 56655 4069
rect 56597 4060 56609 4063
rect 56284 4032 56609 4060
rect 56284 4020 56290 4032
rect 56597 4029 56609 4032
rect 56643 4029 56655 4063
rect 56597 4023 56655 4029
rect 56778 4020 56784 4072
rect 56836 4060 56842 4072
rect 57241 4063 57299 4069
rect 57241 4060 57253 4063
rect 56836 4032 57253 4060
rect 56836 4020 56842 4032
rect 57241 4029 57253 4032
rect 57287 4029 57299 4063
rect 57241 4023 57299 4029
rect 57422 4020 57428 4072
rect 57480 4060 57486 4072
rect 57885 4063 57943 4069
rect 57885 4060 57897 4063
rect 57480 4032 57897 4060
rect 57480 4020 57486 4032
rect 57885 4029 57897 4032
rect 57931 4029 57943 4063
rect 57885 4023 57943 4029
rect 58544 3992 58572 4100
rect 60918 4088 60924 4100
rect 60976 4088 60982 4140
rect 61010 4088 61016 4140
rect 61068 4128 61074 4140
rect 61068 4100 61792 4128
rect 61068 4088 61074 4100
rect 58618 4020 58624 4072
rect 58676 4060 58682 4072
rect 59265 4063 59323 4069
rect 59265 4060 59277 4063
rect 58676 4032 59277 4060
rect 58676 4020 58682 4032
rect 59265 4029 59277 4032
rect 59311 4029 59323 4063
rect 59909 4063 59967 4069
rect 59909 4060 59921 4063
rect 59265 4023 59323 4029
rect 59372 4032 59921 4060
rect 53708 3964 54708 3992
rect 55140 3964 58572 3992
rect 53708 3952 53714 3964
rect 52822 3924 52828 3936
rect 42628 3896 52828 3924
rect 52822 3884 52828 3896
rect 52880 3884 52886 3936
rect 53926 3884 53932 3936
rect 53984 3924 53990 3936
rect 55140 3924 55168 3964
rect 59078 3952 59084 4004
rect 59136 3992 59142 4004
rect 59372 3992 59400 4032
rect 59909 4029 59921 4032
rect 59955 4029 59967 4063
rect 59909 4023 59967 4029
rect 60553 4063 60611 4069
rect 60553 4029 60565 4063
rect 60599 4029 60611 4063
rect 60553 4023 60611 4029
rect 59136 3964 59400 3992
rect 59136 3952 59142 3964
rect 59814 3952 59820 4004
rect 59872 3992 59878 4004
rect 60560 3992 60588 4023
rect 60734 4020 60740 4072
rect 60792 4060 60798 4072
rect 61197 4063 61255 4069
rect 61197 4060 61209 4063
rect 60792 4032 61209 4060
rect 60792 4020 60798 4032
rect 61197 4029 61209 4032
rect 61243 4029 61255 4063
rect 61764 4060 61792 4100
rect 62298 4088 62304 4140
rect 62356 4128 62362 4140
rect 62356 4100 63080 4128
rect 62356 4088 62362 4100
rect 61833 4063 61891 4069
rect 61833 4060 61845 4063
rect 61764 4032 61845 4060
rect 61197 4023 61255 4029
rect 61833 4029 61845 4032
rect 61879 4029 61891 4063
rect 61833 4023 61891 4029
rect 62022 4020 62028 4072
rect 62080 4060 62086 4072
rect 62485 4063 62543 4069
rect 62485 4060 62497 4063
rect 62080 4032 62497 4060
rect 62080 4020 62086 4032
rect 62485 4029 62497 4032
rect 62531 4029 62543 4063
rect 63052 4060 63080 4100
rect 63494 4088 63500 4140
rect 63552 4128 63558 4140
rect 63552 4100 64644 4128
rect 63552 4088 63558 4100
rect 63121 4063 63179 4069
rect 63121 4060 63133 4063
rect 63052 4032 63133 4060
rect 62485 4023 62543 4029
rect 63121 4029 63133 4032
rect 63167 4029 63179 4063
rect 63121 4023 63179 4029
rect 63218 4020 63224 4072
rect 63276 4060 63282 4072
rect 64509 4063 64567 4069
rect 64509 4060 64521 4063
rect 63276 4032 64521 4060
rect 63276 4020 63282 4032
rect 64509 4029 64521 4032
rect 64555 4029 64567 4063
rect 64616 4060 64644 4100
rect 64782 4088 64788 4140
rect 64840 4128 64846 4140
rect 64840 4100 65288 4128
rect 64840 4088 64846 4100
rect 65153 4063 65211 4069
rect 65153 4060 65165 4063
rect 64616 4032 65165 4060
rect 64509 4023 64567 4029
rect 65153 4029 65165 4032
rect 65199 4029 65211 4063
rect 65260 4060 65288 4100
rect 65334 4088 65340 4140
rect 65392 4128 65398 4140
rect 65392 4100 66484 4128
rect 65392 4088 65398 4100
rect 66456 4069 66484 4100
rect 69566 4088 69572 4140
rect 69624 4128 69630 4140
rect 69624 4100 69888 4128
rect 69624 4088 69630 4100
rect 65797 4063 65855 4069
rect 65797 4060 65809 4063
rect 65260 4032 65809 4060
rect 65153 4023 65211 4029
rect 65797 4029 65809 4032
rect 65843 4029 65855 4063
rect 65797 4023 65855 4029
rect 66441 4063 66499 4069
rect 66441 4029 66453 4063
rect 66487 4029 66499 4063
rect 66441 4023 66499 4029
rect 66530 4020 66536 4072
rect 66588 4060 66594 4072
rect 67085 4063 67143 4069
rect 67085 4060 67097 4063
rect 66588 4032 67097 4060
rect 66588 4020 66594 4032
rect 67085 4029 67097 4032
rect 67131 4029 67143 4063
rect 67085 4023 67143 4029
rect 67174 4020 67180 4072
rect 67232 4060 67238 4072
rect 67729 4063 67787 4069
rect 67729 4060 67741 4063
rect 67232 4032 67741 4060
rect 67232 4020 67238 4032
rect 67729 4029 67741 4032
rect 67775 4029 67787 4063
rect 67729 4023 67787 4029
rect 67818 4020 67824 4072
rect 67876 4060 67882 4072
rect 68373 4063 68431 4069
rect 68373 4060 68385 4063
rect 67876 4032 68385 4060
rect 67876 4020 67882 4032
rect 68373 4029 68385 4032
rect 68419 4029 68431 4063
rect 68373 4023 68431 4029
rect 68922 4020 68928 4072
rect 68980 4060 68986 4072
rect 69753 4063 69811 4069
rect 69753 4060 69765 4063
rect 68980 4032 69765 4060
rect 68980 4020 68986 4032
rect 69753 4029 69765 4032
rect 69799 4029 69811 4063
rect 69860 4060 69888 4100
rect 70210 4088 70216 4140
rect 70268 4128 70274 4140
rect 70268 4100 71084 4128
rect 70268 4088 70274 4100
rect 71056 4069 71084 4100
rect 87138 4088 87144 4140
rect 87196 4128 87202 4140
rect 88153 4131 88211 4137
rect 88153 4128 88165 4131
rect 87196 4100 88165 4128
rect 87196 4088 87202 4100
rect 88153 4097 88165 4100
rect 88199 4097 88211 4131
rect 88153 4091 88211 4097
rect 90634 4088 90640 4140
rect 90692 4128 90698 4140
rect 91848 4137 91876 4236
rect 91833 4131 91891 4137
rect 90692 4100 91600 4128
rect 90692 4088 90698 4100
rect 70397 4063 70455 4069
rect 70397 4060 70409 4063
rect 69860 4032 70409 4060
rect 69753 4023 69811 4029
rect 70397 4029 70409 4032
rect 70443 4029 70455 4063
rect 70397 4023 70455 4029
rect 71041 4063 71099 4069
rect 71041 4029 71053 4063
rect 71087 4029 71099 4063
rect 71041 4023 71099 4029
rect 71406 4020 71412 4072
rect 71464 4060 71470 4072
rect 71685 4063 71743 4069
rect 71685 4060 71697 4063
rect 71464 4032 71697 4060
rect 71464 4020 71470 4032
rect 71685 4029 71697 4032
rect 71731 4029 71743 4063
rect 71685 4023 71743 4029
rect 72050 4020 72056 4072
rect 72108 4060 72114 4072
rect 72329 4063 72387 4069
rect 72329 4060 72341 4063
rect 72108 4032 72341 4060
rect 72108 4020 72114 4032
rect 72329 4029 72341 4032
rect 72375 4029 72387 4063
rect 72329 4023 72387 4029
rect 72602 4020 72608 4072
rect 72660 4060 72666 4072
rect 72973 4063 73031 4069
rect 72973 4060 72985 4063
rect 72660 4032 72985 4060
rect 72660 4020 72666 4032
rect 72973 4029 72985 4032
rect 73019 4029 73031 4063
rect 72973 4023 73031 4029
rect 73246 4020 73252 4072
rect 73304 4060 73310 4072
rect 73617 4063 73675 4069
rect 73617 4060 73629 4063
rect 73304 4032 73629 4060
rect 73304 4020 73310 4032
rect 73617 4029 73629 4032
rect 73663 4029 73675 4063
rect 73617 4023 73675 4029
rect 74442 4020 74448 4072
rect 74500 4060 74506 4072
rect 74997 4063 75055 4069
rect 74997 4060 75009 4063
rect 74500 4032 75009 4060
rect 74500 4020 74506 4032
rect 74997 4029 75009 4032
rect 75043 4029 75055 4063
rect 74997 4023 75055 4029
rect 75086 4020 75092 4072
rect 75144 4060 75150 4072
rect 75641 4063 75699 4069
rect 75641 4060 75653 4063
rect 75144 4032 75653 4060
rect 75144 4020 75150 4032
rect 75641 4029 75653 4032
rect 75687 4029 75699 4063
rect 75641 4023 75699 4029
rect 75730 4020 75736 4072
rect 75788 4060 75794 4072
rect 76285 4063 76343 4069
rect 76285 4060 76297 4063
rect 75788 4032 76297 4060
rect 75788 4020 75794 4032
rect 76285 4029 76297 4032
rect 76331 4029 76343 4063
rect 77110 4060 77116 4072
rect 77071 4032 77116 4060
rect 76285 4023 76343 4029
rect 77110 4020 77116 4032
rect 77168 4020 77174 4072
rect 78306 4060 78312 4072
rect 78267 4032 78312 4060
rect 78306 4020 78312 4032
rect 78364 4020 78370 4072
rect 78950 4060 78956 4072
rect 78911 4032 78956 4060
rect 78950 4020 78956 4032
rect 79008 4020 79014 4072
rect 80790 4060 80796 4072
rect 80751 4032 80796 4060
rect 80790 4020 80796 4032
rect 80848 4020 80854 4072
rect 81342 4020 81348 4072
rect 81400 4060 81406 4072
rect 81437 4063 81495 4069
rect 81437 4060 81449 4063
rect 81400 4032 81449 4060
rect 81400 4020 81406 4032
rect 81437 4029 81449 4032
rect 81483 4029 81495 4063
rect 81437 4023 81495 4029
rect 81986 4020 81992 4072
rect 82044 4060 82050 4072
rect 82081 4063 82139 4069
rect 82081 4060 82093 4063
rect 82044 4032 82093 4060
rect 82044 4020 82050 4032
rect 82081 4029 82093 4032
rect 82127 4029 82139 4063
rect 82722 4060 82728 4072
rect 82683 4032 82728 4060
rect 82081 4023 82139 4029
rect 82722 4020 82728 4032
rect 82780 4020 82786 4072
rect 83642 4060 83648 4072
rect 83603 4032 83648 4060
rect 83642 4020 83648 4032
rect 83700 4020 83706 4072
rect 84194 4020 84200 4072
rect 84252 4060 84258 4072
rect 84289 4063 84347 4069
rect 84289 4060 84301 4063
rect 84252 4032 84301 4060
rect 84252 4020 84258 4032
rect 84289 4029 84301 4032
rect 84335 4029 84347 4063
rect 84289 4023 84347 4029
rect 84838 4020 84844 4072
rect 84896 4060 84902 4072
rect 85485 4063 85543 4069
rect 85485 4060 85497 4063
rect 84896 4032 85497 4060
rect 84896 4020 84902 4032
rect 85485 4029 85497 4032
rect 85531 4029 85543 4063
rect 85485 4023 85543 4029
rect 87598 4020 87604 4072
rect 87656 4060 87662 4072
rect 87877 4063 87935 4069
rect 87877 4060 87889 4063
rect 87656 4032 87889 4060
rect 87656 4020 87662 4032
rect 87877 4029 87889 4032
rect 87923 4029 87935 4063
rect 91186 4060 91192 4072
rect 87877 4023 87935 4029
rect 87984 4032 89714 4060
rect 91147 4032 91192 4060
rect 59872 3964 60588 3992
rect 59872 3952 59878 3964
rect 60918 3952 60924 4004
rect 60976 3992 60982 4004
rect 80882 3992 80888 4004
rect 60976 3964 80888 3992
rect 60976 3952 60982 3964
rect 80882 3952 80888 3964
rect 80940 3952 80946 4004
rect 85666 3952 85672 4004
rect 85724 3992 85730 4004
rect 87984 3992 88012 4032
rect 85724 3964 88012 3992
rect 85724 3952 85730 3964
rect 53984 3896 55168 3924
rect 53984 3884 53990 3896
rect 55674 3884 55680 3936
rect 55732 3924 55738 3936
rect 89257 3927 89315 3933
rect 89257 3924 89269 3927
rect 55732 3896 89269 3924
rect 55732 3884 55738 3896
rect 89257 3893 89269 3896
rect 89303 3893 89315 3927
rect 89686 3924 89714 4032
rect 91186 4020 91192 4032
rect 91244 4020 91250 4072
rect 91370 4060 91376 4072
rect 91331 4032 91376 4060
rect 91370 4020 91376 4032
rect 91428 4020 91434 4072
rect 91572 4069 91600 4100
rect 91833 4097 91845 4131
rect 91879 4097 91891 4131
rect 91833 4091 91891 4097
rect 92014 4088 92020 4140
rect 92072 4128 92078 4140
rect 92293 4131 92351 4137
rect 92293 4128 92305 4131
rect 92072 4100 92305 4128
rect 92072 4088 92078 4100
rect 92293 4097 92305 4100
rect 92339 4097 92351 4131
rect 92293 4091 92351 4097
rect 96985 4131 97043 4137
rect 96985 4097 96997 4131
rect 97031 4128 97043 4131
rect 97074 4128 97080 4140
rect 97031 4100 97080 4128
rect 97031 4097 97043 4100
rect 96985 4091 97043 4097
rect 97074 4088 97080 4100
rect 97132 4128 97138 4140
rect 97132 4100 97212 4128
rect 97132 4088 97138 4100
rect 91557 4063 91615 4069
rect 91557 4029 91569 4063
rect 91603 4029 91615 4063
rect 91557 4023 91615 4029
rect 91925 4063 91983 4069
rect 91925 4029 91937 4063
rect 91971 4029 91983 4063
rect 91925 4023 91983 4029
rect 91097 3995 91155 4001
rect 91097 3961 91109 3995
rect 91143 3992 91155 3995
rect 91738 3992 91744 4004
rect 91143 3964 91744 3992
rect 91143 3961 91155 3964
rect 91097 3955 91155 3961
rect 91738 3952 91744 3964
rect 91796 3952 91802 4004
rect 91940 3924 91968 4023
rect 92382 4020 92388 4072
rect 92440 4060 92446 4072
rect 93029 4063 93087 4069
rect 93029 4060 93041 4063
rect 92440 4032 93041 4060
rect 92440 4020 92446 4032
rect 93029 4029 93041 4032
rect 93075 4029 93087 4063
rect 93029 4023 93087 4029
rect 93578 4020 93584 4072
rect 93636 4060 93642 4072
rect 93673 4063 93731 4069
rect 93673 4060 93685 4063
rect 93636 4032 93685 4060
rect 93636 4020 93642 4032
rect 93673 4029 93685 4032
rect 93719 4029 93731 4063
rect 93673 4023 93731 4029
rect 94130 4020 94136 4072
rect 94188 4060 94194 4072
rect 94317 4063 94375 4069
rect 94317 4060 94329 4063
rect 94188 4032 94329 4060
rect 94188 4020 94194 4032
rect 94317 4029 94329 4032
rect 94363 4029 94375 4063
rect 94317 4023 94375 4029
rect 95418 4020 95424 4072
rect 95476 4060 95482 4072
rect 97184 4069 97212 4100
rect 95973 4063 96031 4069
rect 95973 4060 95985 4063
rect 95476 4032 95985 4060
rect 95476 4020 95482 4032
rect 95973 4029 95985 4032
rect 96019 4029 96031 4063
rect 95973 4023 96031 4029
rect 97169 4063 97227 4069
rect 97169 4029 97181 4063
rect 97215 4029 97227 4063
rect 97169 4023 97227 4029
rect 97721 4063 97779 4069
rect 97721 4029 97733 4063
rect 97767 4060 97779 4063
rect 97902 4060 97908 4072
rect 97767 4032 97908 4060
rect 97767 4029 97779 4032
rect 97721 4023 97779 4029
rect 97902 4020 97908 4032
rect 97960 4020 97966 4072
rect 97353 3995 97411 4001
rect 97353 3961 97365 3995
rect 97399 3992 97411 3995
rect 99282 3992 99288 4004
rect 97399 3964 99288 3992
rect 97399 3961 97411 3964
rect 97353 3955 97411 3961
rect 99282 3952 99288 3964
rect 99340 3952 99346 4004
rect 97994 3924 98000 3936
rect 89686 3896 91968 3924
rect 97955 3896 98000 3924
rect 89257 3887 89315 3893
rect 97994 3884 98000 3896
rect 98052 3884 98058 3936
rect 1104 3834 98808 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 50326 3834
rect 50378 3782 50390 3834
rect 50442 3782 50454 3834
rect 50506 3782 50518 3834
rect 50570 3782 81046 3834
rect 81098 3782 81110 3834
rect 81162 3782 81174 3834
rect 81226 3782 81238 3834
rect 81290 3782 98808 3834
rect 1104 3760 98808 3782
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5350 3720 5356 3732
rect 5132 3692 5356 3720
rect 5132 3680 5138 3692
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 11885 3723 11943 3729
rect 11885 3720 11897 3723
rect 11204 3692 11897 3720
rect 11204 3680 11210 3692
rect 11885 3689 11897 3692
rect 11931 3689 11943 3723
rect 19334 3720 19340 3732
rect 11885 3683 11943 3689
rect 12406 3692 14780 3720
rect 3050 3652 3056 3664
rect 3011 3624 3056 3652
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 4709 3655 4767 3661
rect 4709 3621 4721 3655
rect 4755 3652 4767 3655
rect 4798 3652 4804 3664
rect 4755 3624 4804 3652
rect 4755 3621 4767 3624
rect 4709 3615 4767 3621
rect 4798 3612 4804 3624
rect 4856 3612 4862 3664
rect 5534 3652 5540 3664
rect 5495 3624 5540 3652
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 6270 3652 6276 3664
rect 6231 3624 6276 3652
rect 6270 3612 6276 3624
rect 6328 3612 6334 3664
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 8113 3655 8171 3661
rect 8113 3652 8125 3655
rect 8076 3624 8125 3652
rect 8076 3612 8082 3624
rect 8113 3621 8125 3624
rect 8159 3621 8171 3655
rect 9950 3652 9956 3664
rect 8113 3615 8171 3621
rect 8588 3624 9956 3652
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 1946 3584 1952 3596
rect 1903 3556 1952 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2777 3587 2835 3593
rect 2777 3553 2789 3587
rect 2823 3553 2835 3587
rect 2777 3547 2835 3553
rect 106 3476 112 3528
rect 164 3516 170 3528
rect 1118 3516 1124 3528
rect 164 3488 1124 3516
rect 164 3476 170 3488
rect 1118 3476 1124 3488
rect 1176 3476 1182 3528
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3516 2191 3519
rect 2406 3516 2412 3528
rect 2179 3488 2412 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 2792 3448 2820 3547
rect 3878 3544 3884 3596
rect 3936 3584 3942 3596
rect 4341 3587 4399 3593
rect 4341 3584 4353 3587
rect 3936 3556 4353 3584
rect 3936 3544 3942 3556
rect 4341 3553 4353 3556
rect 4387 3553 4399 3587
rect 4341 3547 4399 3553
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 6917 3587 6975 3593
rect 6917 3584 6929 3587
rect 5408 3556 6929 3584
rect 5408 3544 5414 3556
rect 6917 3553 6929 3556
rect 6963 3553 6975 3587
rect 6917 3547 6975 3553
rect 7190 3544 7196 3596
rect 7248 3584 7254 3596
rect 7837 3587 7895 3593
rect 7837 3584 7849 3587
rect 7248 3556 7849 3584
rect 7248 3544 7254 3556
rect 7837 3553 7849 3556
rect 7883 3553 7895 3587
rect 8588 3584 8616 3624
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 11057 3655 11115 3661
rect 11057 3621 11069 3655
rect 11103 3652 11115 3655
rect 12406 3652 12434 3692
rect 13262 3652 13268 3664
rect 11103 3624 12434 3652
rect 13223 3624 13268 3652
rect 11103 3621 11115 3624
rect 11057 3615 11115 3621
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 7837 3547 7895 3553
rect 7944 3556 8616 3584
rect 9585 3587 9643 3593
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7944 3516 7972 3556
rect 9585 3553 9597 3587
rect 9631 3553 9643 3587
rect 10318 3584 10324 3596
rect 10279 3556 10324 3584
rect 9585 3547 9643 3553
rect 7147 3488 7972 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 8018 3476 8024 3528
rect 8076 3516 8082 3528
rect 8938 3516 8944 3528
rect 8076 3488 8944 3516
rect 8076 3476 8082 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 1360 3420 2820 3448
rect 9600 3448 9628 3547
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 11793 3587 11851 3593
rect 11793 3553 11805 3587
rect 11839 3553 11851 3587
rect 11793 3547 11851 3553
rect 12529 3587 12587 3593
rect 12529 3553 12541 3587
rect 12575 3584 12587 3587
rect 13630 3584 13636 3596
rect 12575 3556 13636 3584
rect 12575 3553 12587 3556
rect 12529 3547 12587 3553
rect 11808 3516 11836 3547
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 14752 3584 14780 3692
rect 14844 3692 19340 3720
rect 14844 3661 14872 3692
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 20680 3692 20852 3720
rect 20680 3680 20686 3692
rect 14829 3655 14887 3661
rect 14829 3621 14841 3655
rect 14875 3621 14887 3655
rect 14829 3615 14887 3621
rect 15565 3655 15623 3661
rect 15565 3621 15577 3655
rect 15611 3652 15623 3655
rect 17586 3652 17592 3664
rect 15611 3624 17592 3652
rect 15611 3621 15623 3624
rect 15565 3615 15623 3621
rect 17586 3612 17592 3624
rect 17644 3612 17650 3664
rect 17862 3612 17868 3664
rect 17920 3661 17926 3664
rect 17920 3655 17940 3661
rect 17928 3621 17940 3655
rect 17920 3615 17940 3621
rect 17920 3612 17926 3615
rect 18138 3612 18144 3664
rect 18196 3652 18202 3664
rect 20162 3652 20168 3664
rect 18196 3624 20168 3652
rect 18196 3612 18202 3624
rect 20162 3612 20168 3624
rect 20220 3612 20226 3664
rect 20824 3661 20852 3692
rect 27522 3680 27528 3732
rect 27580 3720 27586 3732
rect 29086 3720 29092 3732
rect 27580 3692 29092 3720
rect 27580 3680 27586 3692
rect 29086 3680 29092 3692
rect 29144 3680 29150 3732
rect 34698 3680 34704 3732
rect 34756 3720 34762 3732
rect 34756 3692 36676 3720
rect 34756 3680 34762 3692
rect 20809 3655 20867 3661
rect 20809 3621 20821 3655
rect 20855 3621 20867 3655
rect 21542 3652 21548 3664
rect 21503 3624 21548 3652
rect 20809 3615 20867 3621
rect 21542 3612 21548 3624
rect 21600 3612 21606 3664
rect 21818 3612 21824 3664
rect 21876 3652 21882 3664
rect 36538 3652 36544 3664
rect 21876 3624 36544 3652
rect 21876 3612 21882 3624
rect 36538 3612 36544 3624
rect 36596 3612 36602 3664
rect 16206 3584 16212 3596
rect 14752 3556 16212 3584
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 16301 3587 16359 3593
rect 16301 3553 16313 3587
rect 16347 3584 16359 3587
rect 17034 3584 17040 3596
rect 16347 3556 17040 3584
rect 16347 3553 16359 3556
rect 16301 3547 16359 3553
rect 17034 3544 17040 3556
rect 17092 3544 17098 3596
rect 17129 3587 17187 3593
rect 17129 3553 17141 3587
rect 17175 3584 17187 3587
rect 17218 3584 17224 3596
rect 17175 3556 17224 3584
rect 17175 3553 17187 3556
rect 17129 3547 17187 3553
rect 16666 3516 16672 3528
rect 11808 3488 16672 3516
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3516 16911 3519
rect 17144 3516 17172 3547
rect 17218 3544 17224 3556
rect 17276 3544 17282 3596
rect 18506 3584 18512 3596
rect 18467 3556 18512 3584
rect 18506 3544 18512 3556
rect 18564 3544 18570 3596
rect 20070 3584 20076 3596
rect 20031 3556 20076 3584
rect 20070 3544 20076 3556
rect 20128 3544 20134 3596
rect 20993 3587 21051 3593
rect 20993 3553 21005 3587
rect 21039 3584 21051 3587
rect 21174 3584 21180 3596
rect 21039 3556 21180 3584
rect 21039 3553 21051 3556
rect 20993 3547 21051 3553
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 21910 3544 21916 3596
rect 21968 3584 21974 3596
rect 22189 3587 22247 3593
rect 22189 3584 22201 3587
rect 21968 3556 22201 3584
rect 21968 3544 21974 3556
rect 22189 3553 22201 3556
rect 22235 3553 22247 3587
rect 22830 3584 22836 3596
rect 22791 3556 22836 3584
rect 22189 3547 22247 3553
rect 22830 3544 22836 3556
rect 22888 3544 22894 3596
rect 24026 3584 24032 3596
rect 23987 3556 24032 3584
rect 24026 3544 24032 3556
rect 24084 3544 24090 3596
rect 24670 3544 24676 3596
rect 24728 3584 24734 3596
rect 25225 3587 25283 3593
rect 25225 3584 25237 3587
rect 24728 3556 25237 3584
rect 24728 3544 24734 3556
rect 25225 3553 25237 3556
rect 25271 3553 25283 3587
rect 25225 3547 25283 3553
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 25869 3587 25927 3593
rect 25869 3584 25881 3587
rect 25372 3556 25881 3584
rect 25372 3544 25378 3556
rect 25869 3553 25881 3556
rect 25915 3553 25927 3587
rect 26786 3584 26792 3596
rect 26747 3556 26792 3584
rect 25869 3547 25927 3553
rect 26786 3544 26792 3556
rect 26844 3544 26850 3596
rect 27706 3584 27712 3596
rect 27667 3556 27712 3584
rect 27706 3544 27712 3556
rect 27764 3544 27770 3596
rect 28902 3584 28908 3596
rect 28863 3556 28908 3584
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 29914 3544 29920 3596
rect 29972 3584 29978 3596
rect 30469 3587 30527 3593
rect 30469 3584 30481 3587
rect 29972 3556 30481 3584
rect 29972 3544 29978 3556
rect 30469 3553 30481 3556
rect 30515 3553 30527 3587
rect 30469 3547 30527 3553
rect 30558 3544 30564 3596
rect 30616 3584 30622 3596
rect 31113 3587 31171 3593
rect 31113 3584 31125 3587
rect 30616 3556 31125 3584
rect 30616 3544 30622 3556
rect 31113 3553 31125 3556
rect 31159 3553 31171 3587
rect 31938 3584 31944 3596
rect 31899 3556 31944 3584
rect 31113 3547 31171 3553
rect 31938 3544 31944 3556
rect 31996 3544 32002 3596
rect 32585 3587 32643 3593
rect 32585 3553 32597 3587
rect 32631 3553 32643 3587
rect 32585 3547 32643 3553
rect 16899 3488 17172 3516
rect 16899 3485 16911 3488
rect 16853 3479 16911 3485
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 20622 3516 20628 3528
rect 17920 3488 20628 3516
rect 17920 3476 17926 3488
rect 13262 3448 13268 3460
rect 9600 3420 13268 3448
rect 1360 3408 1366 3420
rect 13262 3408 13268 3420
rect 13320 3408 13326 3460
rect 13446 3408 13452 3460
rect 13504 3448 13510 3460
rect 14458 3448 14464 3460
rect 13504 3420 14464 3448
rect 13504 3408 13510 3420
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 14734 3408 14740 3460
rect 14792 3448 14798 3460
rect 15749 3451 15807 3457
rect 15749 3448 15761 3451
rect 14792 3420 15761 3448
rect 14792 3408 14798 3420
rect 15749 3417 15761 3420
rect 15795 3417 15807 3451
rect 15749 3411 15807 3417
rect 16482 3408 16488 3460
rect 16540 3448 16546 3460
rect 16945 3451 17003 3457
rect 16945 3448 16957 3451
rect 16540 3420 16957 3448
rect 16540 3408 16546 3420
rect 16945 3417 16957 3420
rect 16991 3417 17003 3451
rect 16945 3411 17003 3417
rect 17126 3408 17132 3460
rect 17184 3448 17190 3460
rect 17681 3451 17739 3457
rect 17681 3448 17693 3451
rect 17184 3420 17693 3448
rect 17184 3408 17190 3420
rect 17681 3417 17693 3420
rect 17727 3417 17739 3451
rect 17681 3411 17739 3417
rect 9214 3340 9220 3392
rect 9272 3380 9278 3392
rect 9677 3383 9735 3389
rect 9677 3380 9689 3383
rect 9272 3352 9689 3380
rect 9272 3340 9278 3352
rect 9677 3349 9689 3352
rect 9723 3349 9735 3383
rect 9677 3343 9735 3349
rect 9858 3340 9864 3392
rect 9916 3380 9922 3392
rect 10413 3383 10471 3389
rect 10413 3380 10425 3383
rect 9916 3352 10425 3380
rect 9916 3340 9922 3352
rect 10413 3349 10425 3352
rect 10459 3349 10471 3383
rect 10413 3343 10471 3349
rect 10502 3340 10508 3392
rect 10560 3380 10566 3392
rect 11149 3383 11207 3389
rect 11149 3380 11161 3383
rect 10560 3352 11161 3380
rect 10560 3340 10566 3352
rect 11149 3349 11161 3352
rect 11195 3349 11207 3383
rect 11149 3343 11207 3349
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 12621 3383 12679 3389
rect 12621 3380 12633 3383
rect 11664 3352 12633 3380
rect 11664 3340 11670 3352
rect 12621 3349 12633 3352
rect 12667 3349 12679 3383
rect 12621 3343 12679 3349
rect 12894 3340 12900 3392
rect 12952 3380 12958 3392
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 12952 3352 13369 3380
rect 12952 3340 12958 3352
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 13357 3343 13415 3349
rect 14090 3340 14096 3392
rect 14148 3380 14154 3392
rect 14921 3383 14979 3389
rect 14921 3380 14933 3383
rect 14148 3352 14933 3380
rect 14148 3340 14154 3352
rect 14921 3349 14933 3352
rect 14967 3349 14979 3383
rect 14921 3343 14979 3349
rect 16022 3340 16028 3392
rect 16080 3380 16086 3392
rect 16393 3383 16451 3389
rect 16393 3380 16405 3383
rect 16080 3352 16405 3380
rect 16080 3340 16086 3352
rect 16393 3349 16405 3352
rect 16439 3349 16451 3383
rect 16393 3343 16451 3349
rect 17589 3383 17647 3389
rect 17589 3349 17601 3383
rect 17635 3380 17647 3383
rect 17972 3380 18000 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 22278 3476 22284 3528
rect 22336 3516 22342 3528
rect 22336 3488 31754 3516
rect 22336 3476 22342 3488
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 18288 3420 20760 3448
rect 18288 3408 18294 3420
rect 17635 3352 18000 3380
rect 17635 3349 17647 3352
rect 17589 3343 17647 3349
rect 18138 3340 18144 3392
rect 18196 3380 18202 3392
rect 18601 3383 18659 3389
rect 18601 3380 18613 3383
rect 18196 3352 18613 3380
rect 18196 3340 18202 3352
rect 18601 3349 18613 3352
rect 18647 3349 18659 3383
rect 18601 3343 18659 3349
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 20165 3383 20223 3389
rect 20165 3380 20177 3383
rect 19484 3352 20177 3380
rect 19484 3340 19490 3352
rect 20165 3349 20177 3352
rect 20211 3349 20223 3383
rect 20732 3380 20760 3420
rect 20806 3408 20812 3460
rect 20864 3448 20870 3460
rect 21729 3451 21787 3457
rect 21729 3448 21741 3451
rect 20864 3420 21741 3448
rect 20864 3408 20870 3420
rect 21729 3417 21741 3420
rect 21775 3417 21787 3451
rect 21729 3411 21787 3417
rect 22002 3408 22008 3460
rect 22060 3448 22066 3460
rect 25590 3448 25596 3460
rect 22060 3420 25596 3448
rect 22060 3408 22066 3420
rect 25590 3408 25596 3420
rect 25648 3408 25654 3460
rect 31726 3448 31754 3488
rect 31846 3476 31852 3528
rect 31904 3516 31910 3528
rect 32600 3516 32628 3547
rect 32858 3544 32864 3596
rect 32916 3584 32922 3596
rect 33229 3587 33287 3593
rect 33229 3584 33241 3587
rect 32916 3556 33241 3584
rect 32916 3544 32922 3556
rect 33229 3553 33241 3556
rect 33275 3553 33287 3587
rect 34422 3584 34428 3596
rect 34383 3556 34428 3584
rect 33229 3547 33287 3553
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 35434 3544 35440 3596
rect 35492 3584 35498 3596
rect 35713 3587 35771 3593
rect 35713 3584 35725 3587
rect 35492 3556 35725 3584
rect 35492 3544 35498 3556
rect 35713 3553 35725 3556
rect 35759 3553 35771 3587
rect 35713 3547 35771 3553
rect 36357 3587 36415 3593
rect 36357 3553 36369 3587
rect 36403 3553 36415 3587
rect 36648 3584 36676 3692
rect 37458 3680 37464 3732
rect 37516 3680 37522 3732
rect 37826 3680 37832 3732
rect 37884 3720 37890 3732
rect 39482 3720 39488 3732
rect 37884 3692 39488 3720
rect 37884 3680 37890 3692
rect 39482 3680 39488 3692
rect 39540 3680 39546 3732
rect 40405 3723 40463 3729
rect 40405 3689 40417 3723
rect 40451 3720 40463 3723
rect 49694 3720 49700 3732
rect 40451 3692 49700 3720
rect 40451 3689 40463 3692
rect 40405 3683 40463 3689
rect 49694 3680 49700 3692
rect 49752 3680 49758 3732
rect 76374 3720 76380 3732
rect 50172 3692 76380 3720
rect 37369 3655 37427 3661
rect 37369 3621 37381 3655
rect 37415 3652 37427 3655
rect 37476 3652 37504 3680
rect 44634 3652 44640 3664
rect 37415 3624 37504 3652
rect 37568 3624 44640 3652
rect 37415 3621 37427 3624
rect 37369 3615 37427 3621
rect 37568 3584 37596 3624
rect 44634 3612 44640 3624
rect 44692 3612 44698 3664
rect 45094 3612 45100 3664
rect 45152 3652 45158 3664
rect 48682 3652 48688 3664
rect 45152 3624 48688 3652
rect 45152 3612 45158 3624
rect 48682 3612 48688 3624
rect 48740 3612 48746 3664
rect 49602 3612 49608 3664
rect 49660 3652 49666 3664
rect 50172 3652 50200 3692
rect 76374 3680 76380 3692
rect 76432 3680 76438 3732
rect 78122 3680 78128 3732
rect 78180 3720 78186 3732
rect 78674 3720 78680 3732
rect 78180 3692 78680 3720
rect 78180 3680 78186 3692
rect 78674 3680 78680 3692
rect 78732 3680 78738 3732
rect 79318 3680 79324 3732
rect 79376 3720 79382 3732
rect 81437 3723 81495 3729
rect 81437 3720 81449 3723
rect 79376 3692 81449 3720
rect 79376 3680 79382 3692
rect 81437 3689 81449 3692
rect 81483 3720 81495 3723
rect 81483 3692 81756 3720
rect 81483 3689 81495 3692
rect 81437 3683 81495 3689
rect 49660 3624 50200 3652
rect 49660 3612 49666 3624
rect 62482 3612 62488 3664
rect 62540 3652 62546 3664
rect 62540 3624 63264 3652
rect 62540 3612 62546 3624
rect 37734 3584 37740 3596
rect 36648 3556 37596 3584
rect 37695 3556 37740 3584
rect 36357 3547 36415 3553
rect 31904 3488 32628 3516
rect 31904 3476 31910 3488
rect 35618 3476 35624 3528
rect 35676 3516 35682 3528
rect 36372 3516 36400 3547
rect 37734 3544 37740 3556
rect 37792 3544 37798 3596
rect 38102 3544 38108 3596
rect 38160 3584 38166 3596
rect 38933 3587 38991 3593
rect 38933 3584 38945 3587
rect 38160 3556 38945 3584
rect 38160 3544 38166 3556
rect 38933 3553 38945 3556
rect 38979 3553 38991 3587
rect 38933 3547 38991 3553
rect 39298 3544 39304 3596
rect 39356 3584 39362 3596
rect 39577 3587 39635 3593
rect 39577 3584 39589 3587
rect 39356 3556 39589 3584
rect 39356 3544 39362 3556
rect 39577 3553 39589 3556
rect 39623 3553 39635 3587
rect 39577 3547 39635 3553
rect 40494 3544 40500 3596
rect 40552 3584 40558 3596
rect 40957 3587 41015 3593
rect 40957 3584 40969 3587
rect 40552 3556 40969 3584
rect 40552 3544 40558 3556
rect 40957 3553 40969 3556
rect 41003 3553 41015 3587
rect 41690 3584 41696 3596
rect 41651 3556 41696 3584
rect 40957 3547 41015 3553
rect 41690 3544 41696 3556
rect 41748 3544 41754 3596
rect 42334 3584 42340 3596
rect 42295 3556 42340 3584
rect 42334 3544 42340 3556
rect 42392 3544 42398 3596
rect 42978 3584 42984 3596
rect 42939 3556 42984 3584
rect 42978 3544 42984 3556
rect 43036 3544 43042 3596
rect 43625 3587 43683 3593
rect 43625 3553 43637 3587
rect 43671 3553 43683 3587
rect 44818 3584 44824 3596
rect 44779 3556 44824 3584
rect 43625 3547 43683 3553
rect 35676 3488 36400 3516
rect 35676 3476 35682 3488
rect 42242 3476 42248 3528
rect 42300 3516 42306 3528
rect 43640 3516 43668 3547
rect 44818 3544 44824 3556
rect 44876 3544 44882 3596
rect 46566 3544 46572 3596
rect 46624 3584 46630 3596
rect 47213 3587 47271 3593
rect 47213 3584 47225 3587
rect 46624 3556 47225 3584
rect 46624 3544 46630 3556
rect 47213 3553 47225 3556
rect 47259 3553 47271 3587
rect 47213 3547 47271 3553
rect 47302 3544 47308 3596
rect 47360 3584 47366 3596
rect 47857 3587 47915 3593
rect 47857 3584 47869 3587
rect 47360 3556 47869 3584
rect 47360 3544 47366 3556
rect 47857 3553 47869 3556
rect 47903 3553 47915 3587
rect 47857 3547 47915 3553
rect 47946 3544 47952 3596
rect 48004 3584 48010 3596
rect 48501 3587 48559 3593
rect 48501 3584 48513 3587
rect 48004 3556 48513 3584
rect 48004 3544 48010 3556
rect 48501 3553 48513 3556
rect 48547 3553 48559 3587
rect 48501 3547 48559 3553
rect 49145 3587 49203 3593
rect 49145 3553 49157 3587
rect 49191 3553 49203 3587
rect 49145 3547 49203 3553
rect 42300 3488 43668 3516
rect 42300 3476 42306 3488
rect 48406 3476 48412 3528
rect 48464 3516 48470 3528
rect 49160 3516 49188 3547
rect 49778 3544 49784 3596
rect 49836 3584 49842 3596
rect 49836 3556 49881 3584
rect 49836 3544 49842 3556
rect 50890 3544 50896 3596
rect 50948 3584 50954 3596
rect 51445 3587 51503 3593
rect 51445 3584 51457 3587
rect 50948 3556 51457 3584
rect 50948 3544 50954 3556
rect 51445 3553 51457 3556
rect 51491 3553 51503 3587
rect 52086 3584 52092 3596
rect 52047 3556 52092 3584
rect 51445 3547 51503 3553
rect 52086 3544 52092 3556
rect 52144 3544 52150 3596
rect 52730 3584 52736 3596
rect 52691 3556 52736 3584
rect 52730 3544 52736 3556
rect 52788 3544 52794 3596
rect 53282 3544 53288 3596
rect 53340 3584 53346 3596
rect 53377 3587 53435 3593
rect 53377 3584 53389 3587
rect 53340 3556 53389 3584
rect 53340 3544 53346 3556
rect 53377 3553 53389 3556
rect 53423 3553 53435 3587
rect 53377 3547 53435 3553
rect 53926 3544 53932 3596
rect 53984 3584 53990 3596
rect 54021 3587 54079 3593
rect 54021 3584 54033 3587
rect 53984 3556 54033 3584
rect 53984 3544 53990 3556
rect 54021 3553 54033 3556
rect 54067 3553 54079 3587
rect 54021 3547 54079 3553
rect 54570 3544 54576 3596
rect 54628 3584 54634 3596
rect 54665 3587 54723 3593
rect 54665 3584 54677 3587
rect 54628 3556 54677 3584
rect 54628 3544 54634 3556
rect 54665 3553 54677 3556
rect 54711 3553 54723 3587
rect 54665 3547 54723 3553
rect 55122 3544 55128 3596
rect 55180 3584 55186 3596
rect 55309 3587 55367 3593
rect 55309 3584 55321 3587
rect 55180 3556 55321 3584
rect 55180 3544 55186 3556
rect 55309 3553 55321 3556
rect 55355 3553 55367 3587
rect 55309 3547 55367 3553
rect 56318 3544 56324 3596
rect 56376 3584 56382 3596
rect 56689 3587 56747 3593
rect 56689 3584 56701 3587
rect 56376 3556 56701 3584
rect 56376 3544 56382 3556
rect 56689 3553 56701 3556
rect 56735 3553 56747 3587
rect 56689 3547 56747 3553
rect 57146 3544 57152 3596
rect 57204 3584 57210 3596
rect 57333 3587 57391 3593
rect 57333 3584 57345 3587
rect 57204 3556 57345 3584
rect 57204 3544 57210 3556
rect 57333 3553 57345 3556
rect 57379 3553 57391 3587
rect 58158 3584 58164 3596
rect 58119 3556 58164 3584
rect 57333 3547 57391 3553
rect 58158 3544 58164 3556
rect 58216 3544 58222 3596
rect 58802 3584 58808 3596
rect 58763 3556 58808 3584
rect 58802 3544 58808 3556
rect 58860 3544 58866 3596
rect 59449 3587 59507 3593
rect 59449 3553 59461 3587
rect 59495 3553 59507 3587
rect 60642 3584 60648 3596
rect 60603 3556 60648 3584
rect 59449 3547 59507 3553
rect 48464 3488 49188 3516
rect 48464 3476 48470 3488
rect 57974 3476 57980 3528
rect 58032 3516 58038 3528
rect 59464 3516 59492 3547
rect 60642 3544 60648 3556
rect 60700 3544 60706 3596
rect 61286 3544 61292 3596
rect 61344 3584 61350 3596
rect 63236 3593 63264 3624
rect 64046 3612 64052 3664
rect 64104 3652 64110 3664
rect 64104 3624 65840 3652
rect 64104 3612 64110 3624
rect 61933 3587 61991 3593
rect 61933 3584 61945 3587
rect 61344 3556 61945 3584
rect 61344 3544 61350 3556
rect 61933 3553 61945 3556
rect 61979 3553 61991 3587
rect 61933 3547 61991 3553
rect 62577 3587 62635 3593
rect 62577 3553 62589 3587
rect 62623 3553 62635 3587
rect 62577 3547 62635 3553
rect 63221 3587 63279 3593
rect 63221 3553 63233 3587
rect 63267 3553 63279 3587
rect 63865 3587 63923 3593
rect 63865 3584 63877 3587
rect 63221 3547 63279 3553
rect 63328 3556 63877 3584
rect 58032 3488 59492 3516
rect 58032 3476 58038 3488
rect 61838 3476 61844 3528
rect 61896 3516 61902 3528
rect 62592 3516 62620 3547
rect 61896 3488 62620 3516
rect 61896 3476 61902 3488
rect 63034 3476 63040 3528
rect 63092 3516 63098 3528
rect 63328 3516 63356 3556
rect 63865 3553 63877 3556
rect 63911 3553 63923 3587
rect 63865 3547 63923 3553
rect 64509 3587 64567 3593
rect 64509 3553 64521 3587
rect 64555 3553 64567 3587
rect 64509 3547 64567 3553
rect 63092 3488 63356 3516
rect 63092 3476 63098 3488
rect 63678 3476 63684 3528
rect 63736 3516 63742 3528
rect 64524 3516 64552 3547
rect 64874 3544 64880 3596
rect 64932 3584 64938 3596
rect 65812 3593 65840 3624
rect 71314 3612 71320 3664
rect 71372 3652 71378 3664
rect 78582 3652 78588 3664
rect 71372 3624 78588 3652
rect 71372 3612 71378 3624
rect 78582 3612 78588 3624
rect 78640 3612 78646 3664
rect 80238 3652 80244 3664
rect 78692 3624 80244 3652
rect 65153 3587 65211 3593
rect 65153 3584 65165 3587
rect 64932 3556 65165 3584
rect 64932 3544 64938 3556
rect 65153 3553 65165 3556
rect 65199 3553 65211 3587
rect 65153 3547 65211 3553
rect 65797 3587 65855 3593
rect 65797 3553 65809 3587
rect 65843 3553 65855 3587
rect 65797 3547 65855 3553
rect 66714 3544 66720 3596
rect 66772 3584 66778 3596
rect 67177 3587 67235 3593
rect 67177 3584 67189 3587
rect 66772 3556 67189 3584
rect 66772 3544 66778 3556
rect 67177 3553 67189 3556
rect 67223 3553 67235 3587
rect 67910 3584 67916 3596
rect 67871 3556 67916 3584
rect 67177 3547 67235 3553
rect 67910 3544 67916 3556
rect 67968 3544 67974 3596
rect 68554 3584 68560 3596
rect 68515 3556 68560 3584
rect 68554 3544 68560 3556
rect 68612 3544 68618 3596
rect 69198 3584 69204 3596
rect 69159 3556 69204 3584
rect 69198 3544 69204 3556
rect 69256 3544 69262 3596
rect 69750 3544 69756 3596
rect 69808 3584 69814 3596
rect 69845 3587 69903 3593
rect 69845 3584 69857 3587
rect 69808 3556 69857 3584
rect 69808 3544 69814 3556
rect 69845 3553 69857 3556
rect 69891 3553 69903 3587
rect 69845 3547 69903 3553
rect 70394 3544 70400 3596
rect 70452 3584 70458 3596
rect 70489 3587 70547 3593
rect 70489 3584 70501 3587
rect 70452 3556 70501 3584
rect 70452 3544 70458 3556
rect 70489 3553 70501 3556
rect 70535 3553 70547 3587
rect 70489 3547 70547 3553
rect 71038 3544 71044 3596
rect 71096 3584 71102 3596
rect 71133 3587 71191 3593
rect 71133 3584 71145 3587
rect 71096 3556 71145 3584
rect 71096 3544 71102 3556
rect 71133 3553 71145 3556
rect 71179 3553 71191 3587
rect 71133 3547 71191 3553
rect 71590 3544 71596 3596
rect 71648 3584 71654 3596
rect 72421 3587 72479 3593
rect 72421 3584 72433 3587
rect 71648 3556 72433 3584
rect 71648 3544 71654 3556
rect 72421 3553 72433 3556
rect 72467 3553 72479 3587
rect 72421 3547 72479 3553
rect 72786 3544 72792 3596
rect 72844 3584 72850 3596
rect 73065 3587 73123 3593
rect 73065 3584 73077 3587
rect 72844 3556 73077 3584
rect 72844 3544 72850 3556
rect 73065 3553 73077 3556
rect 73111 3553 73123 3587
rect 74074 3584 74080 3596
rect 74035 3556 74080 3584
rect 73065 3547 73123 3553
rect 74074 3544 74080 3556
rect 74132 3544 74138 3596
rect 74626 3544 74632 3596
rect 74684 3584 74690 3596
rect 74721 3587 74779 3593
rect 74721 3584 74733 3587
rect 74684 3556 74733 3584
rect 74684 3544 74690 3556
rect 74721 3553 74733 3556
rect 74767 3553 74779 3587
rect 75914 3584 75920 3596
rect 75875 3556 75920 3584
rect 74721 3547 74779 3553
rect 75914 3544 75920 3556
rect 75972 3544 75978 3596
rect 76466 3544 76472 3596
rect 76524 3584 76530 3596
rect 76561 3587 76619 3593
rect 76561 3584 76573 3587
rect 76524 3556 76573 3584
rect 76524 3544 76530 3556
rect 76561 3553 76573 3556
rect 76607 3553 76619 3587
rect 76561 3547 76619 3553
rect 77662 3544 77668 3596
rect 77720 3584 77726 3596
rect 78309 3587 78367 3593
rect 78309 3584 78321 3587
rect 77720 3556 78321 3584
rect 77720 3544 77726 3556
rect 78309 3553 78321 3556
rect 78355 3553 78367 3587
rect 78309 3547 78367 3553
rect 63736 3488 64552 3516
rect 63736 3476 63742 3488
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 74902 3516 74908 3528
rect 65576 3488 74908 3516
rect 65576 3476 65582 3488
rect 74902 3476 74908 3488
rect 74960 3476 74966 3528
rect 78692 3516 78720 3624
rect 80238 3612 80244 3624
rect 80296 3612 80302 3664
rect 81728 3661 81756 3692
rect 82354 3680 82360 3732
rect 82412 3720 82418 3732
rect 83550 3720 83556 3732
rect 82412 3692 83556 3720
rect 82412 3680 82418 3692
rect 83550 3680 83556 3692
rect 83608 3680 83614 3732
rect 87874 3680 87880 3732
rect 87932 3720 87938 3732
rect 88794 3720 88800 3732
rect 87932 3692 88800 3720
rect 87932 3680 87938 3692
rect 88794 3680 88800 3692
rect 88852 3680 88858 3732
rect 89346 3680 89352 3732
rect 89404 3720 89410 3732
rect 89404 3692 93854 3720
rect 89404 3680 89410 3692
rect 81713 3655 81771 3661
rect 81713 3621 81725 3655
rect 81759 3621 81771 3655
rect 81713 3615 81771 3621
rect 88702 3612 88708 3664
rect 88760 3652 88766 3664
rect 88760 3624 89484 3652
rect 88760 3612 88766 3624
rect 79321 3587 79379 3593
rect 79321 3584 79333 3587
rect 75196 3488 78720 3516
rect 78968 3556 79333 3584
rect 40405 3451 40463 3457
rect 40405 3448 40417 3451
rect 31726 3420 40417 3448
rect 40405 3417 40417 3420
rect 40451 3417 40463 3451
rect 40405 3411 40463 3417
rect 43070 3408 43076 3460
rect 43128 3448 43134 3460
rect 43128 3420 55720 3448
rect 43128 3408 43134 3420
rect 21818 3380 21824 3392
rect 20732 3352 21824 3380
rect 20165 3343 20223 3349
rect 21818 3340 21824 3352
rect 21876 3340 21882 3392
rect 23934 3340 23940 3392
rect 23992 3380 23998 3392
rect 26234 3380 26240 3392
rect 23992 3352 26240 3380
rect 23992 3340 23998 3352
rect 26234 3340 26240 3352
rect 26292 3340 26298 3392
rect 26694 3340 26700 3392
rect 26752 3380 26758 3392
rect 26881 3383 26939 3389
rect 26881 3380 26893 3383
rect 26752 3352 26893 3380
rect 26752 3340 26758 3352
rect 26881 3349 26893 3352
rect 26927 3349 26939 3383
rect 26881 3343 26939 3349
rect 32398 3340 32404 3392
rect 32456 3380 32462 3392
rect 32858 3380 32864 3392
rect 32456 3352 32864 3380
rect 32456 3340 32462 3352
rect 32858 3340 32864 3352
rect 32916 3340 32922 3392
rect 35802 3340 35808 3392
rect 35860 3380 35866 3392
rect 38930 3380 38936 3392
rect 35860 3352 38936 3380
rect 35860 3340 35866 3352
rect 38930 3340 38936 3352
rect 38988 3340 38994 3392
rect 46753 3383 46811 3389
rect 46753 3349 46765 3383
rect 46799 3380 46811 3383
rect 54018 3380 54024 3392
rect 46799 3352 54024 3380
rect 46799 3349 46811 3352
rect 46753 3343 46811 3349
rect 54018 3340 54024 3352
rect 54076 3340 54082 3392
rect 55692 3380 55720 3420
rect 55766 3408 55772 3460
rect 55824 3448 55830 3460
rect 75196 3448 75224 3488
rect 78968 3457 78996 3556
rect 79321 3553 79333 3556
rect 79367 3553 79379 3587
rect 79321 3547 79379 3553
rect 79594 3544 79600 3596
rect 79652 3584 79658 3596
rect 79873 3587 79931 3593
rect 79873 3584 79885 3587
rect 79652 3556 79885 3584
rect 79652 3544 79658 3556
rect 79873 3553 79885 3556
rect 79919 3553 79931 3587
rect 79873 3547 79931 3553
rect 80146 3544 80152 3596
rect 80204 3584 80210 3596
rect 80517 3587 80575 3593
rect 80517 3584 80529 3587
rect 80204 3556 80529 3584
rect 80204 3544 80210 3556
rect 80517 3553 80529 3556
rect 80563 3553 80575 3587
rect 82998 3584 83004 3596
rect 82959 3556 83004 3584
rect 80517 3547 80575 3553
rect 82998 3544 83004 3556
rect 83056 3544 83062 3596
rect 83826 3544 83832 3596
rect 83884 3584 83890 3596
rect 84289 3587 84347 3593
rect 84289 3584 84301 3587
rect 83884 3556 84301 3584
rect 83884 3544 83890 3556
rect 84289 3553 84301 3556
rect 84335 3553 84347 3587
rect 84289 3547 84347 3553
rect 84378 3544 84384 3596
rect 84436 3584 84442 3596
rect 84933 3587 84991 3593
rect 84933 3584 84945 3587
rect 84436 3556 84945 3584
rect 84436 3544 84442 3556
rect 84933 3553 84945 3556
rect 84979 3553 84991 3587
rect 84933 3547 84991 3553
rect 85022 3544 85028 3596
rect 85080 3584 85086 3596
rect 85577 3587 85635 3593
rect 85577 3584 85589 3587
rect 85080 3556 85589 3584
rect 85080 3544 85086 3556
rect 85577 3553 85589 3556
rect 85623 3553 85635 3587
rect 86218 3584 86224 3596
rect 86179 3556 86224 3584
rect 85577 3547 85635 3553
rect 86218 3544 86224 3556
rect 86276 3544 86282 3596
rect 86862 3584 86868 3596
rect 86823 3556 86868 3584
rect 86862 3544 86868 3556
rect 86920 3544 86926 3596
rect 87506 3544 87512 3596
rect 87564 3584 87570 3596
rect 89456 3593 89484 3624
rect 89898 3612 89904 3664
rect 89956 3652 89962 3664
rect 89956 3624 90772 3652
rect 89956 3612 89962 3624
rect 90744 3593 90772 3624
rect 91738 3612 91744 3664
rect 91796 3652 91802 3664
rect 93826 3652 93854 3692
rect 96617 3655 96675 3661
rect 91796 3624 93440 3652
rect 93826 3624 95832 3652
rect 91796 3612 91802 3624
rect 93412 3593 93440 3624
rect 88153 3587 88211 3593
rect 88153 3584 88165 3587
rect 87564 3556 88165 3584
rect 87564 3544 87570 3556
rect 88153 3553 88165 3556
rect 88199 3553 88211 3587
rect 88153 3547 88211 3553
rect 88797 3587 88855 3593
rect 88797 3553 88809 3587
rect 88843 3553 88855 3587
rect 88797 3547 88855 3553
rect 89441 3587 89499 3593
rect 89441 3553 89453 3587
rect 89487 3553 89499 3587
rect 89441 3547 89499 3553
rect 90085 3587 90143 3593
rect 90085 3553 90097 3587
rect 90131 3553 90143 3587
rect 90085 3547 90143 3553
rect 90729 3587 90787 3593
rect 90729 3553 90741 3587
rect 90775 3553 90787 3587
rect 91373 3587 91431 3593
rect 91373 3584 91385 3587
rect 90729 3547 90787 3553
rect 90836 3556 91385 3584
rect 88058 3476 88064 3528
rect 88116 3516 88122 3528
rect 88812 3516 88840 3547
rect 88116 3488 88840 3516
rect 88116 3476 88122 3488
rect 78953 3451 79011 3457
rect 78953 3448 78965 3451
rect 55824 3420 75224 3448
rect 76208 3420 78965 3448
rect 55824 3408 55830 3420
rect 56870 3380 56876 3392
rect 55692 3352 56876 3380
rect 56870 3340 56876 3352
rect 56928 3340 56934 3392
rect 61654 3340 61660 3392
rect 61712 3380 61718 3392
rect 62022 3380 62028 3392
rect 61712 3352 62028 3380
rect 61712 3340 61718 3352
rect 62022 3340 62028 3352
rect 62080 3340 62086 3392
rect 62850 3340 62856 3392
rect 62908 3380 62914 3392
rect 63218 3380 63224 3392
rect 62908 3352 63224 3380
rect 62908 3340 62914 3352
rect 63218 3340 63224 3352
rect 63276 3340 63282 3392
rect 74534 3340 74540 3392
rect 74592 3380 74598 3392
rect 76208 3380 76236 3420
rect 78953 3417 78965 3420
rect 78999 3417 79011 3451
rect 79134 3448 79140 3460
rect 79095 3420 79140 3448
rect 78953 3411 79011 3417
rect 79134 3408 79140 3420
rect 79192 3408 79198 3460
rect 81526 3448 81532 3460
rect 81487 3420 81532 3448
rect 81526 3408 81532 3420
rect 81584 3408 81590 3460
rect 83734 3408 83740 3460
rect 83792 3448 83798 3460
rect 83829 3451 83887 3457
rect 83829 3448 83841 3451
rect 83792 3420 83841 3448
rect 83792 3408 83798 3420
rect 83829 3417 83841 3420
rect 83875 3417 83887 3451
rect 83829 3411 83887 3417
rect 89254 3408 89260 3460
rect 89312 3448 89318 3460
rect 90100 3448 90128 3547
rect 90542 3476 90548 3528
rect 90600 3516 90606 3528
rect 90836 3516 90864 3556
rect 91373 3553 91385 3556
rect 91419 3553 91431 3587
rect 91373 3547 91431 3553
rect 92017 3587 92075 3593
rect 92017 3553 92029 3587
rect 92063 3553 92075 3587
rect 92017 3547 92075 3553
rect 93397 3587 93455 3593
rect 93397 3553 93409 3587
rect 93443 3553 93455 3587
rect 94041 3587 94099 3593
rect 94041 3584 94053 3587
rect 93397 3547 93455 3553
rect 93826 3556 94053 3584
rect 90600 3488 90864 3516
rect 90600 3476 90606 3488
rect 91094 3476 91100 3528
rect 91152 3516 91158 3528
rect 92032 3516 92060 3547
rect 91152 3488 92060 3516
rect 91152 3476 91158 3488
rect 93026 3476 93032 3528
rect 93084 3516 93090 3528
rect 93826 3516 93854 3556
rect 94041 3553 94053 3556
rect 94087 3553 94099 3587
rect 94041 3547 94099 3553
rect 94869 3587 94927 3593
rect 94869 3553 94881 3587
rect 94915 3584 94927 3587
rect 95050 3584 95056 3596
rect 94915 3556 95056 3584
rect 94915 3553 94927 3556
rect 94869 3547 94927 3553
rect 95050 3544 95056 3556
rect 95108 3584 95114 3596
rect 95145 3587 95203 3593
rect 95145 3584 95157 3587
rect 95108 3556 95157 3584
rect 95108 3544 95114 3556
rect 95145 3553 95157 3556
rect 95191 3553 95203 3587
rect 95145 3547 95203 3553
rect 95697 3587 95755 3593
rect 95697 3553 95709 3587
rect 95743 3553 95755 3587
rect 95804 3584 95832 3624
rect 96617 3621 96629 3655
rect 96663 3652 96675 3655
rect 96798 3652 96804 3664
rect 96663 3624 96804 3652
rect 96663 3621 96675 3624
rect 96617 3615 96675 3621
rect 96798 3612 96804 3624
rect 96856 3612 96862 3664
rect 97537 3587 97595 3593
rect 97537 3584 97549 3587
rect 95804 3556 97549 3584
rect 95697 3547 95755 3553
rect 97537 3553 97549 3556
rect 97583 3553 97595 3587
rect 97537 3547 97595 3553
rect 93084 3488 93854 3516
rect 93084 3476 93090 3488
rect 94774 3476 94780 3528
rect 94832 3516 94838 3528
rect 95712 3516 95740 3547
rect 94832 3488 95740 3516
rect 94832 3476 94838 3488
rect 96154 3476 96160 3528
rect 96212 3516 96218 3528
rect 99466 3516 99472 3528
rect 96212 3488 99472 3516
rect 96212 3476 96218 3488
rect 99466 3476 99472 3488
rect 99524 3476 99530 3528
rect 94958 3448 94964 3460
rect 89312 3420 90128 3448
rect 94919 3420 94964 3448
rect 89312 3408 89318 3420
rect 94958 3408 94964 3420
rect 95016 3408 95022 3460
rect 96985 3451 97043 3457
rect 96985 3417 96997 3451
rect 97031 3448 97043 3451
rect 98638 3448 98644 3460
rect 97031 3420 98644 3448
rect 97031 3417 97043 3420
rect 96985 3411 97043 3417
rect 98638 3408 98644 3420
rect 98696 3408 98702 3460
rect 74592 3352 76236 3380
rect 77849 3383 77907 3389
rect 74592 3340 74598 3352
rect 77849 3349 77861 3383
rect 77895 3380 77907 3383
rect 78030 3380 78036 3392
rect 77895 3352 78036 3380
rect 77895 3349 77907 3352
rect 77849 3343 77907 3349
rect 78030 3340 78036 3352
rect 78088 3340 78094 3392
rect 97442 3340 97448 3392
rect 97500 3380 97506 3392
rect 97629 3383 97687 3389
rect 97629 3380 97641 3383
rect 97500 3352 97641 3380
rect 97500 3340 97506 3352
rect 97629 3349 97641 3352
rect 97675 3349 97687 3383
rect 97629 3343 97687 3349
rect 1104 3290 98808 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 65686 3290
rect 65738 3238 65750 3290
rect 65802 3238 65814 3290
rect 65866 3238 65878 3290
rect 65930 3238 96406 3290
rect 96458 3238 96470 3290
rect 96522 3238 96534 3290
rect 96586 3238 96598 3290
rect 96650 3238 98808 3290
rect 1104 3216 98808 3238
rect 4249 3179 4307 3185
rect 4249 3145 4261 3179
rect 4295 3176 4307 3179
rect 5166 3176 5172 3188
rect 4295 3148 5172 3176
rect 4295 3145 4307 3148
rect 4249 3139 4307 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 9674 3176 9680 3188
rect 5500 3148 9680 3176
rect 5500 3136 5506 3148
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 14366 3176 14372 3188
rect 13320 3148 13952 3176
rect 14327 3148 14372 3176
rect 13320 3136 13326 3148
rect 5074 3108 5080 3120
rect 5035 3080 5080 3108
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 8202 3108 8208 3120
rect 6886 3080 8208 3108
rect 2130 3040 2136 3052
rect 2091 3012 2136 3040
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 3786 3040 3792 3052
rect 3375 3012 3792 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4890 3040 4896 3052
rect 4212 3012 4896 3040
rect 4212 3000 4218 3012
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 6886 3040 6914 3080
rect 8202 3068 8208 3080
rect 8260 3068 8266 3120
rect 10318 3068 10324 3120
rect 10376 3108 10382 3120
rect 10376 3080 13860 3108
rect 10376 3068 10382 3080
rect 5736 3012 6914 3040
rect 7193 3043 7251 3049
rect 1486 2932 1492 2984
rect 1544 2972 1550 2984
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 1544 2944 1593 2972
rect 1544 2932 1550 2944
rect 1581 2941 1593 2944
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 2314 2932 2320 2984
rect 2372 2972 2378 2984
rect 2777 2975 2835 2981
rect 2777 2972 2789 2975
rect 2372 2944 2789 2972
rect 2372 2932 2378 2944
rect 2777 2941 2789 2944
rect 2823 2941 2835 2975
rect 2777 2935 2835 2941
rect 2866 2932 2872 2984
rect 2924 2972 2930 2984
rect 5736 2981 5764 3012
rect 7193 3009 7205 3043
rect 7239 3040 7251 3043
rect 7466 3040 7472 3052
rect 7239 3012 7472 3040
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 7558 3000 7564 3052
rect 7616 3040 7622 3052
rect 9122 3040 9128 3052
rect 7616 3012 9128 3040
rect 7616 3000 7622 3012
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3040 10931 3043
rect 11790 3040 11796 3052
rect 10919 3012 11796 3040
rect 10919 3009 10931 3012
rect 10873 3003 10931 3009
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 13538 3040 13544 3052
rect 13499 3012 13544 3040
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 2924 2944 3985 2972
rect 2924 2932 2930 2944
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2941 5779 2975
rect 5721 2935 5779 2941
rect 5994 2932 6000 2984
rect 6052 2972 6058 2984
rect 7745 2975 7803 2981
rect 7745 2972 7757 2975
rect 6052 2944 7757 2972
rect 6052 2932 6058 2944
rect 7745 2941 7757 2944
rect 7791 2941 7803 2975
rect 7745 2935 7803 2941
rect 7926 2932 7932 2984
rect 7984 2972 7990 2984
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7984 2944 8033 2972
rect 7984 2932 7990 2944
rect 8021 2941 8033 2944
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 10284 2944 10333 2972
rect 10284 2932 10290 2944
rect 10321 2941 10333 2944
rect 10367 2941 10379 2975
rect 12066 2972 12072 2984
rect 12027 2944 12072 2972
rect 10321 2935 10379 2941
rect 12066 2932 12072 2944
rect 12124 2932 12130 2984
rect 13262 2972 13268 2984
rect 13223 2944 13268 2972
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 4614 2864 4620 2916
rect 4672 2904 4678 2916
rect 4893 2907 4951 2913
rect 4893 2904 4905 2907
rect 4672 2876 4905 2904
rect 4672 2864 4678 2876
rect 4893 2873 4905 2876
rect 4939 2873 4951 2907
rect 4893 2867 4951 2873
rect 6362 2864 6368 2916
rect 6420 2904 6426 2916
rect 6917 2907 6975 2913
rect 6917 2904 6929 2907
rect 6420 2876 6929 2904
rect 6420 2864 6426 2876
rect 6917 2873 6929 2876
rect 6963 2873 6975 2907
rect 6917 2867 6975 2873
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 9125 2907 9183 2913
rect 9125 2904 9137 2907
rect 9088 2876 9137 2904
rect 9088 2864 9094 2876
rect 9125 2873 9137 2876
rect 9171 2873 9183 2907
rect 12342 2904 12348 2916
rect 12303 2876 12348 2904
rect 9125 2867 9183 2873
rect 12342 2864 12348 2876
rect 12400 2864 12406 2916
rect 13832 2904 13860 3080
rect 13924 3040 13952 3148
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 14458 3136 14464 3188
rect 14516 3176 14522 3188
rect 15930 3176 15936 3188
rect 14516 3148 15148 3176
rect 15891 3148 15936 3176
rect 14516 3136 14522 3148
rect 14182 3068 14188 3120
rect 14240 3108 14246 3120
rect 15010 3108 15016 3120
rect 14240 3080 15016 3108
rect 14240 3068 14246 3080
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 15120 3108 15148 3148
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 16666 3136 16672 3188
rect 16724 3176 16730 3188
rect 20162 3176 20168 3188
rect 16724 3148 20168 3176
rect 16724 3136 16730 3148
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 20257 3179 20315 3185
rect 20257 3145 20269 3179
rect 20303 3176 20315 3179
rect 20438 3176 20444 3188
rect 20303 3148 20444 3176
rect 20303 3145 20315 3148
rect 20257 3139 20315 3145
rect 20438 3136 20444 3148
rect 20496 3136 20502 3188
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 20993 3179 21051 3185
rect 20993 3176 21005 3179
rect 20956 3148 21005 3176
rect 20956 3136 20962 3148
rect 20993 3145 21005 3148
rect 21039 3145 21051 3179
rect 20993 3139 21051 3145
rect 21634 3136 21640 3188
rect 21692 3176 21698 3188
rect 21818 3176 21824 3188
rect 21692 3148 21824 3176
rect 21692 3136 21698 3148
rect 21818 3136 21824 3148
rect 21876 3136 21882 3188
rect 35802 3176 35808 3188
rect 21928 3148 35808 3176
rect 19058 3108 19064 3120
rect 15120 3080 19064 3108
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 19150 3068 19156 3120
rect 19208 3108 19214 3120
rect 21928 3108 21956 3148
rect 35802 3136 35808 3148
rect 35860 3136 35866 3188
rect 38010 3136 38016 3188
rect 38068 3176 38074 3188
rect 38105 3179 38163 3185
rect 38105 3176 38117 3179
rect 38068 3148 38117 3176
rect 38068 3136 38074 3148
rect 38105 3145 38117 3148
rect 38151 3145 38163 3179
rect 38105 3139 38163 3145
rect 38194 3136 38200 3188
rect 38252 3176 38258 3188
rect 39482 3176 39488 3188
rect 38252 3148 39488 3176
rect 38252 3136 38258 3148
rect 39482 3136 39488 3148
rect 39540 3136 39546 3188
rect 39574 3136 39580 3188
rect 39632 3176 39638 3188
rect 74534 3176 74540 3188
rect 39632 3148 74540 3176
rect 39632 3136 39638 3148
rect 74534 3136 74540 3148
rect 74592 3136 74598 3188
rect 74810 3176 74816 3188
rect 74771 3148 74816 3176
rect 74810 3136 74816 3148
rect 74868 3136 74874 3188
rect 76374 3176 76380 3188
rect 76287 3148 76380 3176
rect 76374 3136 76380 3148
rect 76432 3176 76438 3188
rect 76469 3179 76527 3185
rect 76469 3176 76481 3179
rect 76432 3148 76481 3176
rect 76432 3136 76438 3148
rect 76469 3145 76481 3148
rect 76515 3145 76527 3179
rect 78490 3176 78496 3188
rect 78451 3148 78496 3176
rect 76469 3139 76527 3145
rect 78490 3136 78496 3148
rect 78548 3136 78554 3188
rect 78582 3136 78588 3188
rect 78640 3176 78646 3188
rect 80701 3179 80759 3185
rect 80701 3176 80713 3179
rect 78640 3148 80713 3176
rect 78640 3136 78646 3148
rect 80701 3145 80713 3148
rect 80747 3176 80759 3179
rect 80793 3179 80851 3185
rect 80793 3176 80805 3179
rect 80747 3148 80805 3176
rect 80747 3145 80759 3148
rect 80701 3139 80759 3145
rect 80793 3145 80805 3148
rect 80839 3145 80851 3179
rect 80793 3139 80851 3145
rect 80882 3136 80888 3188
rect 80940 3176 80946 3188
rect 81529 3179 81587 3185
rect 81529 3176 81541 3179
rect 80940 3148 81541 3176
rect 80940 3136 80946 3148
rect 81529 3145 81541 3148
rect 81575 3145 81587 3179
rect 81529 3139 81587 3145
rect 19208 3080 21956 3108
rect 22005 3111 22063 3117
rect 19208 3068 19214 3080
rect 22005 3077 22017 3111
rect 22051 3108 22063 3111
rect 65518 3108 65524 3120
rect 22051 3080 65524 3108
rect 22051 3077 22063 3080
rect 22005 3071 22063 3077
rect 65518 3068 65524 3080
rect 65576 3068 65582 3120
rect 66806 3108 66812 3120
rect 66767 3080 66812 3108
rect 66806 3068 66812 3080
rect 66864 3068 66870 3120
rect 69290 3068 69296 3120
rect 69348 3108 69354 3120
rect 69477 3111 69535 3117
rect 69477 3108 69489 3111
rect 69348 3080 69489 3108
rect 69348 3068 69354 3080
rect 69477 3077 69489 3080
rect 69523 3108 69535 3111
rect 69569 3111 69627 3117
rect 69569 3108 69581 3111
rect 69523 3080 69581 3108
rect 69523 3077 69535 3080
rect 69477 3071 69535 3077
rect 69569 3077 69581 3080
rect 69615 3077 69627 3111
rect 69569 3071 69627 3077
rect 70026 3068 70032 3120
rect 70084 3108 70090 3120
rect 70084 3080 71820 3108
rect 70084 3068 70090 3080
rect 13924 3012 15332 3040
rect 13906 2932 13912 2984
rect 13964 2972 13970 2984
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13964 2944 14197 2972
rect 13964 2932 13970 2944
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 15010 2972 15016 2984
rect 14971 2944 15016 2972
rect 14185 2935 14243 2941
rect 15010 2932 15016 2944
rect 15068 2932 15074 2984
rect 15304 2904 15332 3012
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 17497 3043 17555 3049
rect 17497 3040 17509 3043
rect 17460 3012 17509 3040
rect 17460 3000 17466 3012
rect 17497 3009 17509 3012
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 18506 3000 18512 3052
rect 18564 3040 18570 3052
rect 34698 3040 34704 3052
rect 18564 3012 34704 3040
rect 18564 3000 18570 3012
rect 34698 3000 34704 3012
rect 34756 3000 34762 3052
rect 35526 3040 35532 3052
rect 35487 3012 35532 3040
rect 35526 3000 35532 3012
rect 35584 3000 35590 3052
rect 42150 3040 42156 3052
rect 36372 3012 42156 3040
rect 15746 2972 15752 2984
rect 15707 2944 15752 2972
rect 15746 2932 15752 2944
rect 15804 2932 15810 2984
rect 16942 2932 16948 2984
rect 17000 2972 17006 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 17000 2944 17325 2972
rect 17000 2932 17006 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 18233 2975 18291 2981
rect 18233 2972 18245 2975
rect 18196 2944 18245 2972
rect 18196 2932 18202 2944
rect 18233 2941 18245 2944
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 18782 2932 18788 2984
rect 18840 2972 18846 2984
rect 19153 2975 19211 2981
rect 19153 2972 19165 2975
rect 18840 2944 19165 2972
rect 18840 2932 18846 2944
rect 19153 2941 19165 2944
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 20073 2975 20131 2981
rect 20073 2972 20085 2975
rect 19392 2944 20085 2972
rect 19392 2932 19398 2944
rect 20073 2941 20085 2944
rect 20119 2941 20131 2975
rect 20073 2935 20131 2941
rect 20162 2932 20168 2984
rect 20220 2972 20226 2984
rect 22094 2972 22100 2984
rect 20220 2944 22100 2972
rect 20220 2932 20226 2944
rect 22094 2932 22100 2944
rect 22152 2932 22158 2984
rect 22186 2932 22192 2984
rect 22244 2972 22250 2984
rect 23293 2975 23351 2981
rect 23293 2972 23305 2975
rect 22244 2944 23305 2972
rect 22244 2932 22250 2944
rect 23293 2941 23305 2944
rect 23339 2941 23351 2975
rect 23293 2935 23351 2941
rect 23474 2932 23480 2984
rect 23532 2972 23538 2984
rect 23937 2975 23995 2981
rect 23937 2972 23949 2975
rect 23532 2944 23949 2972
rect 23532 2932 23538 2944
rect 23937 2941 23949 2944
rect 23983 2941 23995 2975
rect 23937 2935 23995 2941
rect 25041 2975 25099 2981
rect 25041 2941 25053 2975
rect 25087 2972 25099 2975
rect 25130 2972 25136 2984
rect 25087 2944 25136 2972
rect 25087 2941 25099 2944
rect 25041 2935 25099 2941
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 25590 2972 25596 2984
rect 25551 2944 25596 2972
rect 25590 2932 25596 2944
rect 25648 2932 25654 2984
rect 26970 2972 26976 2984
rect 25700 2944 26976 2972
rect 18046 2904 18052 2916
rect 13832 2876 15240 2904
rect 15304 2876 18052 2904
rect 2498 2796 2504 2848
rect 2556 2836 2562 2848
rect 3418 2836 3424 2848
rect 2556 2808 3424 2836
rect 2556 2796 2562 2808
rect 3418 2796 3424 2808
rect 3476 2796 3482 2848
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2836 9275 2839
rect 9306 2836 9312 2848
rect 9263 2808 9312 2836
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 13446 2796 13452 2848
rect 13504 2836 13510 2848
rect 15105 2839 15163 2845
rect 15105 2836 15117 2839
rect 13504 2808 15117 2836
rect 13504 2796 13510 2808
rect 15105 2805 15117 2808
rect 15151 2805 15163 2839
rect 15212 2836 15240 2876
rect 18046 2864 18052 2876
rect 18104 2864 18110 2916
rect 18509 2907 18567 2913
rect 18509 2873 18521 2907
rect 18555 2904 18567 2907
rect 18690 2904 18696 2916
rect 18555 2876 18696 2904
rect 18555 2873 18567 2876
rect 18509 2867 18567 2873
rect 18690 2864 18696 2876
rect 18748 2864 18754 2916
rect 19429 2907 19487 2913
rect 19429 2873 19441 2907
rect 19475 2904 19487 2907
rect 20438 2904 20444 2916
rect 19475 2876 20444 2904
rect 19475 2873 19487 2876
rect 19429 2867 19487 2873
rect 20438 2864 20444 2876
rect 20496 2864 20502 2916
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 20901 2907 20959 2913
rect 20901 2904 20913 2907
rect 20680 2876 20913 2904
rect 20680 2864 20686 2876
rect 20901 2873 20913 2876
rect 20947 2873 20959 2907
rect 22005 2907 22063 2913
rect 22005 2904 22017 2907
rect 20901 2867 20959 2873
rect 21008 2876 22017 2904
rect 19978 2836 19984 2848
rect 15212 2808 19984 2836
rect 15105 2799 15163 2805
rect 19978 2796 19984 2808
rect 20036 2796 20042 2848
rect 20070 2796 20076 2848
rect 20128 2836 20134 2848
rect 21008 2836 21036 2876
rect 22005 2873 22017 2876
rect 22051 2873 22063 2907
rect 22005 2867 22063 2873
rect 22649 2907 22707 2913
rect 22649 2873 22661 2907
rect 22695 2904 22707 2907
rect 22695 2876 24808 2904
rect 22695 2873 22707 2876
rect 22649 2867 22707 2873
rect 20128 2808 21036 2836
rect 20128 2796 20134 2808
rect 21358 2796 21364 2848
rect 21416 2836 21422 2848
rect 22741 2839 22799 2845
rect 22741 2836 22753 2839
rect 21416 2808 22753 2836
rect 21416 2796 21422 2808
rect 22741 2805 22753 2808
rect 22787 2805 22799 2839
rect 24780 2836 24808 2876
rect 24854 2864 24860 2916
rect 24912 2904 24918 2916
rect 25700 2904 25728 2944
rect 26970 2932 26976 2944
rect 27028 2932 27034 2984
rect 27614 2972 27620 2984
rect 27575 2944 27620 2972
rect 27614 2932 27620 2944
rect 27672 2972 27678 2984
rect 27985 2975 28043 2981
rect 27985 2972 27997 2975
rect 27672 2944 27997 2972
rect 27672 2932 27678 2944
rect 27985 2941 27997 2944
rect 28031 2941 28043 2975
rect 27985 2935 28043 2941
rect 28353 2975 28411 2981
rect 28353 2941 28365 2975
rect 28399 2972 28411 2975
rect 28721 2975 28779 2981
rect 28721 2972 28733 2975
rect 28399 2944 28733 2972
rect 28399 2941 28411 2944
rect 28353 2935 28411 2941
rect 28721 2941 28733 2944
rect 28767 2972 28779 2975
rect 28810 2972 28816 2984
rect 28767 2944 28816 2972
rect 28767 2941 28779 2944
rect 28721 2935 28779 2941
rect 28810 2932 28816 2944
rect 28868 2932 28874 2984
rect 29181 2975 29239 2981
rect 29181 2941 29193 2975
rect 29227 2941 29239 2975
rect 29181 2935 29239 2941
rect 24912 2876 25728 2904
rect 24912 2864 24918 2876
rect 26234 2864 26240 2916
rect 26292 2904 26298 2916
rect 26329 2907 26387 2913
rect 26329 2904 26341 2907
rect 26292 2876 26341 2904
rect 26292 2864 26298 2876
rect 26329 2873 26341 2876
rect 26375 2873 26387 2907
rect 26329 2867 26387 2873
rect 27338 2864 27344 2916
rect 27396 2904 27402 2916
rect 27801 2907 27859 2913
rect 27801 2904 27813 2907
rect 27396 2876 27813 2904
rect 27396 2864 27402 2876
rect 27801 2873 27813 2876
rect 27847 2873 27859 2907
rect 27801 2867 27859 2873
rect 28442 2864 28448 2916
rect 28500 2904 28506 2916
rect 29196 2904 29224 2935
rect 29546 2932 29552 2984
rect 29604 2972 29610 2984
rect 29825 2975 29883 2981
rect 29825 2972 29837 2975
rect 29604 2944 29837 2972
rect 29604 2932 29610 2944
rect 29825 2941 29837 2944
rect 29871 2941 29883 2975
rect 29825 2935 29883 2941
rect 30098 2932 30104 2984
rect 30156 2972 30162 2984
rect 30469 2975 30527 2981
rect 30469 2972 30481 2975
rect 30156 2944 30481 2972
rect 30156 2932 30162 2944
rect 30469 2941 30481 2944
rect 30515 2941 30527 2975
rect 30469 2935 30527 2941
rect 30742 2932 30748 2984
rect 30800 2972 30806 2984
rect 31113 2975 31171 2981
rect 31113 2972 31125 2975
rect 30800 2944 31125 2972
rect 30800 2932 30806 2944
rect 31113 2941 31125 2944
rect 31159 2941 31171 2975
rect 31113 2935 31171 2941
rect 31386 2932 31392 2984
rect 31444 2972 31450 2984
rect 31757 2975 31815 2981
rect 31757 2972 31769 2975
rect 31444 2944 31769 2972
rect 31444 2932 31450 2944
rect 31757 2941 31769 2944
rect 31803 2941 31815 2975
rect 31757 2935 31815 2941
rect 32582 2932 32588 2984
rect 32640 2972 32646 2984
rect 33045 2975 33103 2981
rect 33045 2972 33057 2975
rect 32640 2944 33057 2972
rect 32640 2932 32646 2944
rect 33045 2941 33057 2944
rect 33091 2941 33103 2975
rect 33045 2935 33103 2941
rect 33226 2932 33232 2984
rect 33284 2972 33290 2984
rect 33689 2975 33747 2981
rect 33689 2972 33701 2975
rect 33284 2944 33701 2972
rect 33284 2932 33290 2944
rect 33689 2941 33701 2944
rect 33735 2941 33747 2975
rect 33689 2935 33747 2941
rect 33778 2932 33784 2984
rect 33836 2972 33842 2984
rect 34333 2975 34391 2981
rect 34333 2972 34345 2975
rect 33836 2944 34345 2972
rect 33836 2932 33842 2944
rect 34333 2941 34345 2944
rect 34379 2941 34391 2975
rect 35342 2972 35348 2984
rect 35303 2944 35348 2972
rect 34333 2935 34391 2941
rect 35342 2932 35348 2944
rect 35400 2932 35406 2984
rect 36372 2981 36400 3012
rect 42150 3000 42156 3012
rect 42208 3000 42214 3052
rect 42426 3000 42432 3052
rect 42484 3040 42490 3052
rect 46937 3043 46995 3049
rect 42484 3012 45876 3040
rect 42484 3000 42490 3012
rect 36357 2975 36415 2981
rect 36357 2941 36369 2975
rect 36403 2941 36415 2975
rect 36357 2935 36415 2941
rect 37001 2975 37059 2981
rect 37001 2941 37013 2975
rect 37047 2941 37059 2975
rect 37001 2935 37059 2941
rect 28500 2876 29224 2904
rect 28500 2864 28506 2876
rect 34606 2864 34612 2916
rect 34664 2904 34670 2916
rect 36170 2904 36176 2916
rect 34664 2876 36176 2904
rect 34664 2864 34670 2876
rect 36170 2864 36176 2876
rect 36228 2864 36234 2916
rect 36262 2864 36268 2916
rect 36320 2904 36326 2916
rect 37016 2904 37044 2935
rect 37458 2932 37464 2984
rect 37516 2972 37522 2984
rect 39025 2975 39083 2981
rect 39025 2972 39037 2975
rect 37516 2944 39037 2972
rect 37516 2932 37522 2944
rect 39025 2941 39037 2944
rect 39071 2941 39083 2975
rect 39025 2935 39083 2941
rect 39482 2932 39488 2984
rect 39540 2972 39546 2984
rect 40221 2975 40279 2981
rect 40221 2972 40233 2975
rect 39540 2944 40233 2972
rect 39540 2932 39546 2944
rect 40221 2941 40233 2944
rect 40267 2941 40279 2975
rect 40221 2935 40279 2941
rect 41138 2932 41144 2984
rect 41196 2972 41202 2984
rect 42061 2975 42119 2981
rect 42061 2972 42073 2975
rect 41196 2944 42073 2972
rect 41196 2932 41202 2944
rect 42061 2941 42073 2944
rect 42107 2941 42119 2975
rect 42061 2935 42119 2941
rect 43530 2932 43536 2984
rect 43588 2972 43594 2984
rect 44269 2975 44327 2981
rect 44269 2972 44281 2975
rect 43588 2944 44281 2972
rect 43588 2932 43594 2944
rect 44269 2941 44281 2944
rect 44315 2941 44327 2975
rect 44269 2935 44327 2941
rect 44913 2975 44971 2981
rect 44913 2941 44925 2975
rect 44959 2941 44971 2975
rect 44913 2935 44971 2941
rect 45465 2975 45523 2981
rect 45465 2941 45477 2975
rect 45511 2972 45523 2975
rect 45738 2972 45744 2984
rect 45511 2944 45744 2972
rect 45511 2941 45523 2944
rect 45465 2935 45523 2941
rect 36320 2876 37044 2904
rect 36320 2864 36326 2876
rect 37642 2864 37648 2916
rect 37700 2904 37706 2916
rect 38289 2907 38347 2913
rect 38289 2904 38301 2907
rect 37700 2876 38301 2904
rect 37700 2864 37706 2876
rect 38289 2873 38301 2876
rect 38335 2873 38347 2907
rect 38289 2867 38347 2873
rect 38473 2907 38531 2913
rect 38473 2873 38485 2907
rect 38519 2873 38531 2907
rect 38473 2867 38531 2873
rect 41417 2907 41475 2913
rect 41417 2873 41429 2907
rect 41463 2904 41475 2907
rect 41598 2904 41604 2916
rect 41463 2876 41604 2904
rect 41463 2873 41475 2876
rect 41417 2867 41475 2873
rect 25222 2836 25228 2848
rect 24780 2808 25228 2836
rect 22741 2799 22799 2805
rect 25222 2796 25228 2808
rect 25280 2796 25286 2848
rect 25498 2796 25504 2848
rect 25556 2836 25562 2848
rect 25685 2839 25743 2845
rect 25685 2836 25697 2839
rect 25556 2808 25697 2836
rect 25556 2796 25562 2808
rect 25685 2805 25697 2808
rect 25731 2805 25743 2839
rect 25685 2799 25743 2805
rect 26142 2796 26148 2848
rect 26200 2836 26206 2848
rect 26421 2839 26479 2845
rect 26421 2836 26433 2839
rect 26200 2808 26433 2836
rect 26200 2796 26206 2808
rect 26421 2805 26433 2808
rect 26467 2805 26479 2839
rect 26421 2799 26479 2805
rect 35526 2796 35532 2848
rect 35584 2836 35590 2848
rect 35710 2836 35716 2848
rect 35584 2808 35716 2836
rect 35584 2796 35590 2808
rect 35710 2796 35716 2808
rect 35768 2796 35774 2848
rect 35802 2796 35808 2848
rect 35860 2836 35866 2848
rect 36449 2839 36507 2845
rect 36449 2836 36461 2839
rect 35860 2808 36461 2836
rect 35860 2796 35866 2808
rect 36449 2805 36461 2808
rect 36495 2805 36507 2839
rect 36449 2799 36507 2805
rect 38010 2796 38016 2848
rect 38068 2836 38074 2848
rect 38488 2836 38516 2867
rect 41598 2864 41604 2876
rect 41656 2864 41662 2916
rect 43622 2904 43628 2916
rect 43583 2876 43628 2904
rect 43622 2864 43628 2876
rect 43680 2864 43686 2916
rect 44174 2864 44180 2916
rect 44232 2904 44238 2916
rect 44928 2904 44956 2935
rect 45738 2932 45744 2944
rect 45796 2932 45802 2984
rect 45554 2904 45560 2916
rect 44232 2876 44956 2904
rect 45515 2876 45560 2904
rect 44232 2864 44238 2876
rect 45554 2864 45560 2876
rect 45612 2864 45618 2916
rect 45848 2904 45876 3012
rect 46937 3009 46949 3043
rect 46983 3040 46995 3043
rect 46983 3012 47256 3040
rect 46983 3009 46995 3012
rect 46937 3003 46995 3009
rect 46198 2932 46204 2984
rect 46256 2972 46262 2984
rect 46385 2975 46443 2981
rect 46385 2972 46397 2975
rect 46256 2944 46397 2972
rect 46256 2932 46262 2944
rect 46385 2941 46397 2944
rect 46431 2941 46443 2975
rect 46385 2935 46443 2941
rect 46842 2932 46848 2984
rect 46900 2972 46906 2984
rect 47228 2981 47256 3012
rect 49050 3000 49056 3052
rect 49108 3040 49114 3052
rect 49108 3012 50292 3040
rect 49108 3000 49114 3012
rect 47029 2975 47087 2981
rect 47029 2972 47041 2975
rect 46900 2944 47041 2972
rect 46900 2932 46906 2944
rect 47029 2941 47041 2944
rect 47075 2941 47087 2975
rect 47029 2935 47087 2941
rect 47213 2975 47271 2981
rect 47213 2941 47225 2975
rect 47259 2972 47271 2975
rect 48130 2972 48136 2984
rect 47259 2944 48136 2972
rect 47259 2941 47271 2944
rect 47213 2935 47271 2941
rect 48130 2932 48136 2944
rect 48188 2932 48194 2984
rect 48869 2975 48927 2981
rect 48869 2941 48881 2975
rect 48915 2972 48927 2975
rect 49142 2972 49148 2984
rect 48915 2944 49148 2972
rect 48915 2941 48927 2944
rect 48869 2935 48927 2941
rect 49142 2932 49148 2944
rect 49200 2932 49206 2984
rect 49421 2975 49479 2981
rect 49421 2941 49433 2975
rect 49467 2972 49479 2975
rect 49697 2975 49755 2981
rect 49697 2972 49709 2975
rect 49467 2944 49709 2972
rect 49467 2941 49479 2944
rect 49421 2935 49479 2941
rect 49697 2941 49709 2944
rect 49743 2972 49755 2975
rect 49786 2972 49792 2984
rect 49743 2944 49792 2972
rect 49743 2941 49755 2944
rect 49697 2935 49755 2941
rect 49786 2932 49792 2944
rect 49844 2932 49850 2984
rect 50264 2981 50292 3012
rect 50798 3000 50804 3052
rect 50856 3040 50862 3052
rect 50982 3040 50988 3052
rect 50856 3012 50988 3040
rect 50856 3000 50862 3012
rect 50982 3000 50988 3012
rect 51040 3000 51046 3052
rect 55214 3040 55220 3052
rect 55175 3012 55220 3040
rect 55214 3000 55220 3012
rect 55272 3040 55278 3052
rect 58342 3040 58348 3052
rect 55272 3012 55536 3040
rect 55272 3000 55278 3012
rect 50249 2975 50307 2981
rect 50249 2941 50261 2975
rect 50295 2941 50307 2975
rect 51813 2975 51871 2981
rect 51813 2972 51825 2975
rect 50249 2935 50307 2941
rect 51046 2944 51825 2972
rect 45848 2876 49096 2904
rect 38068 2808 38516 2836
rect 38068 2796 38074 2808
rect 40126 2796 40132 2848
rect 40184 2836 40190 2848
rect 40313 2839 40371 2845
rect 40313 2836 40325 2839
rect 40184 2808 40325 2836
rect 40184 2796 40190 2808
rect 40313 2805 40325 2808
rect 40359 2805 40371 2839
rect 40313 2799 40371 2805
rect 41230 2796 41236 2848
rect 41288 2836 41294 2848
rect 41509 2839 41567 2845
rect 41509 2836 41521 2839
rect 41288 2808 41521 2836
rect 41288 2796 41294 2808
rect 41509 2805 41521 2808
rect 41555 2805 41567 2839
rect 41509 2799 41567 2805
rect 43162 2796 43168 2848
rect 43220 2836 43226 2848
rect 43717 2839 43775 2845
rect 43717 2836 43729 2839
rect 43220 2808 43729 2836
rect 43220 2796 43226 2808
rect 43717 2805 43729 2808
rect 43763 2805 43775 2839
rect 43717 2799 43775 2805
rect 44358 2796 44364 2848
rect 44416 2836 44422 2848
rect 46106 2836 46112 2848
rect 44416 2808 46112 2836
rect 44416 2796 44422 2808
rect 46106 2796 46112 2808
rect 46164 2796 46170 2848
rect 46198 2796 46204 2848
rect 46256 2836 46262 2848
rect 46477 2839 46535 2845
rect 46477 2836 46489 2839
rect 46256 2808 46489 2836
rect 46256 2796 46262 2808
rect 46477 2805 46489 2808
rect 46523 2805 46535 2839
rect 46477 2799 46535 2805
rect 48038 2796 48044 2848
rect 48096 2836 48102 2848
rect 48961 2839 49019 2845
rect 48961 2836 48973 2839
rect 48096 2808 48973 2836
rect 48096 2796 48102 2808
rect 48961 2805 48973 2808
rect 49007 2805 49019 2839
rect 49068 2836 49096 2876
rect 49234 2864 49240 2916
rect 49292 2904 49298 2916
rect 49513 2907 49571 2913
rect 49513 2904 49525 2907
rect 49292 2876 49525 2904
rect 49292 2864 49298 2876
rect 49513 2873 49525 2876
rect 49559 2873 49571 2907
rect 49513 2867 49571 2873
rect 50154 2864 50160 2916
rect 50212 2904 50218 2916
rect 51046 2904 51074 2944
rect 51813 2941 51825 2944
rect 51859 2941 51871 2975
rect 51813 2935 51871 2941
rect 52457 2975 52515 2981
rect 52457 2941 52469 2975
rect 52503 2941 52515 2975
rect 52457 2935 52515 2941
rect 50212 2876 51074 2904
rect 51169 2907 51227 2913
rect 50212 2864 50218 2876
rect 51169 2873 51181 2907
rect 51215 2904 51227 2907
rect 51350 2904 51356 2916
rect 51215 2876 51356 2904
rect 51215 2873 51227 2876
rect 51169 2867 51227 2873
rect 51350 2864 51356 2876
rect 51408 2864 51414 2916
rect 51442 2864 51448 2916
rect 51500 2904 51506 2916
rect 52472 2904 52500 2935
rect 54018 2932 54024 2984
rect 54076 2972 54082 2984
rect 55508 2981 55536 3012
rect 55600 3012 58348 3040
rect 54113 2975 54171 2981
rect 54113 2972 54125 2975
rect 54076 2944 54125 2972
rect 54076 2932 54082 2944
rect 54113 2941 54125 2944
rect 54159 2941 54171 2975
rect 54113 2935 54171 2941
rect 55493 2975 55551 2981
rect 55493 2941 55505 2975
rect 55539 2941 55551 2975
rect 55493 2935 55551 2941
rect 55306 2904 55312 2916
rect 51500 2876 52500 2904
rect 55267 2876 55312 2904
rect 51500 2864 51506 2876
rect 55306 2864 55312 2876
rect 55364 2864 55370 2916
rect 49602 2836 49608 2848
rect 49068 2808 49608 2836
rect 48961 2799 49019 2805
rect 49602 2796 49608 2808
rect 49660 2796 49666 2848
rect 49786 2796 49792 2848
rect 49844 2836 49850 2848
rect 49970 2836 49976 2848
rect 49844 2808 49976 2836
rect 49844 2796 49850 2808
rect 49970 2796 49976 2808
rect 50028 2796 50034 2848
rect 51074 2796 51080 2848
rect 51132 2836 51138 2848
rect 51261 2839 51319 2845
rect 51261 2836 51273 2839
rect 51132 2808 51273 2836
rect 51132 2796 51138 2808
rect 51261 2805 51273 2808
rect 51307 2805 51319 2839
rect 51261 2799 51319 2805
rect 53558 2796 53564 2848
rect 53616 2836 53622 2848
rect 54205 2839 54263 2845
rect 54205 2836 54217 2839
rect 53616 2808 54217 2836
rect 53616 2796 53622 2808
rect 54205 2805 54217 2808
rect 54251 2805 54263 2839
rect 54205 2799 54263 2805
rect 54754 2796 54760 2848
rect 54812 2836 54818 2848
rect 55600 2836 55628 3012
rect 58342 3000 58348 3012
rect 58400 3000 58406 3052
rect 60826 3000 60832 3052
rect 60884 3040 60890 3052
rect 64414 3040 64420 3052
rect 60884 3012 64420 3040
rect 60884 3000 60890 3012
rect 64414 3000 64420 3012
rect 64472 3000 64478 3052
rect 56686 2972 56692 2984
rect 56647 2944 56692 2972
rect 56686 2932 56692 2944
rect 56744 2932 56750 2984
rect 57333 2975 57391 2981
rect 57333 2941 57345 2975
rect 57379 2941 57391 2975
rect 57333 2935 57391 2941
rect 55766 2864 55772 2916
rect 55824 2904 55830 2916
rect 57348 2904 57376 2935
rect 57606 2932 57612 2984
rect 57664 2972 57670 2984
rect 57977 2975 58035 2981
rect 57977 2972 57989 2975
rect 57664 2944 57989 2972
rect 57664 2932 57670 2944
rect 57977 2941 57989 2944
rect 58023 2941 58035 2975
rect 59354 2972 59360 2984
rect 59315 2944 59360 2972
rect 57977 2935 58035 2941
rect 59354 2932 59360 2944
rect 59412 2932 59418 2984
rect 59446 2932 59452 2984
rect 59504 2972 59510 2984
rect 60001 2975 60059 2981
rect 60001 2972 60013 2975
rect 59504 2944 60013 2972
rect 59504 2932 59510 2944
rect 60001 2941 60013 2944
rect 60047 2941 60059 2975
rect 60001 2935 60059 2941
rect 60090 2932 60096 2984
rect 60148 2972 60154 2984
rect 60645 2975 60703 2981
rect 60645 2972 60657 2975
rect 60148 2944 60657 2972
rect 60148 2932 60154 2944
rect 60645 2941 60657 2944
rect 60691 2941 60703 2975
rect 60645 2935 60703 2941
rect 60918 2932 60924 2984
rect 60976 2972 60982 2984
rect 62114 2972 62120 2984
rect 60976 2944 62120 2972
rect 60976 2932 60982 2944
rect 62114 2932 62120 2944
rect 62172 2932 62178 2984
rect 62758 2972 62764 2984
rect 62719 2944 62764 2972
rect 62758 2932 62764 2944
rect 62816 2932 62822 2984
rect 63586 2972 63592 2984
rect 63547 2944 63592 2972
rect 63586 2932 63592 2944
rect 63644 2932 63650 2984
rect 64322 2932 64328 2984
rect 64380 2972 64386 2984
rect 65245 2975 65303 2981
rect 65245 2972 65257 2975
rect 64380 2944 65257 2972
rect 64380 2932 64386 2944
rect 65245 2941 65257 2944
rect 65291 2941 65303 2975
rect 65245 2935 65303 2941
rect 65518 2932 65524 2984
rect 65576 2972 65582 2984
rect 65889 2975 65947 2981
rect 65889 2972 65901 2975
rect 65576 2944 65901 2972
rect 65576 2932 65582 2944
rect 65889 2941 65901 2944
rect 65935 2941 65947 2975
rect 66824 2972 66852 3068
rect 67266 3000 67272 3052
rect 67324 3040 67330 3052
rect 67324 3012 70072 3040
rect 67324 3000 67330 3012
rect 67085 2975 67143 2981
rect 67085 2972 67097 2975
rect 66824 2944 67097 2972
rect 65889 2935 65947 2941
rect 67085 2941 67097 2944
rect 67131 2941 67143 2975
rect 67637 2975 67695 2981
rect 67637 2972 67649 2975
rect 67085 2935 67143 2941
rect 67192 2944 67649 2972
rect 55824 2876 57376 2904
rect 55824 2864 55830 2876
rect 57790 2864 57796 2916
rect 57848 2904 57854 2916
rect 60274 2904 60280 2916
rect 57848 2876 60280 2904
rect 57848 2864 57854 2876
rect 60274 2864 60280 2876
rect 60332 2864 60338 2916
rect 61562 2904 61568 2916
rect 61523 2876 61568 2904
rect 61562 2864 61568 2876
rect 61620 2864 61626 2916
rect 64506 2904 64512 2916
rect 64467 2876 64512 2904
rect 64506 2864 64512 2876
rect 64564 2864 64570 2916
rect 64690 2904 64696 2916
rect 64651 2876 64696 2904
rect 64690 2864 64696 2876
rect 64748 2864 64754 2916
rect 66898 2904 66904 2916
rect 66859 2876 66904 2904
rect 66898 2864 66904 2876
rect 66956 2864 66962 2916
rect 54812 2808 55628 2836
rect 54812 2796 54818 2808
rect 56594 2796 56600 2848
rect 56652 2836 56658 2848
rect 56781 2839 56839 2845
rect 56781 2836 56793 2839
rect 56652 2808 56793 2836
rect 56652 2796 56658 2808
rect 56781 2805 56793 2808
rect 56827 2805 56839 2839
rect 56781 2799 56839 2805
rect 58986 2796 58992 2848
rect 59044 2836 59050 2848
rect 59449 2839 59507 2845
rect 59449 2836 59461 2839
rect 59044 2808 59461 2836
rect 59044 2796 59050 2808
rect 59449 2805 59461 2808
rect 59495 2805 59507 2839
rect 59449 2799 59507 2805
rect 61470 2796 61476 2848
rect 61528 2836 61534 2848
rect 61657 2839 61715 2845
rect 61657 2836 61669 2839
rect 61528 2808 61669 2836
rect 61528 2796 61534 2808
rect 61657 2805 61669 2808
rect 61703 2805 61715 2839
rect 61657 2799 61715 2805
rect 62666 2796 62672 2848
rect 62724 2836 62730 2848
rect 62853 2839 62911 2845
rect 62853 2836 62865 2839
rect 62724 2808 62865 2836
rect 62724 2796 62730 2808
rect 62853 2805 62865 2808
rect 62899 2805 62911 2839
rect 62853 2799 62911 2805
rect 64417 2839 64475 2845
rect 64417 2805 64429 2839
rect 64463 2836 64475 2839
rect 64708 2836 64736 2864
rect 64463 2808 64736 2836
rect 64463 2805 64475 2808
rect 64417 2799 64475 2805
rect 66162 2796 66168 2848
rect 66220 2836 66226 2848
rect 67192 2836 67220 2944
rect 67637 2941 67649 2944
rect 67683 2941 67695 2975
rect 67637 2935 67695 2941
rect 68281 2975 68339 2981
rect 68281 2941 68293 2975
rect 68327 2941 68339 2975
rect 68281 2935 68339 2941
rect 69477 2975 69535 2981
rect 69477 2941 69489 2975
rect 69523 2972 69535 2975
rect 69937 2975 69995 2981
rect 69937 2972 69949 2975
rect 69523 2944 69949 2972
rect 69523 2941 69535 2944
rect 69477 2935 69535 2941
rect 69937 2941 69949 2944
rect 69983 2941 69995 2975
rect 70044 2972 70072 3012
rect 70118 3000 70124 3052
rect 70176 3040 70182 3052
rect 71593 3043 71651 3049
rect 71593 3040 71605 3043
rect 70176 3012 71605 3040
rect 70176 3000 70182 3012
rect 71593 3009 71605 3012
rect 71639 3009 71651 3043
rect 71593 3003 71651 3009
rect 70489 2975 70547 2981
rect 70489 2972 70501 2975
rect 70044 2944 70501 2972
rect 69937 2935 69995 2941
rect 70489 2941 70501 2944
rect 70535 2972 70547 2975
rect 70765 2975 70823 2981
rect 70765 2972 70777 2975
rect 70535 2944 70777 2972
rect 70535 2941 70547 2944
rect 70489 2935 70547 2941
rect 70765 2941 70777 2944
rect 70811 2941 70823 2975
rect 71314 2972 71320 2984
rect 71275 2944 71320 2972
rect 70765 2935 70823 2941
rect 67358 2864 67364 2916
rect 67416 2904 67422 2916
rect 68296 2904 68324 2935
rect 71314 2932 71320 2944
rect 71372 2932 71378 2984
rect 71498 2932 71504 2984
rect 71556 2972 71562 2984
rect 71685 2975 71743 2981
rect 71556 2944 71600 2972
rect 71556 2932 71562 2944
rect 71685 2941 71697 2975
rect 71731 2941 71743 2975
rect 71685 2935 71743 2941
rect 67416 2876 68324 2904
rect 67416 2864 67422 2876
rect 69382 2864 69388 2916
rect 69440 2904 69446 2916
rect 69753 2907 69811 2913
rect 69753 2904 69765 2907
rect 69440 2876 69765 2904
rect 69440 2864 69446 2876
rect 69753 2873 69765 2876
rect 69799 2873 69811 2907
rect 70578 2904 70584 2916
rect 70539 2876 70584 2904
rect 69753 2867 69811 2873
rect 70578 2864 70584 2876
rect 70636 2864 70642 2916
rect 70854 2864 70860 2916
rect 70912 2904 70918 2916
rect 71700 2904 71728 2935
rect 70912 2876 71728 2904
rect 71792 2904 71820 3080
rect 74902 3000 74908 3052
rect 74960 3040 74966 3052
rect 78508 3040 78536 3136
rect 81544 3040 81572 3139
rect 81802 3136 81808 3188
rect 81860 3176 81866 3188
rect 82906 3176 82912 3188
rect 81860 3148 82912 3176
rect 81860 3136 81866 3148
rect 82906 3136 82912 3148
rect 82964 3136 82970 3188
rect 83458 3136 83464 3188
rect 83516 3176 83522 3188
rect 85669 3179 85727 3185
rect 85669 3176 85681 3179
rect 83516 3148 85681 3176
rect 83516 3136 83522 3148
rect 85669 3145 85681 3148
rect 85715 3176 85727 3179
rect 85942 3176 85948 3188
rect 85715 3148 85948 3176
rect 85715 3145 85727 3148
rect 85669 3139 85727 3145
rect 85942 3136 85948 3148
rect 86000 3136 86006 3188
rect 88334 3136 88340 3188
rect 88392 3176 88398 3188
rect 89073 3179 89131 3185
rect 89073 3176 89085 3179
rect 88392 3148 89085 3176
rect 88392 3136 88398 3148
rect 89073 3145 89085 3148
rect 89119 3145 89131 3179
rect 89073 3139 89131 3145
rect 89990 3136 89996 3188
rect 90048 3176 90054 3188
rect 90453 3179 90511 3185
rect 90453 3176 90465 3179
rect 90048 3148 90465 3176
rect 90048 3136 90054 3148
rect 90453 3145 90465 3148
rect 90499 3176 90511 3179
rect 90545 3179 90603 3185
rect 90545 3176 90557 3179
rect 90499 3148 90557 3176
rect 90499 3145 90511 3148
rect 90453 3139 90511 3145
rect 90545 3145 90557 3148
rect 90591 3145 90603 3179
rect 94406 3176 94412 3188
rect 94367 3148 94412 3176
rect 90545 3139 90603 3145
rect 94406 3136 94412 3148
rect 94464 3136 94470 3188
rect 95786 3176 95792 3188
rect 95747 3148 95792 3176
rect 95786 3136 95792 3148
rect 95844 3136 95850 3188
rect 96062 3136 96068 3188
rect 96120 3176 96126 3188
rect 97261 3179 97319 3185
rect 97261 3176 97273 3179
rect 96120 3148 97273 3176
rect 96120 3136 96126 3148
rect 97261 3145 97273 3148
rect 97307 3145 97319 3179
rect 97261 3139 97319 3145
rect 92198 3068 92204 3120
rect 92256 3108 92262 3120
rect 92934 3108 92940 3120
rect 92256 3080 92940 3108
rect 92256 3068 92262 3080
rect 92934 3068 92940 3080
rect 92992 3068 92998 3120
rect 94424 3040 94452 3136
rect 74960 3012 76972 3040
rect 78508 3012 78904 3040
rect 81544 3012 81940 3040
rect 74960 3000 74966 3012
rect 71866 2932 71872 2984
rect 71924 2972 71930 2984
rect 71924 2944 71969 2972
rect 71924 2932 71930 2944
rect 72234 2932 72240 2984
rect 72292 2972 72298 2984
rect 73249 2975 73307 2981
rect 73249 2972 73261 2975
rect 72292 2944 73261 2972
rect 72292 2932 72298 2944
rect 73249 2941 73261 2944
rect 73295 2941 73307 2975
rect 73249 2935 73307 2941
rect 73430 2932 73436 2984
rect 73488 2972 73494 2984
rect 73893 2975 73951 2981
rect 73893 2972 73905 2975
rect 73488 2944 73905 2972
rect 73488 2932 73494 2944
rect 73893 2941 73905 2944
rect 73939 2941 73951 2975
rect 73893 2935 73951 2941
rect 74810 2932 74816 2984
rect 74868 2972 74874 2984
rect 75181 2975 75239 2981
rect 75181 2972 75193 2975
rect 74868 2944 75193 2972
rect 74868 2932 74874 2944
rect 75181 2941 75193 2944
rect 75227 2941 75239 2975
rect 75181 2935 75239 2941
rect 75270 2932 75276 2984
rect 75328 2972 75334 2984
rect 75733 2975 75791 2981
rect 75733 2972 75745 2975
rect 75328 2944 75745 2972
rect 75328 2932 75334 2944
rect 75733 2941 75745 2944
rect 75779 2941 75791 2975
rect 75733 2935 75791 2941
rect 76377 2975 76435 2981
rect 76377 2941 76389 2975
rect 76423 2972 76435 2975
rect 76837 2975 76895 2981
rect 76837 2972 76849 2975
rect 76423 2944 76849 2972
rect 76423 2941 76435 2944
rect 76377 2935 76435 2941
rect 76837 2941 76849 2944
rect 76883 2941 76895 2975
rect 76837 2935 76895 2941
rect 72605 2907 72663 2913
rect 72605 2904 72617 2907
rect 71792 2876 72617 2904
rect 70912 2864 70918 2876
rect 72605 2873 72617 2876
rect 72651 2873 72663 2907
rect 72605 2867 72663 2873
rect 74902 2864 74908 2916
rect 74960 2904 74966 2916
rect 74997 2907 75055 2913
rect 74997 2904 75009 2907
rect 74960 2876 75009 2904
rect 74960 2864 74966 2876
rect 74997 2873 75009 2876
rect 75043 2873 75055 2907
rect 76650 2904 76656 2916
rect 76611 2876 76656 2904
rect 74997 2867 75055 2873
rect 76650 2864 76656 2876
rect 76708 2864 76714 2916
rect 76944 2904 76972 3012
rect 77570 2932 77576 2984
rect 77628 2972 77634 2984
rect 78033 2975 78091 2981
rect 78033 2972 78045 2975
rect 77628 2944 78045 2972
rect 77628 2932 77634 2944
rect 78033 2941 78045 2944
rect 78079 2941 78091 2975
rect 78033 2935 78091 2941
rect 78490 2932 78496 2984
rect 78548 2972 78554 2984
rect 78876 2981 78904 3012
rect 78677 2975 78735 2981
rect 78677 2972 78689 2975
rect 78548 2944 78689 2972
rect 78548 2932 78554 2944
rect 78677 2941 78689 2944
rect 78723 2941 78735 2975
rect 78677 2935 78735 2941
rect 78861 2975 78919 2981
rect 78861 2941 78873 2975
rect 78907 2941 78919 2975
rect 80149 2975 80207 2981
rect 80149 2972 80161 2975
rect 78861 2935 78919 2941
rect 78968 2944 80161 2972
rect 78968 2904 78996 2944
rect 80149 2941 80161 2944
rect 80195 2972 80207 2975
rect 80425 2975 80483 2981
rect 80425 2972 80437 2975
rect 80195 2944 80437 2972
rect 80195 2941 80207 2944
rect 80149 2935 80207 2941
rect 80425 2941 80437 2944
rect 80471 2941 80483 2975
rect 80425 2935 80483 2941
rect 80882 2932 80888 2984
rect 80940 2972 80946 2984
rect 81912 2981 81940 3012
rect 82556 3012 94360 3040
rect 94424 3012 94820 3040
rect 82556 2981 82584 3012
rect 81713 2975 81771 2981
rect 81713 2972 81725 2975
rect 80940 2944 81725 2972
rect 80940 2932 80946 2944
rect 81713 2941 81725 2944
rect 81759 2941 81771 2975
rect 81713 2935 81771 2941
rect 81897 2975 81955 2981
rect 81897 2941 81909 2975
rect 81943 2941 81955 2975
rect 81897 2935 81955 2941
rect 82541 2975 82599 2981
rect 82541 2941 82553 2975
rect 82587 2941 82599 2975
rect 82541 2935 82599 2941
rect 82630 2932 82636 2984
rect 82688 2972 82694 2984
rect 83185 2975 83243 2981
rect 83185 2972 83197 2975
rect 82688 2944 83197 2972
rect 82688 2932 82694 2944
rect 83185 2941 83197 2944
rect 83231 2941 83243 2975
rect 83185 2935 83243 2941
rect 83274 2932 83280 2984
rect 83332 2972 83338 2984
rect 83829 2975 83887 2981
rect 83829 2972 83841 2975
rect 83332 2944 83841 2972
rect 83332 2932 83338 2944
rect 83829 2941 83841 2944
rect 83875 2941 83887 2975
rect 83829 2935 83887 2941
rect 85666 2932 85672 2984
rect 85724 2972 85730 2984
rect 86589 2975 86647 2981
rect 86589 2972 86601 2975
rect 85724 2944 86601 2972
rect 85724 2932 85730 2944
rect 86589 2941 86601 2944
rect 86635 2941 86647 2975
rect 86589 2935 86647 2941
rect 87598 2932 87604 2984
rect 87656 2972 87662 2984
rect 87693 2975 87751 2981
rect 87693 2972 87705 2975
rect 87656 2944 87705 2972
rect 87656 2932 87662 2944
rect 87693 2941 87705 2944
rect 87739 2941 87751 2975
rect 87966 2972 87972 2984
rect 87927 2944 87972 2972
rect 87693 2935 87751 2941
rect 87966 2932 87972 2944
rect 88024 2932 88030 2984
rect 90453 2975 90511 2981
rect 90453 2941 90465 2975
rect 90499 2972 90511 2975
rect 90913 2975 90971 2981
rect 90913 2972 90925 2975
rect 90499 2944 90925 2972
rect 90499 2941 90511 2944
rect 90453 2935 90511 2941
rect 90913 2941 90925 2944
rect 90959 2941 90971 2975
rect 91554 2972 91560 2984
rect 91515 2944 91560 2972
rect 90913 2935 90971 2941
rect 91554 2932 91560 2944
rect 91612 2932 91618 2984
rect 92290 2972 92296 2984
rect 92251 2944 92296 2972
rect 92290 2932 92296 2944
rect 92348 2932 92354 2984
rect 93946 2972 93952 2984
rect 93907 2944 93952 2972
rect 93946 2932 93952 2944
rect 94004 2932 94010 2984
rect 76944 2876 78996 2904
rect 79778 2864 79784 2916
rect 79836 2904 79842 2916
rect 80241 2907 80299 2913
rect 80241 2904 80253 2907
rect 79836 2876 80253 2904
rect 79836 2864 79842 2876
rect 80241 2873 80253 2876
rect 80287 2873 80299 2907
rect 80241 2867 80299 2873
rect 80330 2864 80336 2916
rect 80388 2904 80394 2916
rect 80977 2907 81035 2913
rect 80977 2904 80989 2907
rect 80388 2876 80989 2904
rect 80388 2864 80394 2876
rect 80977 2873 80989 2876
rect 81023 2873 81035 2907
rect 80977 2867 81035 2873
rect 81161 2907 81219 2913
rect 81161 2873 81173 2907
rect 81207 2873 81219 2907
rect 85850 2904 85856 2916
rect 85811 2876 85856 2904
rect 81161 2867 81219 2873
rect 66220 2808 67220 2836
rect 66220 2796 66226 2808
rect 68186 2796 68192 2848
rect 68244 2836 68250 2848
rect 69290 2836 69296 2848
rect 68244 2808 69296 2836
rect 68244 2796 68250 2808
rect 69290 2796 69296 2808
rect 69348 2796 69354 2848
rect 71958 2836 71964 2848
rect 71919 2808 71964 2836
rect 71958 2796 71964 2808
rect 72016 2796 72022 2848
rect 72418 2796 72424 2848
rect 72476 2836 72482 2848
rect 72697 2839 72755 2845
rect 72697 2836 72709 2839
rect 72476 2808 72709 2836
rect 72476 2796 72482 2808
rect 72697 2805 72709 2808
rect 72743 2805 72755 2839
rect 72697 2799 72755 2805
rect 77938 2796 77944 2848
rect 77996 2836 78002 2848
rect 78125 2839 78183 2845
rect 78125 2836 78137 2839
rect 77996 2808 78137 2836
rect 77996 2796 78002 2808
rect 78125 2805 78137 2808
rect 78171 2805 78183 2839
rect 78125 2799 78183 2805
rect 80701 2839 80759 2845
rect 80701 2805 80713 2839
rect 80747 2836 80759 2839
rect 81176 2836 81204 2867
rect 85850 2864 85856 2876
rect 85908 2864 85914 2916
rect 85942 2864 85948 2916
rect 86000 2904 86006 2916
rect 86037 2907 86095 2913
rect 86037 2904 86049 2907
rect 86000 2876 86049 2904
rect 86000 2864 86006 2876
rect 86037 2873 86049 2876
rect 86083 2873 86095 2907
rect 86037 2867 86095 2873
rect 90082 2864 90088 2916
rect 90140 2904 90146 2916
rect 90729 2907 90787 2913
rect 90729 2904 90741 2907
rect 90140 2876 90741 2904
rect 90140 2864 90146 2876
rect 90729 2873 90741 2876
rect 90775 2873 90787 2907
rect 93118 2904 93124 2916
rect 93079 2876 93124 2904
rect 90729 2867 90787 2873
rect 93118 2864 93124 2876
rect 93176 2864 93182 2916
rect 93305 2907 93363 2913
rect 93305 2873 93317 2907
rect 93351 2873 93363 2907
rect 93305 2867 93363 2873
rect 80747 2808 81204 2836
rect 80747 2805 80759 2808
rect 80701 2799 80759 2805
rect 82170 2796 82176 2848
rect 82228 2836 82234 2848
rect 82633 2839 82691 2845
rect 82633 2836 82645 2839
rect 82228 2808 82645 2836
rect 82228 2796 82234 2808
rect 82633 2805 82645 2808
rect 82679 2805 82691 2839
rect 82633 2799 82691 2805
rect 87046 2796 87052 2848
rect 87104 2836 87110 2848
rect 88794 2836 88800 2848
rect 87104 2808 88800 2836
rect 87104 2796 87110 2808
rect 88794 2796 88800 2808
rect 88852 2796 88858 2848
rect 90818 2796 90824 2848
rect 90876 2836 90882 2848
rect 91649 2839 91707 2845
rect 91649 2836 91661 2839
rect 90876 2808 91661 2836
rect 90876 2796 90882 2808
rect 91649 2805 91661 2808
rect 91695 2805 91707 2839
rect 91649 2799 91707 2805
rect 91922 2796 91928 2848
rect 91980 2836 91986 2848
rect 92385 2839 92443 2845
rect 92385 2836 92397 2839
rect 91980 2808 92397 2836
rect 91980 2796 91986 2808
rect 92385 2805 92397 2808
rect 92431 2805 92443 2839
rect 92385 2799 92443 2805
rect 92842 2796 92848 2848
rect 92900 2836 92906 2848
rect 92937 2839 92995 2845
rect 92937 2836 92949 2839
rect 92900 2808 92949 2836
rect 92900 2796 92906 2808
rect 92937 2805 92949 2808
rect 92983 2836 92995 2839
rect 93320 2836 93348 2867
rect 93394 2864 93400 2916
rect 93452 2904 93458 2916
rect 93854 2904 93860 2916
rect 93452 2876 93860 2904
rect 93452 2864 93458 2876
rect 93854 2864 93860 2876
rect 93912 2864 93918 2916
rect 94332 2904 94360 3012
rect 94406 2932 94412 2984
rect 94464 2972 94470 2984
rect 94792 2981 94820 3012
rect 96154 3000 96160 3052
rect 96212 3040 96218 3052
rect 96709 3043 96767 3049
rect 96709 3040 96721 3043
rect 96212 3012 96721 3040
rect 96212 3000 96218 3012
rect 96709 3009 96721 3012
rect 96755 3009 96767 3043
rect 97276 3040 97304 3139
rect 97276 3012 97672 3040
rect 96709 3003 96767 3009
rect 94593 2975 94651 2981
rect 94593 2972 94605 2975
rect 94464 2944 94605 2972
rect 94464 2932 94470 2944
rect 94593 2941 94605 2944
rect 94639 2941 94651 2975
rect 94593 2935 94651 2941
rect 94777 2975 94835 2981
rect 94777 2941 94789 2975
rect 94823 2941 94835 2975
rect 94777 2935 94835 2941
rect 95786 2932 95792 2984
rect 95844 2972 95850 2984
rect 95844 2944 96200 2972
rect 95844 2932 95850 2944
rect 94332 2876 95464 2904
rect 92983 2808 93348 2836
rect 92983 2805 92995 2808
rect 92937 2799 92995 2805
rect 93762 2796 93768 2848
rect 93820 2836 93826 2848
rect 94041 2839 94099 2845
rect 94041 2836 94053 2839
rect 93820 2808 94053 2836
rect 93820 2796 93826 2808
rect 94041 2805 94053 2808
rect 94087 2805 94099 2839
rect 94041 2799 94099 2805
rect 94590 2796 94596 2848
rect 94648 2836 94654 2848
rect 95326 2836 95332 2848
rect 94648 2808 95332 2836
rect 94648 2796 94654 2808
rect 95326 2796 95332 2808
rect 95384 2796 95390 2848
rect 95436 2836 95464 2876
rect 95602 2864 95608 2916
rect 95660 2904 95666 2916
rect 96172 2913 96200 2944
rect 96798 2932 96804 2984
rect 96856 2972 96862 2984
rect 97644 2981 97672 3012
rect 97718 3000 97724 3052
rect 97776 3040 97782 3052
rect 98822 3040 98828 3052
rect 97776 3012 98828 3040
rect 97776 3000 97782 3012
rect 98822 3000 98828 3012
rect 98880 3000 98886 3052
rect 97445 2975 97503 2981
rect 97445 2972 97457 2975
rect 96856 2944 97457 2972
rect 96856 2932 96862 2944
rect 97445 2941 97457 2944
rect 97491 2941 97503 2975
rect 97445 2935 97503 2941
rect 97629 2975 97687 2981
rect 97629 2941 97641 2975
rect 97675 2941 97687 2975
rect 97629 2935 97687 2941
rect 95973 2907 96031 2913
rect 95973 2904 95985 2907
rect 95660 2876 95985 2904
rect 95660 2864 95666 2876
rect 95973 2873 95985 2876
rect 96019 2873 96031 2907
rect 95973 2867 96031 2873
rect 96157 2907 96215 2913
rect 96157 2873 96169 2907
rect 96203 2873 96215 2907
rect 96157 2867 96215 2873
rect 96617 2907 96675 2913
rect 96617 2873 96629 2907
rect 96663 2904 96675 2907
rect 96890 2904 96896 2916
rect 96663 2876 96896 2904
rect 96663 2873 96675 2876
rect 96617 2867 96675 2873
rect 96890 2864 96896 2876
rect 96948 2864 96954 2916
rect 98362 2904 98368 2916
rect 97000 2876 98368 2904
rect 97000 2836 97028 2876
rect 98362 2864 98368 2876
rect 98420 2864 98426 2916
rect 95436 2808 97028 2836
rect 97718 2796 97724 2848
rect 97776 2836 97782 2848
rect 99834 2836 99840 2848
rect 97776 2808 99840 2836
rect 97776 2796 97782 2808
rect 99834 2796 99840 2808
rect 99892 2796 99898 2848
rect 1104 2746 98808 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 50326 2746
rect 50378 2694 50390 2746
rect 50442 2694 50454 2746
rect 50506 2694 50518 2746
rect 50570 2694 81046 2746
rect 81098 2694 81110 2746
rect 81162 2694 81174 2746
rect 81226 2694 81238 2746
rect 81290 2694 98808 2746
rect 1104 2672 98808 2694
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 11054 2632 11060 2644
rect 11015 2604 11060 2632
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 15289 2635 15347 2641
rect 13228 2604 13584 2632
rect 13228 2592 13234 2604
rect 7377 2567 7435 2573
rect 7377 2533 7389 2567
rect 7423 2564 7435 2567
rect 7650 2564 7656 2576
rect 7423 2536 7656 2564
rect 7423 2533 7435 2536
rect 7377 2527 7435 2533
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 10134 2564 10140 2576
rect 10095 2536 10140 2564
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 13354 2524 13360 2576
rect 13412 2564 13418 2576
rect 13449 2567 13507 2573
rect 13449 2564 13461 2567
rect 13412 2536 13461 2564
rect 13412 2524 13418 2536
rect 13449 2533 13461 2536
rect 13495 2533 13507 2567
rect 13556 2564 13584 2604
rect 15289 2601 15301 2635
rect 15335 2632 15347 2635
rect 15838 2632 15844 2644
rect 15335 2604 15844 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 15838 2592 15844 2604
rect 15896 2592 15902 2644
rect 16546 2604 28580 2632
rect 16546 2564 16574 2604
rect 13556 2536 16574 2564
rect 13449 2527 13507 2533
rect 17770 2524 17776 2576
rect 17828 2564 17834 2576
rect 17865 2567 17923 2573
rect 17865 2564 17877 2567
rect 17828 2536 17877 2564
rect 17828 2524 17834 2536
rect 17865 2533 17877 2536
rect 17911 2533 17923 2567
rect 17865 2527 17923 2533
rect 18785 2567 18843 2573
rect 18785 2533 18797 2567
rect 18831 2564 18843 2567
rect 18874 2564 18880 2576
rect 18831 2536 18880 2564
rect 18831 2533 18843 2536
rect 18785 2527 18843 2533
rect 18874 2524 18880 2536
rect 18932 2524 18938 2576
rect 20530 2564 20536 2576
rect 20491 2536 20536 2564
rect 20530 2524 20536 2536
rect 20588 2524 20594 2576
rect 21637 2567 21695 2573
rect 21637 2533 21649 2567
rect 21683 2564 21695 2567
rect 21726 2564 21732 2576
rect 21683 2536 21732 2564
rect 21683 2533 21695 2536
rect 21637 2527 21695 2533
rect 21726 2524 21732 2536
rect 21784 2524 21790 2576
rect 22833 2567 22891 2573
rect 22833 2533 22845 2567
rect 22879 2564 22891 2567
rect 23106 2564 23112 2576
rect 22879 2536 23112 2564
rect 22879 2533 22891 2536
rect 22833 2527 22891 2533
rect 23106 2524 23112 2536
rect 23164 2524 23170 2576
rect 23750 2564 23756 2576
rect 23711 2536 23756 2564
rect 23750 2524 23756 2536
rect 23808 2524 23814 2576
rect 25409 2567 25467 2573
rect 25409 2564 25421 2567
rect 23860 2536 25421 2564
rect 290 2456 296 2508
rect 348 2496 354 2508
rect 1765 2499 1823 2505
rect 1765 2496 1777 2499
rect 348 2468 1777 2496
rect 348 2456 354 2468
rect 1765 2465 1777 2468
rect 1811 2465 1823 2499
rect 1765 2459 1823 2465
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 4341 2499 4399 2505
rect 4341 2496 4353 2499
rect 3752 2468 4353 2496
rect 3752 2456 3758 2468
rect 4341 2465 4353 2468
rect 4387 2465 4399 2499
rect 4341 2459 4399 2465
rect 5166 2456 5172 2508
rect 5224 2496 5230 2508
rect 5537 2499 5595 2505
rect 5537 2496 5549 2499
rect 5224 2468 5549 2496
rect 5224 2456 5230 2468
rect 5537 2465 5549 2468
rect 5583 2465 5595 2499
rect 5537 2459 5595 2465
rect 5718 2456 5724 2508
rect 5776 2496 5782 2508
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 5776 2468 7021 2496
rect 5776 2456 5782 2468
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 8297 2499 8355 2505
rect 8297 2465 8309 2499
rect 8343 2496 8355 2499
rect 8386 2496 8392 2508
rect 8343 2468 8392 2496
rect 8343 2465 8355 2468
rect 8297 2459 8355 2465
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 9582 2456 9588 2508
rect 9640 2496 9646 2508
rect 9677 2499 9735 2505
rect 9677 2496 9689 2499
rect 9640 2468 9689 2496
rect 9640 2456 9646 2468
rect 9677 2465 9689 2468
rect 9723 2465 9735 2499
rect 10870 2496 10876 2508
rect 10831 2468 10876 2496
rect 9677 2459 9735 2465
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 11422 2456 11428 2508
rect 11480 2496 11486 2508
rect 12345 2499 12403 2505
rect 12345 2496 12357 2499
rect 11480 2468 12357 2496
rect 11480 2456 11486 2468
rect 12345 2465 12357 2468
rect 12391 2465 12403 2499
rect 12345 2459 12403 2465
rect 12618 2456 12624 2508
rect 12676 2496 12682 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12676 2468 13185 2496
rect 12676 2456 12682 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 15013 2499 15071 2505
rect 15013 2496 15025 2499
rect 14516 2468 15025 2496
rect 14516 2456 14522 2468
rect 15013 2465 15025 2468
rect 15059 2465 15071 2499
rect 15013 2459 15071 2465
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 15160 2468 15853 2496
rect 15160 2456 15166 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 16298 2456 16304 2508
rect 16356 2496 16362 2508
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 16356 2468 17601 2496
rect 16356 2456 16362 2468
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 17589 2459 17647 2465
rect 17678 2456 17684 2508
rect 17736 2496 17742 2508
rect 18509 2499 18567 2505
rect 18509 2496 18521 2499
rect 17736 2468 18521 2496
rect 17736 2456 17742 2468
rect 18509 2465 18521 2468
rect 18555 2465 18567 2499
rect 18509 2459 18567 2465
rect 19978 2456 19984 2508
rect 20036 2496 20042 2508
rect 20257 2499 20315 2505
rect 20257 2496 20269 2499
rect 20036 2468 20269 2496
rect 20036 2456 20042 2468
rect 20257 2465 20269 2468
rect 20303 2465 20315 2499
rect 20257 2459 20315 2465
rect 21174 2456 21180 2508
rect 21232 2496 21238 2508
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 21232 2468 21281 2496
rect 21232 2456 21238 2468
rect 21269 2465 21281 2468
rect 21315 2465 21327 2499
rect 23860 2496 23888 2536
rect 25409 2533 25421 2536
rect 25455 2564 25467 2567
rect 25777 2567 25835 2573
rect 25777 2564 25789 2567
rect 25455 2536 25789 2564
rect 25455 2533 25467 2536
rect 25409 2527 25467 2533
rect 25777 2533 25789 2536
rect 25823 2533 25835 2567
rect 25777 2527 25835 2533
rect 26970 2524 26976 2576
rect 27028 2564 27034 2576
rect 27065 2567 27123 2573
rect 27065 2564 27077 2567
rect 27028 2536 27077 2564
rect 27028 2524 27034 2536
rect 27065 2533 27077 2536
rect 27111 2533 27123 2567
rect 27065 2527 27123 2533
rect 28169 2567 28227 2573
rect 28169 2533 28181 2567
rect 28215 2564 28227 2567
rect 28442 2564 28448 2576
rect 28215 2536 28448 2564
rect 28215 2533 28227 2536
rect 28169 2527 28227 2533
rect 28442 2524 28448 2536
rect 28500 2524 28506 2576
rect 28552 2564 28580 2604
rect 28626 2592 28632 2644
rect 28684 2632 28690 2644
rect 33134 2632 33140 2644
rect 28684 2604 33140 2632
rect 28684 2592 28690 2604
rect 33134 2592 33140 2604
rect 33192 2592 33198 2644
rect 33410 2592 33416 2644
rect 33468 2632 33474 2644
rect 36357 2635 36415 2641
rect 36357 2632 36369 2635
rect 33468 2604 36369 2632
rect 33468 2592 33474 2604
rect 36357 2601 36369 2604
rect 36403 2601 36415 2635
rect 37921 2635 37979 2641
rect 37921 2632 37933 2635
rect 36357 2595 36415 2601
rect 36464 2604 37933 2632
rect 31018 2564 31024 2576
rect 28552 2536 29960 2564
rect 30979 2536 31024 2564
rect 21269 2459 21327 2465
rect 21744 2468 23888 2496
rect 24489 2499 24547 2505
rect 2590 2428 2596 2440
rect 2551 2400 2596 2428
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 11514 2428 11520 2440
rect 4939 2400 11520 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2428 16175 2431
rect 16206 2428 16212 2440
rect 16163 2400 16212 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 16206 2388 16212 2400
rect 16264 2388 16270 2440
rect 6086 2320 6092 2372
rect 6144 2360 6150 2372
rect 21266 2360 21272 2372
rect 6144 2332 21272 2360
rect 6144 2320 6150 2332
rect 21266 2320 21272 2332
rect 21324 2320 21330 2372
rect 5813 2295 5871 2301
rect 5813 2261 5825 2295
rect 5859 2292 5871 2295
rect 12158 2292 12164 2304
rect 5859 2264 12164 2292
rect 5859 2261 5871 2264
rect 5813 2255 5871 2261
rect 12158 2252 12164 2264
rect 12216 2252 12222 2304
rect 12621 2295 12679 2301
rect 12621 2261 12633 2295
rect 12667 2292 12679 2295
rect 13630 2292 13636 2304
rect 12667 2264 13636 2292
rect 12667 2261 12679 2264
rect 12621 2255 12679 2261
rect 13630 2252 13636 2264
rect 13688 2252 13694 2304
rect 15562 2252 15568 2304
rect 15620 2292 15626 2304
rect 21744 2292 21772 2468
rect 24489 2465 24501 2499
rect 24535 2496 24547 2499
rect 25314 2496 25320 2508
rect 24535 2468 25320 2496
rect 24535 2465 24547 2468
rect 24489 2459 24547 2465
rect 25314 2456 25320 2468
rect 25372 2456 25378 2508
rect 26234 2456 26240 2508
rect 26292 2496 26298 2508
rect 26513 2499 26571 2505
rect 26513 2496 26525 2499
rect 26292 2468 26525 2496
rect 26292 2456 26298 2468
rect 26513 2465 26525 2468
rect 26559 2465 26571 2499
rect 26513 2459 26571 2465
rect 26881 2499 26939 2505
rect 26881 2465 26893 2499
rect 26927 2496 26939 2499
rect 27246 2496 27252 2508
rect 26927 2468 27252 2496
rect 26927 2465 26939 2468
rect 26881 2459 26939 2465
rect 27246 2456 27252 2468
rect 27304 2456 27310 2508
rect 29089 2499 29147 2505
rect 29089 2465 29101 2499
rect 29135 2496 29147 2499
rect 29730 2496 29736 2508
rect 29135 2468 29736 2496
rect 29135 2465 29147 2468
rect 29089 2459 29147 2465
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 29825 2499 29883 2505
rect 29825 2465 29837 2499
rect 29871 2465 29883 2499
rect 29932 2496 29960 2536
rect 31018 2524 31024 2536
rect 31076 2524 31082 2576
rect 32490 2564 32496 2576
rect 31128 2536 31984 2564
rect 32451 2536 32496 2564
rect 31128 2496 31156 2536
rect 31754 2496 31760 2508
rect 29932 2468 31156 2496
rect 31715 2468 31760 2496
rect 29825 2459 29883 2465
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 23716 2400 25605 2428
rect 23716 2388 23722 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 28166 2388 28172 2440
rect 28224 2428 28230 2440
rect 29840 2428 29868 2459
rect 31754 2456 31760 2468
rect 31812 2456 31818 2508
rect 31956 2496 31984 2536
rect 32490 2524 32496 2536
rect 32548 2524 32554 2576
rect 33686 2564 33692 2576
rect 33647 2536 33692 2564
rect 33686 2524 33692 2536
rect 33744 2524 33750 2576
rect 34054 2524 34060 2576
rect 34112 2564 34118 2576
rect 34425 2567 34483 2573
rect 34425 2564 34437 2567
rect 34112 2536 34437 2564
rect 34112 2524 34118 2536
rect 34425 2533 34437 2536
rect 34471 2533 34483 2567
rect 34425 2527 34483 2533
rect 35161 2567 35219 2573
rect 35161 2533 35173 2567
rect 35207 2564 35219 2567
rect 35250 2564 35256 2576
rect 35207 2536 35256 2564
rect 35207 2533 35219 2536
rect 35161 2527 35219 2533
rect 35250 2524 35256 2536
rect 35308 2524 35314 2576
rect 35986 2524 35992 2576
rect 36044 2564 36050 2576
rect 36081 2567 36139 2573
rect 36081 2564 36093 2567
rect 36044 2536 36093 2564
rect 36044 2524 36050 2536
rect 36081 2533 36093 2536
rect 36127 2533 36139 2567
rect 36081 2527 36139 2533
rect 36096 2496 36124 2527
rect 36170 2524 36176 2576
rect 36228 2564 36234 2576
rect 36464 2564 36492 2604
rect 37921 2601 37933 2604
rect 37967 2601 37979 2635
rect 37921 2595 37979 2601
rect 38286 2592 38292 2644
rect 38344 2632 38350 2644
rect 41785 2635 41843 2641
rect 41785 2632 41797 2635
rect 38344 2604 41797 2632
rect 38344 2592 38350 2604
rect 41785 2601 41797 2604
rect 41831 2601 41843 2635
rect 43257 2635 43315 2641
rect 43257 2632 43269 2635
rect 41785 2595 41843 2601
rect 42260 2604 43269 2632
rect 37829 2567 37887 2573
rect 36228 2536 36492 2564
rect 36556 2536 37780 2564
rect 36228 2524 36234 2536
rect 36446 2496 36452 2508
rect 31956 2468 35894 2496
rect 36096 2468 36452 2496
rect 28224 2400 29868 2428
rect 28224 2388 28230 2400
rect 30926 2388 30932 2440
rect 30984 2428 30990 2440
rect 32677 2431 32735 2437
rect 32677 2428 32689 2431
rect 30984 2400 32689 2428
rect 30984 2388 30990 2400
rect 32677 2397 32689 2400
rect 32723 2397 32735 2431
rect 35866 2428 35894 2468
rect 36446 2456 36452 2468
rect 36504 2456 36510 2508
rect 36556 2428 36584 2536
rect 36906 2496 36912 2508
rect 36867 2468 36912 2496
rect 36906 2456 36912 2468
rect 36964 2496 36970 2508
rect 37185 2499 37243 2505
rect 37185 2496 37197 2499
rect 36964 2468 37197 2496
rect 36964 2456 36970 2468
rect 37185 2465 37197 2468
rect 37231 2465 37243 2499
rect 37752 2496 37780 2536
rect 37829 2533 37841 2567
rect 37875 2564 37887 2567
rect 38746 2564 38752 2576
rect 37875 2536 38752 2564
rect 37875 2533 37887 2536
rect 37829 2527 37887 2533
rect 38746 2524 38752 2536
rect 38804 2524 38810 2576
rect 38841 2567 38899 2573
rect 38841 2533 38853 2567
rect 38887 2564 38899 2567
rect 39114 2564 39120 2576
rect 38887 2536 39120 2564
rect 38887 2533 38899 2536
rect 38841 2527 38899 2533
rect 39114 2524 39120 2536
rect 39172 2524 39178 2576
rect 39577 2567 39635 2573
rect 39577 2533 39589 2567
rect 39623 2564 39635 2567
rect 39850 2564 39856 2576
rect 39623 2536 39856 2564
rect 39623 2533 39635 2536
rect 39577 2527 39635 2533
rect 39850 2524 39856 2536
rect 39908 2524 39914 2576
rect 40313 2567 40371 2573
rect 40313 2533 40325 2567
rect 40359 2564 40371 2567
rect 40586 2564 40592 2576
rect 40359 2536 40592 2564
rect 40359 2533 40371 2536
rect 40313 2527 40371 2533
rect 40586 2524 40592 2536
rect 40644 2564 40650 2576
rect 40773 2567 40831 2573
rect 40773 2564 40785 2567
rect 40644 2536 40785 2564
rect 40644 2524 40650 2536
rect 40773 2533 40785 2536
rect 40819 2533 40831 2567
rect 42260 2564 42288 2604
rect 43257 2601 43269 2604
rect 43303 2601 43315 2635
rect 43257 2595 43315 2601
rect 44726 2592 44732 2644
rect 44784 2632 44790 2644
rect 44821 2635 44879 2641
rect 44821 2632 44833 2635
rect 44784 2604 44833 2632
rect 44784 2592 44790 2604
rect 44821 2601 44833 2604
rect 44867 2632 44879 2635
rect 44867 2604 45232 2632
rect 44867 2601 44879 2604
rect 44821 2595 44879 2601
rect 42426 2564 42432 2576
rect 40773 2527 40831 2533
rect 40880 2536 42288 2564
rect 42387 2536 42432 2564
rect 39390 2496 39396 2508
rect 37752 2468 39396 2496
rect 37185 2459 37243 2465
rect 39390 2456 39396 2468
rect 39448 2456 39454 2508
rect 39482 2456 39488 2508
rect 39540 2496 39546 2508
rect 40880 2496 40908 2536
rect 42426 2524 42432 2536
rect 42484 2524 42490 2576
rect 43165 2567 43223 2573
rect 43165 2533 43177 2567
rect 43211 2564 43223 2567
rect 44082 2564 44088 2576
rect 43211 2536 44088 2564
rect 43211 2533 43223 2536
rect 43165 2527 43223 2533
rect 44082 2524 44088 2536
rect 44140 2524 44146 2576
rect 44177 2567 44235 2573
rect 44177 2533 44189 2567
rect 44223 2564 44235 2567
rect 44450 2564 44456 2576
rect 44223 2536 44456 2564
rect 44223 2533 44235 2536
rect 44177 2527 44235 2533
rect 44450 2524 44456 2536
rect 44508 2524 44514 2576
rect 45204 2573 45232 2604
rect 46106 2592 46112 2644
rect 46164 2632 46170 2644
rect 47857 2635 47915 2641
rect 47857 2632 47869 2635
rect 46164 2604 47869 2632
rect 46164 2592 46170 2604
rect 47857 2601 47869 2604
rect 47903 2601 47915 2635
rect 48314 2632 48320 2644
rect 48275 2604 48320 2632
rect 47857 2595 47915 2601
rect 48314 2592 48320 2604
rect 48372 2632 48378 2644
rect 48372 2604 48636 2632
rect 48372 2592 48378 2604
rect 45189 2567 45247 2573
rect 45189 2533 45201 2567
rect 45235 2533 45247 2567
rect 45189 2527 45247 2533
rect 45833 2567 45891 2573
rect 45833 2533 45845 2567
rect 45879 2564 45891 2567
rect 46750 2564 46756 2576
rect 45879 2536 46756 2564
rect 45879 2533 45891 2536
rect 45833 2527 45891 2533
rect 46750 2524 46756 2536
rect 46808 2524 46814 2576
rect 47762 2564 47768 2576
rect 47723 2536 47768 2564
rect 47762 2524 47768 2536
rect 47820 2524 47826 2576
rect 48608 2573 48636 2604
rect 49786 2592 49792 2644
rect 49844 2632 49850 2644
rect 49881 2635 49939 2641
rect 49881 2632 49893 2635
rect 49844 2604 49893 2632
rect 49844 2592 49850 2604
rect 49881 2601 49893 2604
rect 49927 2601 49939 2635
rect 49881 2595 49939 2601
rect 49970 2592 49976 2644
rect 50028 2632 50034 2644
rect 53193 2635 53251 2641
rect 53193 2632 53205 2635
rect 50028 2604 53205 2632
rect 50028 2592 50034 2604
rect 53193 2601 53205 2604
rect 53239 2601 53251 2635
rect 53193 2595 53251 2601
rect 54018 2592 54024 2644
rect 54076 2632 54082 2644
rect 56597 2635 56655 2641
rect 56597 2632 56609 2635
rect 54076 2604 56609 2632
rect 54076 2592 54082 2604
rect 56597 2601 56609 2604
rect 56643 2601 56655 2635
rect 56597 2595 56655 2601
rect 57330 2592 57336 2644
rect 57388 2632 57394 2644
rect 57425 2635 57483 2641
rect 57425 2632 57437 2635
rect 57388 2604 57437 2632
rect 57388 2592 57394 2604
rect 57425 2601 57437 2604
rect 57471 2632 57483 2635
rect 57471 2604 57836 2632
rect 57471 2601 57483 2604
rect 57425 2595 57483 2601
rect 48593 2567 48651 2573
rect 48593 2533 48605 2567
rect 48639 2564 48651 2567
rect 48777 2567 48835 2573
rect 48777 2564 48789 2567
rect 48639 2536 48789 2564
rect 48639 2533 48651 2536
rect 48593 2527 48651 2533
rect 48777 2533 48789 2536
rect 48823 2533 48835 2567
rect 51534 2564 51540 2576
rect 48777 2527 48835 2533
rect 50356 2536 51540 2564
rect 39540 2468 40908 2496
rect 41693 2499 41751 2505
rect 39540 2456 39546 2468
rect 41693 2465 41705 2499
rect 41739 2496 41751 2499
rect 42242 2496 42248 2508
rect 41739 2468 42248 2496
rect 41739 2465 41751 2468
rect 41693 2459 41751 2465
rect 42242 2456 42248 2468
rect 42300 2456 42306 2508
rect 42518 2456 42524 2508
rect 42576 2496 42582 2508
rect 46017 2499 46075 2505
rect 46017 2496 46029 2499
rect 42576 2468 46029 2496
rect 42576 2456 42582 2468
rect 46017 2465 46029 2468
rect 46063 2465 46075 2499
rect 46017 2459 46075 2465
rect 47029 2499 47087 2505
rect 47029 2465 47041 2499
rect 47075 2496 47087 2499
rect 47670 2496 47676 2508
rect 47075 2468 47676 2496
rect 47075 2465 47087 2468
rect 47029 2459 47087 2465
rect 47670 2456 47676 2468
rect 47728 2456 47734 2508
rect 49878 2456 49884 2508
rect 49936 2496 49942 2508
rect 50356 2505 50384 2536
rect 51534 2524 51540 2536
rect 51592 2524 51598 2576
rect 52362 2564 52368 2576
rect 52323 2536 52368 2564
rect 52362 2524 52368 2536
rect 52420 2524 52426 2576
rect 53101 2567 53159 2573
rect 53101 2533 53113 2567
rect 53147 2564 53159 2567
rect 53742 2564 53748 2576
rect 53147 2536 53748 2564
rect 53147 2533 53159 2536
rect 53101 2527 53159 2533
rect 53742 2524 53748 2536
rect 53800 2524 53806 2576
rect 53837 2567 53895 2573
rect 53837 2533 53849 2567
rect 53883 2564 53895 2567
rect 54110 2564 54116 2576
rect 53883 2536 54116 2564
rect 53883 2533 53895 2536
rect 53837 2527 53895 2533
rect 54110 2524 54116 2536
rect 54168 2524 54174 2576
rect 55030 2564 55036 2576
rect 54991 2536 55036 2564
rect 55030 2524 55036 2536
rect 55088 2524 55094 2576
rect 55398 2524 55404 2576
rect 55456 2564 55462 2576
rect 55769 2567 55827 2573
rect 55769 2564 55781 2567
rect 55456 2536 55781 2564
rect 55456 2524 55462 2536
rect 55769 2533 55781 2536
rect 55815 2533 55827 2567
rect 55769 2527 55827 2533
rect 55953 2567 56011 2573
rect 55953 2533 55965 2567
rect 55999 2533 56011 2567
rect 55953 2527 56011 2533
rect 50065 2499 50123 2505
rect 50065 2496 50077 2499
rect 49936 2468 50077 2496
rect 49936 2456 49942 2468
rect 50065 2465 50077 2468
rect 50111 2465 50123 2499
rect 50249 2499 50307 2505
rect 50249 2496 50261 2499
rect 50065 2459 50123 2465
rect 50172 2468 50261 2496
rect 35866 2400 36584 2428
rect 32677 2391 32735 2397
rect 37918 2388 37924 2440
rect 37976 2428 37982 2440
rect 39669 2431 39727 2437
rect 39669 2428 39681 2431
rect 37976 2400 39681 2428
rect 37976 2388 37982 2400
rect 39669 2397 39681 2400
rect 39715 2397 39727 2431
rect 39669 2391 39727 2397
rect 40678 2388 40684 2440
rect 40736 2428 40742 2440
rect 44269 2431 44327 2437
rect 44269 2428 44281 2431
rect 40736 2400 44281 2428
rect 40736 2388 40742 2400
rect 44269 2397 44281 2400
rect 44315 2397 44327 2431
rect 44269 2391 44327 2397
rect 45002 2388 45008 2440
rect 45060 2428 45066 2440
rect 48409 2431 48467 2437
rect 48409 2428 48421 2431
rect 45060 2400 48421 2428
rect 45060 2388 45066 2400
rect 48409 2397 48421 2400
rect 48455 2397 48467 2431
rect 48409 2391 48467 2397
rect 21818 2320 21824 2372
rect 21876 2360 21882 2372
rect 22925 2363 22983 2369
rect 22925 2360 22937 2363
rect 21876 2332 22937 2360
rect 21876 2320 21882 2332
rect 22925 2329 22937 2332
rect 22971 2329 22983 2363
rect 22925 2323 22983 2329
rect 23014 2320 23020 2372
rect 23072 2360 23078 2372
rect 24673 2363 24731 2369
rect 24673 2360 24685 2363
rect 23072 2332 24685 2360
rect 23072 2320 23078 2332
rect 24673 2329 24685 2332
rect 24719 2329 24731 2363
rect 26329 2363 26387 2369
rect 26329 2360 26341 2363
rect 24673 2323 24731 2329
rect 24872 2332 26341 2360
rect 15620 2264 21772 2292
rect 15620 2252 15626 2264
rect 22462 2252 22468 2304
rect 22520 2292 22526 2304
rect 23845 2295 23903 2301
rect 23845 2292 23857 2295
rect 22520 2264 23857 2292
rect 22520 2252 22526 2264
rect 23845 2261 23857 2264
rect 23891 2261 23903 2295
rect 23845 2255 23903 2261
rect 24210 2252 24216 2304
rect 24268 2292 24274 2304
rect 24872 2292 24900 2332
rect 26329 2329 26341 2332
rect 26375 2329 26387 2363
rect 26329 2323 26387 2329
rect 27890 2320 27896 2372
rect 27948 2360 27954 2372
rect 28261 2363 28319 2369
rect 28261 2360 28273 2363
rect 27948 2332 28273 2360
rect 27948 2320 27954 2332
rect 28261 2329 28273 2332
rect 28307 2329 28319 2363
rect 28261 2323 28319 2329
rect 29086 2320 29092 2372
rect 29144 2360 29150 2372
rect 30009 2363 30067 2369
rect 30009 2360 30021 2363
rect 29144 2332 30021 2360
rect 29144 2320 29150 2332
rect 30009 2329 30021 2332
rect 30055 2329 30067 2363
rect 30009 2323 30067 2329
rect 30374 2320 30380 2372
rect 30432 2360 30438 2372
rect 31941 2363 31999 2369
rect 31941 2360 31953 2363
rect 30432 2332 31953 2360
rect 30432 2320 30438 2332
rect 31941 2329 31953 2332
rect 31987 2329 31999 2363
rect 31941 2323 31999 2329
rect 32214 2320 32220 2372
rect 32272 2360 32278 2372
rect 34609 2363 34667 2369
rect 34609 2360 34621 2363
rect 32272 2332 34621 2360
rect 32272 2320 32278 2332
rect 34609 2329 34621 2332
rect 34655 2329 34667 2363
rect 34609 2323 34667 2329
rect 34698 2320 34704 2372
rect 34756 2360 34762 2372
rect 37001 2363 37059 2369
rect 37001 2360 37013 2363
rect 34756 2332 37013 2360
rect 34756 2320 34762 2332
rect 37001 2329 37013 2332
rect 37047 2329 37059 2363
rect 37001 2323 37059 2329
rect 37182 2320 37188 2372
rect 37240 2360 37246 2372
rect 38933 2363 38991 2369
rect 38933 2360 38945 2363
rect 37240 2332 38945 2360
rect 37240 2320 37246 2332
rect 38933 2329 38945 2332
rect 38979 2329 38991 2363
rect 38933 2323 38991 2329
rect 39022 2320 39028 2372
rect 39080 2360 39086 2372
rect 42613 2363 42671 2369
rect 42613 2360 42625 2363
rect 39080 2332 40724 2360
rect 39080 2320 39086 2332
rect 24268 2264 24900 2292
rect 24268 2252 24274 2264
rect 28534 2252 28540 2304
rect 28592 2292 28598 2304
rect 29181 2295 29239 2301
rect 29181 2292 29193 2295
rect 28592 2264 29193 2292
rect 28592 2252 28598 2264
rect 29181 2261 29193 2264
rect 29227 2261 29239 2295
rect 29181 2255 29239 2261
rect 29730 2252 29736 2304
rect 29788 2292 29794 2304
rect 31113 2295 31171 2301
rect 31113 2292 31125 2295
rect 29788 2264 31125 2292
rect 29788 2252 29794 2264
rect 31113 2261 31125 2264
rect 31159 2261 31171 2295
rect 31113 2255 31171 2261
rect 31570 2252 31576 2304
rect 31628 2292 31634 2304
rect 33781 2295 33839 2301
rect 33781 2292 33793 2295
rect 31628 2264 33793 2292
rect 31628 2252 31634 2264
rect 33781 2261 33793 2264
rect 33827 2261 33839 2295
rect 33781 2255 33839 2261
rect 33962 2252 33968 2304
rect 34020 2292 34026 2304
rect 35253 2295 35311 2301
rect 35253 2292 35265 2295
rect 34020 2264 35265 2292
rect 34020 2252 34026 2264
rect 35253 2261 35265 2264
rect 35299 2261 35311 2295
rect 35253 2255 35311 2261
rect 36446 2252 36452 2304
rect 36504 2292 36510 2304
rect 36633 2295 36691 2301
rect 36633 2292 36645 2295
rect 36504 2264 36645 2292
rect 36504 2252 36510 2264
rect 36633 2261 36645 2264
rect 36679 2261 36691 2295
rect 36633 2255 36691 2261
rect 37090 2252 37096 2304
rect 37148 2292 37154 2304
rect 40497 2295 40555 2301
rect 40497 2292 40509 2295
rect 37148 2264 40509 2292
rect 37148 2252 37154 2264
rect 40497 2261 40509 2264
rect 40543 2261 40555 2295
rect 40696 2292 40724 2332
rect 41386 2332 42625 2360
rect 41386 2292 41414 2332
rect 42613 2329 42625 2332
rect 42659 2329 42671 2363
rect 42613 2323 42671 2329
rect 43806 2320 43812 2372
rect 43864 2360 43870 2372
rect 47213 2363 47271 2369
rect 47213 2360 47225 2363
rect 43864 2332 47225 2360
rect 43864 2320 43870 2332
rect 47213 2329 47225 2332
rect 47259 2329 47271 2363
rect 50172 2360 50200 2468
rect 50249 2465 50261 2468
rect 50295 2465 50307 2499
rect 50249 2459 50307 2465
rect 50341 2499 50399 2505
rect 50341 2465 50353 2499
rect 50387 2465 50399 2499
rect 50341 2459 50399 2465
rect 50893 2499 50951 2505
rect 50893 2465 50905 2499
rect 50939 2496 50951 2499
rect 51626 2496 51632 2508
rect 50939 2468 51632 2496
rect 50939 2465 50951 2468
rect 50893 2459 50951 2465
rect 51626 2456 51632 2468
rect 51684 2456 51690 2508
rect 52454 2456 52460 2508
rect 52512 2496 52518 2508
rect 55968 2496 55996 2527
rect 56134 2524 56140 2576
rect 56192 2564 56198 2576
rect 57808 2573 57836 2604
rect 60274 2592 60280 2644
rect 60332 2632 60338 2644
rect 61105 2635 61163 2641
rect 61105 2632 61117 2635
rect 60332 2604 61117 2632
rect 60332 2592 60338 2604
rect 61105 2601 61117 2604
rect 61151 2601 61163 2635
rect 61105 2595 61163 2601
rect 61378 2592 61384 2644
rect 61436 2632 61442 2644
rect 61565 2635 61623 2641
rect 61565 2632 61577 2635
rect 61436 2604 61577 2632
rect 61436 2592 61442 2604
rect 61565 2601 61577 2604
rect 61611 2601 61623 2635
rect 61565 2595 61623 2601
rect 62114 2592 62120 2644
rect 62172 2632 62178 2644
rect 64601 2635 64659 2641
rect 64601 2632 64613 2635
rect 62172 2604 64613 2632
rect 62172 2592 62178 2604
rect 64601 2601 64613 2604
rect 64647 2601 64659 2635
rect 66622 2632 66628 2644
rect 64601 2595 64659 2601
rect 66548 2604 66628 2632
rect 56505 2567 56563 2573
rect 56505 2564 56517 2567
rect 56192 2536 56517 2564
rect 56192 2524 56198 2536
rect 56505 2533 56517 2536
rect 56551 2533 56563 2567
rect 56505 2527 56563 2533
rect 57793 2567 57851 2573
rect 57793 2533 57805 2567
rect 57839 2533 57851 2567
rect 58342 2564 58348 2576
rect 58303 2536 58348 2564
rect 57793 2527 57851 2533
rect 58342 2524 58348 2536
rect 58400 2524 58406 2576
rect 59170 2564 59176 2576
rect 59131 2536 59176 2564
rect 59170 2524 59176 2536
rect 59228 2524 59234 2576
rect 60185 2567 60243 2573
rect 60185 2533 60197 2567
rect 60231 2564 60243 2567
rect 60458 2564 60464 2576
rect 60231 2536 60464 2564
rect 60231 2533 60243 2536
rect 60185 2527 60243 2533
rect 60458 2524 60464 2536
rect 60516 2524 60522 2576
rect 60734 2524 60740 2576
rect 60792 2564 60798 2576
rect 62853 2567 62911 2573
rect 60792 2536 62068 2564
rect 60792 2524 60798 2536
rect 52512 2468 55996 2496
rect 52512 2456 52518 2468
rect 58066 2456 58072 2508
rect 58124 2496 58130 2508
rect 58529 2499 58587 2505
rect 58529 2496 58541 2499
rect 58124 2468 58541 2496
rect 58124 2456 58130 2468
rect 58529 2465 58541 2468
rect 58575 2465 58587 2499
rect 58529 2459 58587 2465
rect 60921 2499 60979 2505
rect 60921 2465 60933 2499
rect 60967 2496 60979 2499
rect 61194 2496 61200 2508
rect 60967 2468 61200 2496
rect 60967 2465 60979 2468
rect 60921 2459 60979 2465
rect 61194 2456 61200 2468
rect 61252 2456 61258 2508
rect 61378 2456 61384 2508
rect 61436 2496 61442 2508
rect 61933 2499 61991 2505
rect 61933 2496 61945 2499
rect 61436 2468 61945 2496
rect 61436 2456 61442 2468
rect 61933 2465 61945 2468
rect 61979 2465 61991 2499
rect 62040 2496 62068 2536
rect 62853 2533 62865 2567
rect 62899 2564 62911 2567
rect 63126 2564 63132 2576
rect 62899 2536 63132 2564
rect 62899 2533 62911 2536
rect 62853 2527 62911 2533
rect 63126 2524 63132 2536
rect 63184 2524 63190 2576
rect 63770 2564 63776 2576
rect 63731 2536 63776 2564
rect 63770 2524 63776 2536
rect 63828 2524 63834 2576
rect 63862 2524 63868 2576
rect 63920 2564 63926 2576
rect 63920 2536 64874 2564
rect 63920 2524 63926 2536
rect 62945 2499 63003 2505
rect 62945 2496 62957 2499
rect 62040 2468 62957 2496
rect 61933 2459 61991 2465
rect 62945 2465 62957 2468
rect 62991 2465 63003 2499
rect 62945 2459 63003 2465
rect 64414 2456 64420 2508
rect 64472 2496 64478 2508
rect 64509 2499 64567 2505
rect 64509 2496 64521 2499
rect 64472 2468 64521 2496
rect 64472 2456 64478 2468
rect 64509 2465 64521 2468
rect 64555 2465 64567 2499
rect 64846 2496 64874 2536
rect 65426 2524 65432 2576
rect 65484 2564 65490 2576
rect 66548 2573 66576 2604
rect 66622 2592 66628 2604
rect 66680 2632 66686 2644
rect 66717 2635 66775 2641
rect 66717 2632 66729 2635
rect 66680 2604 66729 2632
rect 66680 2592 66686 2604
rect 66717 2601 66729 2604
rect 66763 2601 66775 2635
rect 66990 2632 66996 2644
rect 66951 2604 66996 2632
rect 66717 2595 66775 2601
rect 66990 2592 66996 2604
rect 67048 2632 67054 2644
rect 68094 2632 68100 2644
rect 67048 2604 67312 2632
rect 68055 2604 68100 2632
rect 67048 2592 67054 2604
rect 67284 2573 67312 2604
rect 68094 2592 68100 2604
rect 68152 2632 68158 2644
rect 68830 2632 68836 2644
rect 68152 2604 68508 2632
rect 68791 2604 68836 2632
rect 68152 2592 68158 2604
rect 68480 2573 68508 2604
rect 68830 2592 68836 2604
rect 68888 2632 68894 2644
rect 68888 2604 69244 2632
rect 68888 2592 68894 2604
rect 69216 2573 69244 2604
rect 71682 2592 71688 2644
rect 71740 2632 71746 2644
rect 74166 2632 74172 2644
rect 71740 2604 73752 2632
rect 74127 2604 74172 2632
rect 71740 2592 71746 2604
rect 65705 2567 65763 2573
rect 65705 2564 65717 2567
rect 65484 2536 65717 2564
rect 65484 2524 65490 2536
rect 65705 2533 65717 2536
rect 65751 2533 65763 2567
rect 65705 2527 65763 2533
rect 66257 2567 66315 2573
rect 66257 2533 66269 2567
rect 66303 2564 66315 2567
rect 66533 2567 66591 2573
rect 66533 2564 66545 2567
rect 66303 2536 66545 2564
rect 66303 2533 66315 2536
rect 66257 2527 66315 2533
rect 66533 2533 66545 2536
rect 66579 2533 66591 2567
rect 66533 2527 66591 2533
rect 67269 2567 67327 2573
rect 67269 2533 67281 2567
rect 67315 2564 67327 2567
rect 67453 2567 67511 2573
rect 67453 2564 67465 2567
rect 67315 2536 67465 2564
rect 67315 2533 67327 2536
rect 67269 2527 67327 2533
rect 67453 2533 67465 2536
rect 67499 2533 67511 2567
rect 67453 2527 67511 2533
rect 68465 2567 68523 2573
rect 68465 2533 68477 2567
rect 68511 2533 68523 2567
rect 68465 2527 68523 2533
rect 69201 2567 69259 2573
rect 69201 2533 69213 2567
rect 69247 2533 69259 2567
rect 69201 2527 69259 2533
rect 69845 2567 69903 2573
rect 69845 2533 69857 2567
rect 69891 2564 69903 2567
rect 70302 2564 70308 2576
rect 69891 2536 70308 2564
rect 69891 2533 69903 2536
rect 69845 2527 69903 2533
rect 70302 2524 70308 2536
rect 70360 2524 70366 2576
rect 71041 2567 71099 2573
rect 71041 2533 71053 2567
rect 71087 2564 71099 2567
rect 71222 2564 71228 2576
rect 71087 2536 71228 2564
rect 71087 2533 71099 2536
rect 71041 2527 71099 2533
rect 71222 2524 71228 2536
rect 71280 2524 71286 2576
rect 73724 2573 73752 2604
rect 74166 2592 74172 2604
rect 74224 2632 74230 2644
rect 74224 2604 74580 2632
rect 74224 2592 74230 2604
rect 74552 2573 74580 2604
rect 74718 2592 74724 2644
rect 74776 2632 74782 2644
rect 77941 2635 77999 2641
rect 77941 2632 77953 2635
rect 74776 2604 77953 2632
rect 74776 2592 74782 2604
rect 77941 2601 77953 2604
rect 77987 2601 77999 2635
rect 79502 2632 79508 2644
rect 79463 2604 79508 2632
rect 77941 2595 77999 2601
rect 79502 2592 79508 2604
rect 79560 2632 79566 2644
rect 80238 2632 80244 2644
rect 79560 2604 79916 2632
rect 80199 2604 80244 2632
rect 79560 2592 79566 2604
rect 71961 2567 72019 2573
rect 71961 2564 71973 2567
rect 71332 2536 71973 2564
rect 67085 2499 67143 2505
rect 67085 2496 67097 2499
rect 64846 2468 67097 2496
rect 64509 2459 64567 2465
rect 67085 2465 67097 2468
rect 67131 2465 67143 2499
rect 67085 2459 67143 2465
rect 69290 2456 69296 2508
rect 69348 2496 69354 2508
rect 71332 2496 71360 2536
rect 71961 2533 71973 2536
rect 72007 2533 72019 2567
rect 73709 2567 73767 2573
rect 71961 2527 72019 2533
rect 72068 2536 73200 2564
rect 71774 2496 71780 2508
rect 69348 2468 71360 2496
rect 71735 2468 71780 2496
rect 69348 2456 69354 2468
rect 71774 2456 71780 2468
rect 71832 2456 71838 2508
rect 71866 2456 71872 2508
rect 71924 2496 71930 2508
rect 72068 2496 72096 2536
rect 71924 2468 72096 2496
rect 71924 2456 71930 2468
rect 72142 2456 72148 2508
rect 72200 2496 72206 2508
rect 72605 2499 72663 2505
rect 72605 2496 72617 2499
rect 72200 2468 72617 2496
rect 72200 2456 72206 2468
rect 72605 2465 72617 2468
rect 72651 2465 72663 2499
rect 73172 2496 73200 2536
rect 73709 2533 73721 2567
rect 73755 2533 73767 2567
rect 73709 2527 73767 2533
rect 74537 2567 74595 2573
rect 74537 2533 74549 2567
rect 74583 2533 74595 2567
rect 74537 2527 74595 2533
rect 74997 2567 75055 2573
rect 74997 2533 75009 2567
rect 75043 2564 75055 2567
rect 75273 2567 75331 2573
rect 75273 2564 75285 2567
rect 75043 2536 75285 2564
rect 75043 2533 75055 2536
rect 74997 2527 75055 2533
rect 75273 2533 75285 2536
rect 75319 2564 75331 2567
rect 75362 2564 75368 2576
rect 75319 2536 75368 2564
rect 75319 2533 75331 2536
rect 75273 2527 75331 2533
rect 75362 2524 75368 2536
rect 75420 2524 75426 2576
rect 76098 2524 76104 2576
rect 76156 2564 76162 2576
rect 77846 2564 77852 2576
rect 76156 2536 77432 2564
rect 77807 2536 77852 2564
rect 76156 2524 76162 2536
rect 75089 2499 75147 2505
rect 75089 2496 75101 2499
rect 73172 2468 75101 2496
rect 72605 2459 72663 2465
rect 75089 2465 75101 2468
rect 75135 2465 75147 2499
rect 76374 2496 76380 2508
rect 76335 2468 76380 2496
rect 75089 2459 75147 2465
rect 76374 2456 76380 2468
rect 76432 2456 76438 2508
rect 76558 2456 76564 2508
rect 76616 2496 76622 2508
rect 77113 2499 77171 2505
rect 77113 2496 77125 2499
rect 76616 2468 77125 2496
rect 76616 2456 76622 2468
rect 77113 2465 77125 2468
rect 77159 2465 77171 2499
rect 77404 2496 77432 2536
rect 77846 2524 77852 2536
rect 77904 2524 77910 2576
rect 79888 2573 79916 2604
rect 80238 2592 80244 2604
rect 80296 2632 80302 2644
rect 85758 2632 85764 2644
rect 80296 2604 80652 2632
rect 85719 2604 85764 2632
rect 80296 2592 80302 2604
rect 80624 2573 80652 2604
rect 85758 2592 85764 2604
rect 85816 2592 85822 2644
rect 86402 2592 86408 2644
rect 86460 2632 86466 2644
rect 86460 2604 87920 2632
rect 86460 2592 86466 2604
rect 79873 2567 79931 2573
rect 79873 2533 79885 2567
rect 79919 2533 79931 2567
rect 79873 2527 79931 2533
rect 80609 2567 80667 2573
rect 80609 2533 80621 2567
rect 80655 2533 80667 2567
rect 80609 2527 80667 2533
rect 81989 2567 82047 2573
rect 81989 2533 82001 2567
rect 82035 2564 82047 2567
rect 82173 2567 82231 2573
rect 82173 2564 82185 2567
rect 82035 2536 82185 2564
rect 82035 2533 82047 2536
rect 81989 2527 82047 2533
rect 82173 2533 82185 2536
rect 82219 2564 82231 2567
rect 82446 2564 82452 2576
rect 82219 2536 82452 2564
rect 82219 2533 82231 2536
rect 82173 2527 82231 2533
rect 82446 2524 82452 2536
rect 82504 2524 82510 2576
rect 82725 2567 82783 2573
rect 82725 2533 82737 2567
rect 82771 2564 82783 2567
rect 83001 2567 83059 2573
rect 83001 2564 83013 2567
rect 82771 2536 83013 2564
rect 82771 2533 82783 2536
rect 82725 2527 82783 2533
rect 83001 2533 83013 2536
rect 83047 2564 83059 2567
rect 83090 2564 83096 2576
rect 83047 2536 83096 2564
rect 83047 2533 83059 2536
rect 83001 2527 83059 2533
rect 83090 2524 83096 2536
rect 83148 2524 83154 2576
rect 86954 2524 86960 2576
rect 87012 2564 87018 2576
rect 87049 2567 87107 2573
rect 87049 2564 87061 2567
rect 87012 2536 87061 2564
rect 87012 2524 87018 2536
rect 87049 2533 87061 2536
rect 87095 2533 87107 2567
rect 87782 2564 87788 2576
rect 87743 2536 87788 2564
rect 87049 2527 87107 2533
rect 87782 2524 87788 2536
rect 87840 2524 87846 2576
rect 87892 2564 87920 2604
rect 88886 2592 88892 2644
rect 88944 2632 88950 2644
rect 89441 2635 89499 2641
rect 89441 2632 89453 2635
rect 88944 2604 89453 2632
rect 88944 2592 88950 2604
rect 89441 2601 89453 2604
rect 89487 2632 89499 2635
rect 90174 2632 90180 2644
rect 89487 2604 89852 2632
rect 90135 2604 90180 2632
rect 89487 2601 89499 2604
rect 89441 2595 89499 2601
rect 89824 2573 89852 2604
rect 90174 2592 90180 2604
rect 90232 2632 90238 2644
rect 90910 2632 90916 2644
rect 90232 2604 90588 2632
rect 90871 2604 90916 2632
rect 90232 2592 90238 2604
rect 90560 2573 90588 2604
rect 90910 2592 90916 2604
rect 90968 2632 90974 2644
rect 92106 2632 92112 2644
rect 90968 2604 91324 2632
rect 92067 2604 92112 2632
rect 90968 2592 90974 2604
rect 91296 2573 91324 2604
rect 92106 2592 92112 2604
rect 92164 2632 92170 2644
rect 92164 2604 92520 2632
rect 92164 2592 92170 2604
rect 92492 2573 92520 2604
rect 94498 2592 94504 2644
rect 94556 2632 94562 2644
rect 94777 2635 94835 2641
rect 94777 2632 94789 2635
rect 94556 2604 94789 2632
rect 94556 2592 94562 2604
rect 94777 2601 94789 2604
rect 94823 2632 94835 2635
rect 94823 2604 95188 2632
rect 94823 2601 94835 2604
rect 94777 2595 94835 2601
rect 89625 2567 89683 2573
rect 89625 2564 89637 2567
rect 87892 2536 89637 2564
rect 89625 2533 89637 2536
rect 89671 2533 89683 2567
rect 89625 2527 89683 2533
rect 89809 2567 89867 2573
rect 89809 2533 89821 2567
rect 89855 2533 89867 2567
rect 89809 2527 89867 2533
rect 90545 2567 90603 2573
rect 90545 2533 90557 2567
rect 90591 2533 90603 2567
rect 90545 2527 90603 2533
rect 91281 2567 91339 2573
rect 91281 2533 91293 2567
rect 91327 2533 91339 2567
rect 91281 2527 91339 2533
rect 92477 2567 92535 2573
rect 92477 2533 92489 2567
rect 92523 2533 92535 2567
rect 92477 2527 92535 2533
rect 93840 2567 93898 2573
rect 93840 2533 93852 2567
rect 93886 2564 93898 2567
rect 94038 2564 94044 2576
rect 93886 2536 94044 2564
rect 93886 2533 93898 2536
rect 93840 2527 93898 2533
rect 94038 2524 94044 2536
rect 94096 2524 94102 2576
rect 95160 2573 95188 2604
rect 95145 2567 95203 2573
rect 95145 2533 95157 2567
rect 95191 2533 95203 2567
rect 95145 2527 95203 2533
rect 96709 2567 96767 2573
rect 96709 2533 96721 2567
rect 96755 2564 96767 2567
rect 97718 2564 97724 2576
rect 96755 2536 97724 2564
rect 96755 2533 96767 2536
rect 96709 2527 96767 2533
rect 97718 2524 97724 2536
rect 97776 2524 97782 2576
rect 78677 2499 78735 2505
rect 77404 2468 77892 2496
rect 77113 2459 77171 2465
rect 50522 2388 50528 2440
rect 50580 2428 50586 2440
rect 52549 2431 52607 2437
rect 52549 2428 52561 2431
rect 50580 2400 52561 2428
rect 50580 2388 50586 2400
rect 52549 2397 52561 2400
rect 52595 2397 52607 2431
rect 52549 2391 52607 2397
rect 55950 2388 55956 2440
rect 56008 2428 56014 2440
rect 59357 2431 59415 2437
rect 59357 2428 59369 2431
rect 56008 2400 59369 2428
rect 56008 2388 56014 2400
rect 59357 2397 59369 2400
rect 59403 2397 59415 2431
rect 59357 2391 59415 2397
rect 63402 2388 63408 2440
rect 63460 2428 63466 2440
rect 63460 2400 71636 2428
rect 63460 2388 63466 2400
rect 47213 2323 47271 2329
rect 47320 2332 50200 2360
rect 40696 2264 41414 2292
rect 40497 2255 40555 2261
rect 41966 2252 41972 2304
rect 42024 2292 42030 2304
rect 45097 2295 45155 2301
rect 45097 2292 45109 2295
rect 42024 2264 45109 2292
rect 42024 2252 42030 2264
rect 45097 2261 45109 2264
rect 45143 2261 45155 2295
rect 45097 2255 45155 2261
rect 45462 2252 45468 2304
rect 45520 2292 45526 2304
rect 47320 2292 47348 2332
rect 50430 2320 50436 2372
rect 50488 2360 50494 2372
rect 54021 2363 54079 2369
rect 54021 2360 54033 2363
rect 50488 2332 54033 2360
rect 50488 2320 50494 2332
rect 54021 2329 54033 2332
rect 54067 2329 54079 2363
rect 54021 2323 54079 2329
rect 54110 2320 54116 2372
rect 54168 2360 54174 2372
rect 54168 2332 56732 2360
rect 54168 2320 54174 2332
rect 45520 2264 47348 2292
rect 45520 2252 45526 2264
rect 47394 2252 47400 2304
rect 47452 2292 47458 2304
rect 50985 2295 51043 2301
rect 50985 2292 50997 2295
rect 47452 2264 50997 2292
rect 47452 2252 47458 2264
rect 50985 2261 50997 2264
rect 51031 2261 51043 2295
rect 50985 2255 51043 2261
rect 51718 2252 51724 2304
rect 51776 2292 51782 2304
rect 55125 2295 55183 2301
rect 55125 2292 55137 2295
rect 51776 2264 55137 2292
rect 51776 2252 51782 2264
rect 55125 2261 55137 2264
rect 55171 2261 55183 2295
rect 56704 2292 56732 2332
rect 57146 2320 57152 2372
rect 57204 2360 57210 2372
rect 60277 2363 60335 2369
rect 60277 2360 60289 2363
rect 57204 2332 60289 2360
rect 57204 2320 57210 2332
rect 60277 2329 60289 2332
rect 60323 2329 60335 2363
rect 60277 2323 60335 2329
rect 60366 2320 60372 2372
rect 60424 2360 60430 2372
rect 61749 2363 61807 2369
rect 61749 2360 61761 2363
rect 60424 2332 61761 2360
rect 60424 2320 60430 2332
rect 61749 2329 61761 2332
rect 61795 2329 61807 2363
rect 61749 2323 61807 2329
rect 63310 2320 63316 2372
rect 63368 2360 63374 2372
rect 66349 2363 66407 2369
rect 66349 2360 66361 2363
rect 63368 2332 66361 2360
rect 63368 2320 63374 2332
rect 66349 2329 66361 2332
rect 66395 2329 66407 2363
rect 66349 2323 66407 2329
rect 66806 2320 66812 2372
rect 66864 2360 66870 2372
rect 68281 2363 68339 2369
rect 68281 2360 68293 2363
rect 66864 2332 68293 2360
rect 66864 2320 66870 2332
rect 68281 2329 68293 2332
rect 68327 2329 68339 2363
rect 68281 2323 68339 2329
rect 68462 2320 68468 2372
rect 68520 2360 68526 2372
rect 70029 2363 70087 2369
rect 70029 2360 70041 2363
rect 68520 2332 70041 2360
rect 68520 2320 68526 2332
rect 70029 2329 70041 2332
rect 70075 2329 70087 2363
rect 71225 2363 71283 2369
rect 71225 2360 71237 2363
rect 70029 2323 70087 2329
rect 70366 2332 71237 2360
rect 57701 2295 57759 2301
rect 57701 2292 57713 2295
rect 56704 2264 57713 2292
rect 55125 2255 55183 2261
rect 57701 2261 57713 2264
rect 57747 2261 57759 2295
rect 57701 2255 57759 2261
rect 58066 2252 58072 2304
rect 58124 2292 58130 2304
rect 58161 2295 58219 2301
rect 58161 2292 58173 2295
rect 58124 2264 58173 2292
rect 58124 2252 58130 2264
rect 58161 2261 58173 2264
rect 58207 2261 58219 2295
rect 58161 2255 58219 2261
rect 59630 2252 59636 2304
rect 59688 2292 59694 2304
rect 60734 2292 60740 2304
rect 59688 2264 60740 2292
rect 59688 2252 59694 2264
rect 60734 2252 60740 2264
rect 60792 2252 60798 2304
rect 62022 2252 62028 2304
rect 62080 2292 62086 2304
rect 63865 2295 63923 2301
rect 63865 2292 63877 2295
rect 62080 2264 63877 2292
rect 62080 2252 62086 2264
rect 63865 2261 63877 2264
rect 63911 2261 63923 2295
rect 63865 2255 63923 2261
rect 63954 2252 63960 2304
rect 64012 2292 64018 2304
rect 65797 2295 65855 2301
rect 65797 2292 65809 2295
rect 64012 2264 65809 2292
rect 64012 2252 64018 2264
rect 65797 2261 65809 2264
rect 65843 2261 65855 2295
rect 65797 2255 65855 2261
rect 66254 2252 66260 2304
rect 66312 2292 66318 2304
rect 69109 2295 69167 2301
rect 69109 2292 69121 2295
rect 66312 2264 69121 2292
rect 66312 2252 66318 2264
rect 69109 2261 69121 2264
rect 69155 2261 69167 2295
rect 69109 2255 69167 2261
rect 69290 2252 69296 2304
rect 69348 2292 69354 2304
rect 70366 2292 70394 2332
rect 71225 2329 71237 2332
rect 71271 2329 71283 2363
rect 71608 2360 71636 2400
rect 71682 2388 71688 2440
rect 71740 2428 71746 2440
rect 73893 2431 73951 2437
rect 73893 2428 73905 2431
rect 71740 2400 73905 2428
rect 71740 2388 71746 2400
rect 73893 2397 73905 2400
rect 73939 2397 73951 2431
rect 73893 2391 73951 2397
rect 74994 2388 75000 2440
rect 75052 2428 75058 2440
rect 77297 2431 77355 2437
rect 77297 2428 77309 2431
rect 75052 2400 77309 2428
rect 75052 2388 75058 2400
rect 77297 2397 77309 2400
rect 77343 2397 77355 2431
rect 77864 2428 77892 2468
rect 78677 2465 78689 2499
rect 78723 2496 78735 2499
rect 79137 2499 79195 2505
rect 79137 2496 79149 2499
rect 78723 2468 79149 2496
rect 78723 2465 78735 2468
rect 78677 2459 78735 2465
rect 79137 2465 79149 2468
rect 79183 2465 79195 2499
rect 79137 2459 79195 2465
rect 79226 2456 79232 2508
rect 79284 2496 79290 2508
rect 80425 2499 80483 2505
rect 80425 2496 80437 2499
rect 79284 2468 80437 2496
rect 79284 2456 79290 2468
rect 80425 2465 80437 2468
rect 80471 2465 80483 2499
rect 80425 2459 80483 2465
rect 84286 2456 84292 2508
rect 84344 2496 84350 2508
rect 84381 2499 84439 2505
rect 84381 2496 84393 2499
rect 84344 2468 84393 2496
rect 84344 2456 84350 2468
rect 84381 2465 84393 2468
rect 84427 2465 84439 2499
rect 84654 2496 84660 2508
rect 84615 2468 84660 2496
rect 84381 2459 84439 2465
rect 84654 2456 84660 2468
rect 84712 2456 84718 2508
rect 85298 2456 85304 2508
rect 85356 2496 85362 2508
rect 88429 2499 88487 2505
rect 88429 2496 88441 2499
rect 85356 2468 88441 2496
rect 85356 2456 85362 2468
rect 88429 2465 88441 2468
rect 88475 2465 88487 2499
rect 88610 2496 88616 2508
rect 88571 2468 88616 2496
rect 88429 2459 88487 2465
rect 88610 2456 88616 2468
rect 88668 2456 88674 2508
rect 88794 2456 88800 2508
rect 88852 2496 88858 2508
rect 90361 2499 90419 2505
rect 90361 2496 90373 2499
rect 88852 2468 90373 2496
rect 88852 2456 88858 2468
rect 90361 2465 90373 2468
rect 90407 2465 90419 2499
rect 92293 2499 92351 2505
rect 92293 2496 92305 2499
rect 90361 2459 90419 2465
rect 90468 2468 92305 2496
rect 79689 2431 79747 2437
rect 79689 2428 79701 2431
rect 77864 2400 79701 2428
rect 77297 2391 77355 2397
rect 79689 2397 79701 2400
rect 79735 2397 79747 2431
rect 79689 2391 79747 2397
rect 84746 2388 84752 2440
rect 84804 2428 84810 2440
rect 87969 2431 88027 2437
rect 87969 2428 87981 2431
rect 84804 2400 87981 2428
rect 84804 2388 84810 2400
rect 87969 2397 87981 2400
rect 88015 2397 88027 2431
rect 87969 2391 88027 2397
rect 88242 2388 88248 2440
rect 88300 2428 88306 2440
rect 90468 2428 90496 2468
rect 92293 2465 92305 2468
rect 92339 2465 92351 2499
rect 92293 2459 92351 2465
rect 92658 2456 92664 2508
rect 92716 2496 92722 2508
rect 93121 2499 93179 2505
rect 93121 2496 93133 2499
rect 92716 2468 93133 2496
rect 92716 2456 92722 2468
rect 93121 2465 93133 2468
rect 93167 2465 93179 2499
rect 94961 2499 95019 2505
rect 94961 2496 94973 2499
rect 93121 2459 93179 2465
rect 93826 2468 94973 2496
rect 88300 2400 90496 2428
rect 88300 2388 88306 2400
rect 91278 2388 91284 2440
rect 91336 2428 91342 2440
rect 93826 2428 93854 2468
rect 94961 2465 94973 2468
rect 95007 2465 95019 2499
rect 95786 2496 95792 2508
rect 95747 2468 95792 2496
rect 94961 2459 95019 2465
rect 95786 2456 95792 2468
rect 95844 2456 95850 2508
rect 96525 2499 96583 2505
rect 96525 2496 96537 2499
rect 96264 2468 96537 2496
rect 91336 2400 93854 2428
rect 91336 2388 91342 2400
rect 93946 2388 93952 2440
rect 94004 2428 94010 2440
rect 94222 2428 94228 2440
rect 94004 2400 94228 2428
rect 94004 2388 94010 2400
rect 94222 2388 94228 2400
rect 94280 2388 94286 2440
rect 94314 2388 94320 2440
rect 94372 2428 94378 2440
rect 96264 2437 96292 2468
rect 96525 2465 96537 2468
rect 96571 2465 96583 2499
rect 96525 2459 96583 2465
rect 97534 2456 97540 2508
rect 97592 2496 97598 2508
rect 97905 2499 97963 2505
rect 97905 2496 97917 2499
rect 97592 2468 97917 2496
rect 97592 2456 97598 2468
rect 97905 2465 97917 2468
rect 97951 2465 97963 2499
rect 97905 2459 97963 2465
rect 96249 2431 96307 2437
rect 96249 2428 96261 2431
rect 94372 2400 96261 2428
rect 94372 2388 94378 2400
rect 96249 2397 96261 2400
rect 96295 2397 96307 2431
rect 96249 2391 96307 2397
rect 72694 2360 72700 2372
rect 71608 2332 72700 2360
rect 71225 2323 71283 2329
rect 72694 2320 72700 2332
rect 72752 2320 72758 2372
rect 72878 2320 72884 2372
rect 72936 2360 72942 2372
rect 74353 2363 74411 2369
rect 74353 2360 74365 2363
rect 72936 2332 74365 2360
rect 72936 2320 72942 2332
rect 74353 2329 74365 2332
rect 74399 2329 74411 2363
rect 74353 2323 74411 2329
rect 74460 2332 75316 2360
rect 69348 2264 70394 2292
rect 69348 2252 69354 2264
rect 72142 2252 72148 2304
rect 72200 2292 72206 2304
rect 72237 2295 72295 2301
rect 72237 2292 72249 2295
rect 72200 2264 72249 2292
rect 72200 2252 72206 2264
rect 72237 2261 72249 2264
rect 72283 2261 72295 2295
rect 72510 2292 72516 2304
rect 72471 2264 72516 2292
rect 72237 2255 72295 2261
rect 72510 2252 72516 2264
rect 72568 2252 72574 2304
rect 73062 2252 73068 2304
rect 73120 2292 73126 2304
rect 74460 2292 74488 2332
rect 73120 2264 74488 2292
rect 75288 2292 75316 2332
rect 75454 2320 75460 2372
rect 75512 2360 75518 2372
rect 78953 2363 79011 2369
rect 78953 2360 78965 2363
rect 75512 2332 78965 2360
rect 75512 2320 75518 2332
rect 78953 2329 78965 2332
rect 78999 2329 79011 2363
rect 82814 2360 82820 2372
rect 82775 2332 82820 2360
rect 78953 2323 79011 2329
rect 82814 2320 82820 2332
rect 82872 2320 82878 2372
rect 87690 2320 87696 2372
rect 87748 2360 87754 2372
rect 91097 2363 91155 2369
rect 91097 2360 91109 2363
rect 87748 2332 91109 2360
rect 87748 2320 87754 2332
rect 91097 2329 91109 2332
rect 91143 2329 91155 2363
rect 91097 2323 91155 2329
rect 91204 2332 92520 2360
rect 76469 2295 76527 2301
rect 76469 2292 76481 2295
rect 75288 2264 76481 2292
rect 73120 2252 73126 2264
rect 76469 2261 76481 2264
rect 76515 2261 76527 2295
rect 78674 2292 78680 2304
rect 78587 2264 78680 2292
rect 76469 2255 76527 2261
rect 78674 2252 78680 2264
rect 78732 2292 78738 2304
rect 78769 2295 78827 2301
rect 78769 2292 78781 2295
rect 78732 2264 78781 2292
rect 78732 2252 78738 2264
rect 78769 2261 78781 2264
rect 78815 2261 78827 2295
rect 78769 2255 78827 2261
rect 82265 2295 82323 2301
rect 82265 2261 82277 2295
rect 82311 2292 82323 2295
rect 83366 2292 83372 2304
rect 82311 2264 83372 2292
rect 82311 2261 82323 2264
rect 82265 2255 82323 2261
rect 83366 2252 83372 2264
rect 83424 2252 83430 2304
rect 84010 2252 84016 2304
rect 84068 2292 84074 2304
rect 87141 2295 87199 2301
rect 87141 2292 87153 2295
rect 84068 2264 87153 2292
rect 84068 2252 84074 2264
rect 87141 2261 87153 2264
rect 87187 2261 87199 2295
rect 88334 2292 88340 2304
rect 88295 2264 88340 2292
rect 87141 2255 87199 2261
rect 88334 2252 88340 2264
rect 88392 2292 88398 2304
rect 88610 2292 88616 2304
rect 88392 2264 88616 2292
rect 88392 2252 88398 2264
rect 88610 2252 88616 2264
rect 88668 2292 88674 2304
rect 88797 2295 88855 2301
rect 88797 2292 88809 2295
rect 88668 2264 88809 2292
rect 88668 2252 88674 2264
rect 88797 2261 88809 2264
rect 88843 2261 88855 2295
rect 88797 2255 88855 2261
rect 88886 2252 88892 2304
rect 88944 2292 88950 2304
rect 91204 2292 91232 2332
rect 88944 2264 91232 2292
rect 92492 2292 92520 2332
rect 92566 2320 92572 2372
rect 92624 2360 92630 2372
rect 95973 2363 96031 2369
rect 95973 2360 95985 2363
rect 92624 2332 95985 2360
rect 92624 2320 92630 2332
rect 95973 2329 95985 2332
rect 96019 2329 96031 2363
rect 95973 2323 96031 2329
rect 98089 2363 98147 2369
rect 98089 2329 98101 2363
rect 98135 2360 98147 2363
rect 99650 2360 99656 2372
rect 98135 2332 99656 2360
rect 98135 2329 98147 2332
rect 98089 2323 98147 2329
rect 99650 2320 99656 2332
rect 99708 2320 99714 2372
rect 93213 2295 93271 2301
rect 93213 2292 93225 2295
rect 92492 2264 93225 2292
rect 88944 2252 88950 2264
rect 93213 2261 93225 2264
rect 93259 2261 93271 2295
rect 93213 2255 93271 2261
rect 93302 2252 93308 2304
rect 93360 2292 93366 2304
rect 93949 2295 94007 2301
rect 93949 2292 93961 2295
rect 93360 2264 93961 2292
rect 93360 2252 93366 2264
rect 93949 2261 93961 2264
rect 93995 2261 94007 2295
rect 93949 2255 94007 2261
rect 1104 2202 98808 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 65686 2202
rect 65738 2150 65750 2202
rect 65802 2150 65814 2202
rect 65866 2150 65878 2202
rect 65930 2150 96406 2202
rect 96458 2150 96470 2202
rect 96522 2150 96534 2202
rect 96586 2150 96598 2202
rect 96650 2150 98808 2202
rect 1104 2128 98808 2150
rect 18414 2048 18420 2100
rect 18472 2088 18478 2100
rect 31754 2088 31760 2100
rect 18472 2060 31760 2088
rect 18472 2048 18478 2060
rect 31754 2048 31760 2060
rect 31812 2048 31818 2100
rect 48682 2048 48688 2100
rect 48740 2088 48746 2100
rect 51537 2091 51595 2097
rect 51537 2088 51549 2091
rect 48740 2060 51549 2088
rect 48740 2048 48746 2060
rect 51537 2057 51549 2060
rect 51583 2057 51595 2091
rect 51537 2051 51595 2057
rect 51626 2048 51632 2100
rect 51684 2088 51690 2100
rect 56410 2088 56416 2100
rect 51684 2060 56416 2088
rect 51684 2048 51690 2060
rect 56410 2048 56416 2060
rect 56468 2048 56474 2100
rect 61194 2048 61200 2100
rect 61252 2088 61258 2100
rect 61746 2088 61752 2100
rect 61252 2060 61752 2088
rect 61252 2048 61258 2060
rect 61746 2048 61752 2060
rect 61804 2048 61810 2100
rect 62114 2048 62120 2100
rect 62172 2088 62178 2100
rect 63954 2088 63960 2100
rect 62172 2060 63960 2088
rect 62172 2048 62178 2060
rect 63954 2048 63960 2060
rect 64012 2048 64018 2100
rect 67542 2048 67548 2100
rect 67600 2088 67606 2100
rect 69290 2088 69296 2100
rect 67600 2060 69296 2088
rect 67600 2048 67606 2060
rect 69290 2048 69296 2060
rect 69348 2048 69354 2100
rect 70026 2048 70032 2100
rect 70084 2088 70090 2100
rect 71682 2088 71688 2100
rect 70084 2060 71688 2088
rect 70084 2048 70090 2060
rect 71682 2048 71688 2060
rect 71740 2048 71746 2100
rect 76374 2048 76380 2100
rect 76432 2088 76438 2100
rect 80422 2088 80428 2100
rect 76432 2060 80428 2088
rect 76432 2048 76438 2060
rect 80422 2048 80428 2060
rect 80480 2048 80486 2100
rect 81158 2048 81164 2100
rect 81216 2088 81222 2100
rect 82722 2088 82728 2100
rect 81216 2060 82728 2088
rect 81216 2048 81222 2060
rect 82722 2048 82728 2060
rect 82780 2048 82786 2100
rect 89530 2048 89536 2100
rect 89588 2088 89594 2100
rect 93302 2088 93308 2100
rect 89588 2060 93308 2088
rect 89588 2048 89594 2060
rect 93302 2048 93308 2060
rect 93360 2048 93366 2100
rect 2038 1980 2044 2032
rect 2096 2020 2102 2032
rect 2096 1992 26740 2020
rect 2096 1980 2102 1992
rect 3970 1912 3976 1964
rect 4028 1952 4034 1964
rect 4338 1952 4344 1964
rect 4028 1924 4344 1952
rect 4028 1912 4034 1924
rect 4338 1912 4344 1924
rect 4396 1912 4402 1964
rect 21266 1912 21272 1964
rect 21324 1952 21330 1964
rect 26234 1952 26240 1964
rect 21324 1924 26240 1952
rect 21324 1912 21330 1924
rect 26234 1912 26240 1924
rect 26292 1912 26298 1964
rect 25314 1844 25320 1896
rect 25372 1884 25378 1896
rect 26712 1884 26740 1992
rect 27246 1980 27252 2032
rect 27304 2020 27310 2032
rect 31294 2020 31300 2032
rect 27304 1992 31300 2020
rect 27304 1980 27310 1992
rect 31294 1980 31300 1992
rect 31352 1980 31358 2032
rect 31662 1980 31668 2032
rect 31720 2020 31726 2032
rect 33042 2020 33048 2032
rect 31720 1992 33048 2020
rect 31720 1980 31726 1992
rect 33042 1980 33048 1992
rect 33100 1980 33106 2032
rect 38562 2020 38568 2032
rect 35866 1992 38568 2020
rect 26786 1912 26792 1964
rect 26844 1952 26850 1964
rect 35866 1952 35894 1992
rect 38562 1980 38568 1992
rect 38620 1980 38626 2032
rect 54386 1980 54392 2032
rect 54444 2020 54450 2032
rect 63402 2020 63408 2032
rect 54444 1992 63408 2020
rect 54444 1980 54450 1992
rect 63402 1980 63408 1992
rect 63460 1980 63466 2032
rect 68738 1980 68744 2032
rect 68796 2020 68802 2032
rect 72510 2020 72516 2032
rect 68796 1992 72516 2020
rect 68796 1980 68802 1992
rect 72510 1980 72516 1992
rect 72568 1980 72574 2032
rect 72694 1980 72700 2032
rect 72752 2020 72758 2032
rect 78674 2020 78680 2032
rect 72752 1992 78680 2020
rect 72752 1980 72758 1992
rect 78674 1980 78680 1992
rect 78732 1980 78738 2032
rect 26844 1924 35894 1952
rect 26844 1912 26850 1924
rect 47670 1912 47676 1964
rect 47728 1952 47734 1964
rect 53834 1952 53840 1964
rect 47728 1924 53840 1952
rect 47728 1912 47734 1924
rect 53834 1912 53840 1924
rect 53892 1912 53898 1964
rect 71774 1912 71780 1964
rect 71832 1952 71838 1964
rect 82262 1952 82268 1964
rect 71832 1924 82268 1952
rect 71832 1912 71838 1924
rect 82262 1912 82268 1924
rect 82320 1912 82326 1964
rect 33502 1884 33508 1896
rect 25372 1856 26234 1884
rect 26712 1856 33508 1884
rect 25372 1844 25378 1856
rect 26206 1816 26234 1856
rect 33502 1844 33508 1856
rect 33560 1844 33566 1896
rect 51902 1844 51908 1896
rect 51960 1884 51966 1896
rect 52638 1884 52644 1896
rect 51960 1856 52644 1884
rect 51960 1844 51966 1856
rect 52638 1844 52644 1856
rect 52696 1844 52702 1896
rect 66346 1844 66352 1896
rect 66404 1884 66410 1896
rect 76558 1884 76564 1896
rect 66404 1856 76564 1884
rect 66404 1844 66410 1856
rect 76558 1844 76564 1856
rect 76616 1844 76622 1896
rect 31478 1816 31484 1828
rect 26206 1788 31484 1816
rect 31478 1776 31484 1788
rect 31536 1776 31542 1828
rect 18046 1708 18052 1760
rect 18104 1748 18110 1760
rect 33318 1748 33324 1760
rect 18104 1720 33324 1748
rect 18104 1708 18110 1720
rect 33318 1708 33324 1720
rect 33376 1708 33382 1760
rect 35250 1436 35256 1488
rect 35308 1476 35314 1488
rect 37182 1476 37188 1488
rect 35308 1448 37188 1476
rect 35308 1436 35314 1448
rect 37182 1436 37188 1448
rect 37240 1436 37246 1488
rect 58434 1436 58440 1488
rect 58492 1476 58498 1488
rect 60366 1476 60372 1488
rect 58492 1448 60372 1476
rect 58492 1436 58498 1448
rect 60366 1436 60372 1448
rect 60424 1436 60430 1488
rect 65702 1436 65708 1488
rect 65760 1476 65766 1488
rect 66254 1476 66260 1488
rect 65760 1448 66260 1476
rect 65760 1436 65766 1448
rect 66254 1436 66260 1448
rect 66312 1436 66318 1488
rect 66346 1436 66352 1488
rect 66404 1476 66410 1488
rect 68462 1476 68468 1488
rect 66404 1448 68468 1476
rect 66404 1436 66410 1448
rect 68462 1436 68468 1448
rect 68520 1436 68526 1488
rect 74258 1436 74264 1488
rect 74316 1476 74322 1488
rect 74718 1476 74724 1488
rect 74316 1448 74724 1476
rect 74316 1436 74322 1448
rect 74718 1436 74724 1448
rect 74776 1436 74782 1488
rect 32766 1368 32772 1420
rect 32824 1408 32830 1420
rect 33962 1408 33968 1420
rect 32824 1380 33968 1408
rect 32824 1368 32830 1380
rect 33962 1368 33968 1380
rect 34020 1368 34026 1420
rect 34054 1368 34060 1420
rect 34112 1408 34118 1420
rect 34698 1408 34704 1420
rect 34112 1380 34704 1408
rect 34112 1368 34118 1380
rect 34698 1368 34704 1380
rect 34756 1368 34762 1420
rect 36446 1368 36452 1420
rect 36504 1408 36510 1420
rect 37918 1408 37924 1420
rect 36504 1380 37924 1408
rect 36504 1368 36510 1380
rect 37918 1368 37924 1380
rect 37976 1368 37982 1420
rect 48682 1368 48688 1420
rect 48740 1408 48746 1420
rect 50522 1408 50528 1420
rect 48740 1380 50528 1408
rect 48740 1368 48746 1380
rect 50522 1368 50528 1380
rect 50580 1368 50586 1420
rect 52914 1368 52920 1420
rect 52972 1408 52978 1420
rect 54018 1408 54024 1420
rect 52972 1380 54024 1408
rect 52972 1368 52978 1380
rect 54018 1368 54024 1380
rect 54076 1368 54082 1420
rect 60182 1368 60188 1420
rect 60240 1408 60246 1420
rect 62022 1408 62028 1420
rect 60240 1380 62028 1408
rect 60240 1368 60246 1380
rect 62022 1368 62028 1380
rect 62080 1368 62086 1420
rect 65058 1368 65064 1420
rect 65116 1408 65122 1420
rect 66806 1408 66812 1420
rect 65116 1380 66812 1408
rect 65116 1368 65122 1380
rect 66806 1368 66812 1380
rect 66864 1368 66870 1420
rect 71222 1368 71228 1420
rect 71280 1408 71286 1420
rect 72878 1408 72884 1420
rect 71280 1380 72884 1408
rect 71280 1368 71286 1380
rect 72878 1368 72884 1380
rect 72936 1368 72942 1420
rect 73614 1368 73620 1420
rect 73672 1408 73678 1420
rect 74994 1408 75000 1420
rect 73672 1380 75000 1408
rect 73672 1368 73678 1380
rect 74994 1368 75000 1380
rect 75052 1368 75058 1420
rect 77294 1368 77300 1420
rect 77352 1408 77358 1420
rect 79226 1408 79232 1420
rect 77352 1380 79232 1408
rect 77352 1368 77358 1380
rect 79226 1368 79232 1380
rect 79284 1368 79290 1420
rect 16390 1300 16396 1352
rect 16448 1340 16454 1352
rect 30282 1340 30288 1352
rect 16448 1312 30288 1340
rect 16448 1300 16454 1312
rect 30282 1300 30288 1312
rect 30340 1300 30346 1352
rect 31754 1300 31760 1352
rect 31812 1340 31818 1352
rect 43622 1340 43628 1352
rect 31812 1312 43628 1340
rect 31812 1300 31818 1312
rect 43622 1300 43628 1312
rect 43680 1300 43686 1352
rect 48958 1300 48964 1352
rect 49016 1340 49022 1352
rect 58066 1340 58072 1352
rect 49016 1312 58072 1340
rect 49016 1300 49022 1312
rect 58066 1300 58072 1312
rect 58124 1300 58130 1352
rect 58161 1343 58219 1349
rect 58161 1309 58173 1343
rect 58207 1340 58219 1343
rect 59722 1340 59728 1352
rect 58207 1312 59728 1340
rect 58207 1309 58219 1312
rect 58161 1303 58219 1309
rect 59722 1300 59728 1312
rect 59780 1300 59786 1352
rect 62390 1300 62396 1352
rect 62448 1340 62454 1352
rect 91370 1340 91376 1352
rect 62448 1312 91376 1340
rect 62448 1300 62454 1312
rect 91370 1300 91376 1312
rect 91428 1300 91434 1352
rect 38562 1232 38568 1284
rect 38620 1272 38626 1284
rect 43070 1272 43076 1284
rect 38620 1244 43076 1272
rect 38620 1232 38626 1244
rect 43070 1232 43076 1244
rect 43128 1232 43134 1284
rect 43254 1232 43260 1284
rect 43312 1272 43318 1284
rect 49421 1275 49479 1281
rect 49421 1272 49433 1275
rect 43312 1244 49433 1272
rect 43312 1232 43318 1244
rect 49421 1241 49433 1244
rect 49467 1241 49479 1275
rect 65242 1272 65248 1284
rect 49421 1235 49479 1241
rect 51046 1244 65248 1272
rect 25866 1164 25872 1216
rect 25924 1204 25930 1216
rect 25924 1176 26234 1204
rect 25924 1164 25930 1176
rect 26206 1136 26234 1176
rect 36722 1164 36728 1216
rect 36780 1204 36786 1216
rect 51046 1204 51074 1244
rect 65242 1232 65248 1244
rect 65300 1232 65306 1284
rect 36780 1176 51074 1204
rect 51537 1207 51595 1213
rect 36780 1164 36786 1176
rect 51537 1173 51549 1207
rect 51583 1204 51595 1207
rect 72142 1204 72148 1216
rect 51583 1176 72148 1204
rect 51583 1173 51595 1176
rect 51537 1167 51595 1173
rect 72142 1164 72148 1176
rect 72200 1164 72206 1216
rect 40589 1139 40647 1145
rect 40589 1136 40601 1139
rect 26206 1108 40601 1136
rect 40589 1105 40601 1108
rect 40635 1105 40647 1139
rect 40589 1099 40647 1105
rect 40681 1139 40739 1145
rect 40681 1105 40693 1139
rect 40727 1136 40739 1139
rect 58342 1136 58348 1148
rect 40727 1108 58348 1136
rect 40727 1105 40739 1108
rect 40681 1099 40739 1105
rect 58342 1096 58348 1108
rect 58400 1096 58406 1148
rect 63586 1096 63592 1148
rect 63644 1136 63650 1148
rect 95786 1136 95792 1148
rect 63644 1108 95792 1136
rect 63644 1096 63650 1108
rect 95786 1096 95792 1108
rect 95844 1096 95850 1148
rect 12342 1028 12348 1080
rect 12400 1068 12406 1080
rect 58161 1071 58219 1077
rect 58161 1068 58173 1071
rect 12400 1040 58173 1068
rect 12400 1028 12406 1040
rect 58161 1037 58173 1040
rect 58207 1037 58219 1071
rect 58161 1031 58219 1037
rect 58250 1028 58256 1080
rect 58308 1068 58314 1080
rect 92658 1068 92664 1080
rect 58308 1040 92664 1068
rect 58308 1028 58314 1040
rect 92658 1028 92664 1040
rect 92716 1028 92722 1080
rect 26050 960 26056 1012
rect 26108 1000 26114 1012
rect 70670 1000 70676 1012
rect 26108 972 70676 1000
rect 26108 960 26114 972
rect 70670 960 70676 972
rect 70728 960 70734 1012
rect 9306 892 9312 944
rect 9364 932 9370 944
rect 31021 935 31079 941
rect 31021 932 31033 935
rect 9364 904 31033 932
rect 9364 892 9370 904
rect 31021 901 31033 904
rect 31067 901 31079 935
rect 31021 895 31079 901
rect 33870 892 33876 944
rect 33928 932 33934 944
rect 40681 935 40739 941
rect 40681 932 40693 935
rect 33928 904 40693 932
rect 33928 892 33934 904
rect 40681 901 40693 904
rect 40727 901 40739 935
rect 40681 895 40739 901
rect 40773 935 40831 941
rect 40773 901 40785 935
rect 40819 932 40831 935
rect 44266 932 44272 944
rect 40819 904 44272 932
rect 40819 901 40831 904
rect 40773 895 40831 901
rect 44266 892 44272 904
rect 44324 892 44330 944
rect 46658 892 46664 944
rect 46716 932 46722 944
rect 89806 932 89812 944
rect 46716 904 89812 932
rect 46716 892 46722 904
rect 89806 892 89812 904
rect 89864 892 89870 944
rect 13630 824 13636 876
rect 13688 864 13694 876
rect 53006 864 53012 876
rect 13688 836 53012 864
rect 13688 824 13694 836
rect 53006 824 53012 836
rect 53064 824 53070 876
rect 59262 824 59268 876
rect 59320 864 59326 876
rect 88334 864 88340 876
rect 59320 836 88340 864
rect 59320 824 59326 836
rect 88334 824 88340 836
rect 88392 824 88398 876
rect 34514 756 34520 808
rect 34572 796 34578 808
rect 73522 796 73528 808
rect 34572 768 73528 796
rect 34572 756 34578 768
rect 73522 756 73528 768
rect 73580 756 73586 808
rect 25590 688 25596 740
rect 25648 728 25654 740
rect 62206 728 62212 740
rect 25648 700 62212 728
rect 25648 688 25654 700
rect 62206 688 62212 700
rect 62264 688 62270 740
rect 20438 620 20444 672
rect 20496 660 20502 672
rect 20496 632 40724 660
rect 20496 620 20502 632
rect 2590 552 2596 604
rect 2648 592 2654 604
rect 37734 592 37740 604
rect 2648 564 37740 592
rect 2648 552 2654 564
rect 37734 552 37740 564
rect 37792 592 37798 604
rect 38562 592 38568 604
rect 37792 564 38568 592
rect 37792 552 37798 564
rect 38562 552 38568 564
rect 38620 552 38626 604
rect 40696 592 40724 632
rect 42242 620 42248 672
rect 42300 660 42306 672
rect 78030 660 78036 672
rect 42300 632 78036 660
rect 42300 620 42306 632
rect 78030 620 78036 632
rect 78088 620 78094 672
rect 44910 592 44916 604
rect 40696 564 44916 592
rect 44910 552 44916 564
rect 44968 552 44974 604
rect 46109 595 46167 601
rect 46109 561 46121 595
rect 46155 592 46167 595
rect 50798 592 50804 604
rect 46155 564 50804 592
rect 46155 561 46167 564
rect 46109 555 46167 561
rect 50798 552 50804 564
rect 50856 552 50862 604
rect 71498 592 71504 604
rect 51046 564 71504 592
rect 15654 484 15660 536
rect 15712 524 15718 536
rect 45005 527 45063 533
rect 15712 496 44864 524
rect 15712 484 15718 496
rect 38378 416 38384 468
rect 38436 456 38442 468
rect 44729 459 44787 465
rect 44729 456 44741 459
rect 38436 428 44741 456
rect 38436 416 38442 428
rect 44729 425 44741 428
rect 44775 425 44787 459
rect 44836 456 44864 496
rect 45005 493 45017 527
rect 45051 524 45063 527
rect 51046 524 51074 564
rect 71498 552 71504 564
rect 71556 552 71562 604
rect 45051 496 51074 524
rect 45051 493 45063 496
rect 45005 487 45063 493
rect 54846 484 54852 536
rect 54904 524 54910 536
rect 71314 524 71320 536
rect 54904 496 71320 524
rect 54904 484 54910 496
rect 71314 484 71320 496
rect 71372 484 71378 536
rect 49326 456 49332 468
rect 44836 428 49332 456
rect 44729 419 44787 425
rect 49326 416 49332 428
rect 49384 416 49390 468
rect 49421 459 49479 465
rect 49421 425 49433 459
rect 49467 456 49479 459
rect 72326 456 72332 468
rect 49467 428 72332 456
rect 49467 425 49479 428
rect 49421 419 49479 425
rect 72326 416 72332 428
rect 72384 416 72390 468
rect 6454 348 6460 400
rect 6512 388 6518 400
rect 92474 388 92480 400
rect 6512 360 92480 388
rect 6512 348 6518 360
rect 92474 348 92480 360
rect 92532 348 92538 400
rect 25958 280 25964 332
rect 26016 320 26022 332
rect 92842 320 92848 332
rect 26016 292 92848 320
rect 26016 280 26022 292
rect 92842 280 92848 292
rect 92900 280 92906 332
rect 5258 212 5264 264
rect 5316 252 5322 264
rect 62390 252 62396 264
rect 5316 224 62396 252
rect 5316 212 5322 224
rect 62390 212 62396 224
rect 62448 212 62454 264
rect 20254 144 20260 196
rect 20312 184 20318 196
rect 73706 184 73712 196
rect 20312 156 73712 184
rect 20312 144 20318 156
rect 73706 144 73712 156
rect 73764 144 73770 196
rect 16206 76 16212 128
rect 16264 116 16270 128
rect 46109 119 46167 125
rect 46109 116 46121 119
rect 16264 88 46121 116
rect 16264 76 16270 88
rect 46109 85 46121 88
rect 46155 85 46167 119
rect 46109 79 46167 85
rect 48774 76 48780 128
rect 48832 116 48838 128
rect 87138 116 87144 128
rect 48832 88 87144 116
rect 48832 76 48838 88
rect 87138 76 87144 88
rect 87196 76 87202 128
rect 31021 51 31079 57
rect 31021 17 31033 51
rect 31067 48 31079 51
rect 37550 48 37556 60
rect 31067 20 37556 48
rect 31067 17 31079 20
rect 31021 11 31079 17
rect 37550 8 37556 20
rect 37608 48 37614 60
rect 38378 48 38384 60
rect 37608 20 38384 48
rect 37608 8 37614 20
rect 38378 8 38384 20
rect 38436 8 38442 60
rect 39758 8 39764 60
rect 39816 48 39822 60
rect 70854 48 70860 60
rect 39816 20 70860 48
rect 39816 8 39822 20
rect 70854 8 70860 20
rect 70912 8 70918 60
<< via1 >>
rect 37464 39584 37516 39636
rect 40776 39380 40828 39432
rect 55496 39380 55548 39432
rect 44732 39312 44784 39364
rect 46480 39312 46532 39364
rect 61108 39312 61160 39364
rect 21916 39244 21968 39296
rect 89444 39244 89496 39296
rect 13728 39176 13780 39228
rect 41972 39176 42024 39228
rect 30104 39108 30156 39160
rect 59452 39108 59504 39160
rect 32864 39040 32916 39092
rect 25688 38972 25740 39024
rect 23940 38904 23992 38956
rect 10784 38836 10836 38888
rect 38476 38836 38528 38888
rect 48688 38904 48740 38956
rect 50068 38904 50120 38956
rect 76288 38836 76340 38888
rect 19984 38768 20036 38820
rect 13912 38700 13964 38752
rect 90456 38700 90508 38752
rect 93124 38632 93176 38684
rect 27988 38564 28040 38616
rect 36636 38564 36688 38616
rect 68836 38564 68888 38616
rect 23296 38496 23348 38548
rect 54300 38496 54352 38548
rect 18696 38428 18748 38480
rect 74816 38428 74868 38480
rect 16488 38360 16540 38412
rect 75736 38360 75788 38412
rect 88984 38360 89036 38412
rect 89628 38360 89680 38412
rect 32588 38292 32640 38344
rect 90916 38292 90968 38344
rect 17500 38224 17552 38276
rect 81992 38224 82044 38276
rect 15384 38156 15436 38208
rect 86224 38156 86276 38208
rect 4344 38088 4396 38140
rect 16856 38088 16908 38140
rect 10416 38020 10468 38072
rect 17960 38088 18012 38140
rect 19248 38088 19300 38140
rect 93584 38088 93636 38140
rect 24952 38020 25004 38072
rect 26148 38020 26200 38072
rect 30564 38020 30616 38072
rect 31576 38020 31628 38072
rect 47860 38020 47912 38072
rect 57796 38020 57848 38072
rect 71504 38020 71556 38072
rect 15108 37952 15160 38004
rect 42248 37952 42300 38004
rect 45284 37952 45336 38004
rect 11060 37884 11112 37936
rect 3332 37816 3384 37868
rect 37372 37816 37424 37868
rect 39120 37884 39172 37936
rect 50712 37952 50764 38004
rect 70400 37952 70452 38004
rect 40316 37816 40368 37868
rect 7012 37748 7064 37800
rect 13820 37748 13872 37800
rect 14924 37748 14976 37800
rect 34704 37748 34756 37800
rect 37096 37748 37148 37800
rect 41696 37791 41748 37800
rect 5724 37723 5776 37732
rect 5724 37689 5733 37723
rect 5733 37689 5767 37723
rect 5767 37689 5776 37723
rect 5724 37680 5776 37689
rect 12348 37680 12400 37732
rect 17684 37680 17736 37732
rect 25504 37680 25556 37732
rect 26516 37723 26568 37732
rect 26516 37689 26525 37723
rect 26525 37689 26559 37723
rect 26559 37689 26568 37723
rect 26516 37680 26568 37689
rect 27068 37680 27120 37732
rect 31208 37680 31260 37732
rect 31392 37723 31444 37732
rect 31392 37689 31401 37723
rect 31401 37689 31435 37723
rect 31435 37689 31444 37723
rect 31392 37680 31444 37689
rect 40040 37723 40092 37732
rect 40040 37689 40049 37723
rect 40049 37689 40083 37723
rect 40083 37689 40092 37723
rect 40040 37680 40092 37689
rect 41696 37757 41705 37791
rect 41705 37757 41739 37791
rect 41739 37757 41748 37791
rect 41696 37748 41748 37757
rect 42340 37791 42392 37800
rect 42340 37757 42349 37791
rect 42349 37757 42383 37791
rect 42383 37757 42392 37791
rect 42340 37748 42392 37757
rect 86040 37884 86092 37936
rect 48412 37816 48464 37868
rect 56048 37816 56100 37868
rect 66444 37816 66496 37868
rect 66536 37748 66588 37800
rect 75368 37748 75420 37800
rect 96068 37748 96120 37800
rect 70124 37680 70176 37732
rect 74264 37723 74316 37732
rect 74264 37689 74273 37723
rect 74273 37689 74307 37723
rect 74307 37689 74316 37723
rect 74264 37680 74316 37689
rect 75460 37680 75512 37732
rect 79048 37680 79100 37732
rect 81808 37680 81860 37732
rect 4712 37612 4764 37664
rect 8392 37612 8444 37664
rect 8484 37612 8536 37664
rect 15936 37612 15988 37664
rect 23020 37612 23072 37664
rect 36176 37612 36228 37664
rect 38936 37612 38988 37664
rect 42524 37612 42576 37664
rect 43076 37612 43128 37664
rect 48504 37655 48556 37664
rect 48504 37621 48513 37655
rect 48513 37621 48547 37655
rect 48547 37621 48556 37655
rect 48504 37612 48556 37621
rect 52368 37655 52420 37664
rect 52368 37621 52377 37655
rect 52377 37621 52411 37655
rect 52411 37621 52420 37655
rect 52368 37612 52420 37621
rect 54944 37612 54996 37664
rect 63776 37655 63828 37664
rect 63776 37621 63785 37655
rect 63785 37621 63819 37655
rect 63819 37621 63828 37655
rect 63776 37612 63828 37621
rect 64880 37612 64932 37664
rect 76932 37612 76984 37664
rect 80244 37612 80296 37664
rect 85212 37612 85264 37664
rect 86960 37680 87012 37732
rect 97632 37680 97684 37732
rect 87052 37612 87104 37664
rect 87880 37612 87932 37664
rect 90548 37612 90600 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 50326 37510 50378 37562
rect 50390 37510 50442 37562
rect 50454 37510 50506 37562
rect 50518 37510 50570 37562
rect 81046 37510 81098 37562
rect 81110 37510 81162 37562
rect 81174 37510 81226 37562
rect 81238 37510 81290 37562
rect 1400 37408 1452 37460
rect 6460 37408 6512 37460
rect 8392 37408 8444 37460
rect 388 37340 440 37392
rect 3884 37340 3936 37392
rect 7012 37383 7064 37392
rect 2964 37315 3016 37324
rect 2964 37281 2973 37315
rect 2973 37281 3007 37315
rect 3007 37281 3016 37315
rect 2964 37272 3016 37281
rect 4344 37315 4396 37324
rect 4344 37281 4353 37315
rect 4353 37281 4387 37315
rect 4387 37281 4396 37315
rect 4344 37272 4396 37281
rect 5448 37272 5500 37324
rect 5724 37315 5776 37324
rect 5724 37281 5733 37315
rect 5733 37281 5767 37315
rect 5767 37281 5776 37315
rect 5724 37272 5776 37281
rect 7012 37349 7021 37383
rect 7021 37349 7055 37383
rect 7055 37349 7064 37383
rect 7012 37340 7064 37349
rect 8484 37383 8536 37392
rect 8484 37349 8493 37383
rect 8493 37349 8527 37383
rect 8527 37349 8536 37383
rect 8484 37340 8536 37349
rect 9128 37340 9180 37392
rect 10784 37408 10836 37460
rect 11060 37451 11112 37460
rect 11060 37417 11069 37451
rect 11069 37417 11103 37451
rect 11103 37417 11112 37451
rect 11060 37408 11112 37417
rect 11704 37408 11756 37460
rect 16488 37451 16540 37460
rect 16488 37417 16497 37451
rect 16497 37417 16531 37451
rect 16531 37417 16540 37451
rect 16488 37408 16540 37417
rect 17040 37408 17092 37460
rect 17960 37408 18012 37460
rect 22284 37408 22336 37460
rect 23204 37408 23256 37460
rect 2320 37204 2372 37256
rect 11152 37340 11204 37392
rect 12348 37383 12400 37392
rect 12348 37349 12357 37383
rect 12357 37349 12391 37383
rect 12391 37349 12400 37383
rect 12348 37340 12400 37349
rect 13912 37340 13964 37392
rect 14372 37340 14424 37392
rect 15108 37383 15160 37392
rect 15108 37349 15117 37383
rect 15117 37349 15151 37383
rect 15151 37349 15160 37383
rect 15108 37340 15160 37349
rect 16120 37340 16172 37392
rect 17684 37383 17736 37392
rect 17684 37349 17693 37383
rect 17693 37349 17727 37383
rect 17727 37349 17736 37383
rect 17684 37340 17736 37349
rect 18788 37340 18840 37392
rect 19248 37383 19300 37392
rect 19248 37349 19257 37383
rect 19257 37349 19291 37383
rect 19291 37349 19300 37383
rect 19248 37340 19300 37349
rect 19892 37340 19944 37392
rect 21364 37340 21416 37392
rect 23020 37383 23072 37392
rect 23020 37349 23029 37383
rect 23029 37349 23063 37383
rect 23063 37349 23072 37383
rect 23020 37340 23072 37349
rect 10968 37272 11020 37324
rect 13544 37315 13596 37324
rect 13544 37281 13553 37315
rect 13553 37281 13587 37315
rect 13587 37281 13596 37315
rect 13544 37272 13596 37281
rect 20812 37272 20864 37324
rect 24032 37340 24084 37392
rect 24860 37408 24912 37460
rect 25872 37408 25924 37460
rect 28448 37408 28500 37460
rect 30196 37408 30248 37460
rect 31208 37408 31260 37460
rect 32772 37408 32824 37460
rect 34704 37451 34756 37460
rect 34704 37417 34713 37451
rect 34713 37417 34747 37451
rect 34747 37417 34756 37451
rect 34704 37408 34756 37417
rect 35440 37408 35492 37460
rect 37372 37451 37424 37460
rect 37372 37417 37381 37451
rect 37381 37417 37415 37451
rect 37415 37417 37424 37451
rect 37372 37408 37424 37417
rect 38108 37408 38160 37460
rect 40040 37451 40092 37460
rect 40040 37417 40049 37451
rect 40049 37417 40083 37451
rect 40083 37417 40092 37451
rect 40040 37408 40092 37417
rect 40684 37408 40736 37460
rect 42524 37451 42576 37460
rect 42524 37417 42533 37451
rect 42533 37417 42567 37451
rect 42567 37417 42576 37451
rect 42524 37408 42576 37417
rect 26516 37383 26568 37392
rect 26516 37349 26525 37383
rect 26525 37349 26559 37383
rect 26559 37349 26568 37383
rect 26516 37340 26568 37349
rect 27528 37340 27580 37392
rect 30932 37340 30984 37392
rect 31392 37340 31444 37392
rect 31944 37340 31996 37392
rect 34520 37340 34572 37392
rect 41328 37340 41380 37392
rect 41604 37340 41656 37392
rect 45284 37451 45336 37460
rect 45284 37417 45293 37451
rect 45293 37417 45327 37451
rect 45327 37417 45336 37451
rect 45284 37408 45336 37417
rect 45928 37408 45980 37460
rect 47860 37451 47912 37460
rect 47860 37417 47869 37451
rect 47869 37417 47903 37451
rect 47903 37417 47912 37451
rect 47860 37408 47912 37417
rect 48596 37451 48648 37460
rect 48596 37417 48605 37451
rect 48605 37417 48639 37451
rect 48639 37417 48648 37451
rect 48596 37408 48648 37417
rect 50712 37408 50764 37460
rect 51264 37451 51316 37460
rect 51264 37417 51273 37451
rect 51273 37417 51307 37451
rect 51307 37417 51316 37451
rect 51264 37408 51316 37417
rect 52092 37408 52144 37460
rect 56508 37408 56560 37460
rect 57796 37451 57848 37460
rect 57796 37417 57805 37451
rect 57805 37417 57839 37451
rect 57839 37417 57848 37451
rect 57796 37408 57848 37417
rect 59084 37408 59136 37460
rect 61844 37408 61896 37460
rect 64512 37408 64564 37460
rect 67180 37408 67232 37460
rect 69756 37408 69808 37460
rect 43352 37383 43404 37392
rect 43352 37349 43361 37383
rect 43361 37349 43395 37383
rect 43395 37349 43404 37383
rect 43352 37340 43404 37349
rect 47676 37340 47728 37392
rect 48504 37383 48556 37392
rect 48504 37349 48513 37383
rect 48513 37349 48547 37383
rect 48547 37349 48556 37383
rect 48504 37340 48556 37349
rect 49424 37340 49476 37392
rect 24124 37315 24176 37324
rect 24124 37281 24133 37315
rect 24133 37281 24167 37315
rect 24167 37281 24176 37315
rect 24124 37272 24176 37281
rect 26148 37272 26200 37324
rect 27160 37315 27212 37324
rect 27160 37281 27169 37315
rect 27169 37281 27203 37315
rect 27203 37281 27212 37315
rect 27160 37272 27212 37281
rect 28356 37315 28408 37324
rect 28356 37281 28365 37315
rect 28365 37281 28399 37315
rect 28399 37281 28408 37315
rect 28356 37272 28408 37281
rect 29644 37272 29696 37324
rect 31484 37272 31536 37324
rect 34060 37272 34112 37324
rect 36084 37272 36136 37324
rect 36636 37272 36688 37324
rect 37188 37315 37240 37324
rect 37188 37281 37197 37315
rect 37197 37281 37231 37315
rect 37231 37281 37240 37315
rect 37188 37272 37240 37281
rect 38660 37272 38712 37324
rect 39856 37315 39908 37324
rect 39856 37281 39865 37315
rect 39865 37281 39899 37315
rect 39899 37281 39908 37315
rect 39856 37272 39908 37281
rect 41696 37315 41748 37324
rect 41696 37281 41705 37315
rect 41705 37281 41739 37315
rect 41739 37281 41748 37315
rect 41696 37272 41748 37281
rect 42340 37272 42392 37324
rect 42892 37272 42944 37324
rect 44364 37315 44416 37324
rect 44364 37281 44373 37315
rect 44373 37281 44407 37315
rect 44407 37281 44416 37315
rect 44364 37272 44416 37281
rect 45100 37315 45152 37324
rect 45100 37281 45109 37315
rect 45109 37281 45143 37315
rect 45143 37281 45152 37315
rect 45100 37272 45152 37281
rect 47952 37272 48004 37324
rect 49700 37315 49752 37324
rect 49700 37281 49709 37315
rect 49709 37281 49743 37315
rect 49743 37281 49752 37315
rect 49700 37272 49752 37281
rect 49884 37315 49936 37324
rect 49884 37281 49893 37315
rect 49893 37281 49927 37315
rect 49927 37281 49936 37315
rect 49884 37272 49936 37281
rect 50160 37340 50212 37392
rect 53012 37340 53064 37392
rect 53840 37340 53892 37392
rect 55404 37340 55456 37392
rect 51172 37315 51224 37324
rect 51172 37281 51181 37315
rect 51181 37281 51215 37315
rect 51215 37281 51224 37315
rect 51172 37272 51224 37281
rect 52368 37315 52420 37324
rect 52368 37281 52377 37315
rect 52377 37281 52411 37315
rect 52411 37281 52420 37315
rect 52368 37272 52420 37281
rect 53472 37315 53524 37324
rect 53472 37281 53481 37315
rect 53481 37281 53515 37315
rect 53515 37281 53524 37315
rect 53472 37272 53524 37281
rect 54668 37272 54720 37324
rect 55680 37272 55732 37324
rect 58256 37340 58308 37392
rect 60832 37340 60884 37392
rect 61108 37383 61160 37392
rect 61108 37349 61117 37383
rect 61117 37349 61151 37383
rect 61151 37349 61160 37383
rect 61108 37340 61160 37349
rect 63500 37340 63552 37392
rect 63776 37383 63828 37392
rect 63776 37349 63785 37383
rect 63785 37349 63819 37383
rect 63819 37349 63828 37383
rect 63776 37340 63828 37349
rect 66168 37340 66220 37392
rect 66444 37383 66496 37392
rect 66444 37349 66453 37383
rect 66453 37349 66487 37383
rect 66487 37349 66496 37383
rect 66444 37340 66496 37349
rect 71412 37340 71464 37392
rect 77576 37408 77628 37460
rect 80152 37408 80204 37460
rect 81348 37408 81400 37460
rect 73988 37340 74040 37392
rect 58440 37315 58492 37324
rect 58440 37281 58449 37315
rect 58449 37281 58483 37315
rect 58483 37281 58492 37315
rect 58440 37272 58492 37281
rect 58900 37315 58952 37324
rect 58900 37281 58909 37315
rect 58909 37281 58943 37315
rect 58943 37281 58952 37315
rect 58900 37272 58952 37281
rect 61660 37315 61712 37324
rect 61660 37281 61669 37315
rect 61669 37281 61703 37315
rect 61703 37281 61712 37315
rect 61660 37272 61712 37281
rect 64328 37315 64380 37324
rect 64328 37281 64337 37315
rect 64337 37281 64371 37315
rect 64371 37281 64380 37315
rect 64328 37272 64380 37281
rect 66996 37315 67048 37324
rect 66996 37281 67005 37315
rect 67005 37281 67039 37315
rect 67039 37281 67048 37315
rect 66996 37272 67048 37281
rect 68744 37315 68796 37324
rect 68744 37281 68753 37315
rect 68753 37281 68787 37315
rect 68787 37281 68796 37315
rect 68744 37272 68796 37281
rect 22100 37204 22152 37256
rect 41052 37204 41104 37256
rect 64972 37204 65024 37256
rect 65064 37204 65116 37256
rect 68560 37204 68612 37256
rect 28540 37136 28592 37188
rect 68928 37179 68980 37188
rect 68928 37145 68937 37179
rect 68937 37145 68971 37179
rect 68971 37145 68980 37179
rect 68928 37136 68980 37145
rect 69480 37272 69532 37324
rect 71688 37272 71740 37324
rect 72332 37272 72384 37324
rect 76656 37340 76708 37392
rect 76840 37340 76892 37392
rect 81808 37340 81860 37392
rect 81900 37340 81952 37392
rect 82820 37408 82872 37460
rect 83648 37408 83700 37460
rect 85212 37383 85264 37392
rect 85212 37349 85221 37383
rect 85221 37349 85255 37383
rect 85255 37349 85264 37383
rect 85212 37340 85264 37349
rect 85396 37383 85448 37392
rect 85396 37349 85405 37383
rect 85405 37349 85439 37383
rect 85439 37349 85448 37383
rect 85396 37340 85448 37349
rect 85488 37340 85540 37392
rect 86316 37408 86368 37460
rect 74264 37315 74316 37324
rect 74264 37281 74273 37315
rect 74273 37281 74307 37315
rect 74307 37281 74316 37315
rect 74264 37272 74316 37281
rect 74724 37272 74776 37324
rect 74908 37272 74960 37324
rect 77484 37315 77536 37324
rect 70676 37204 70728 37256
rect 73252 37204 73304 37256
rect 73528 37204 73580 37256
rect 76196 37204 76248 37256
rect 76932 37247 76984 37256
rect 76932 37213 76941 37247
rect 76941 37213 76975 37247
rect 76975 37213 76984 37247
rect 76932 37204 76984 37213
rect 77484 37281 77493 37315
rect 77493 37281 77527 37315
rect 77527 37281 77536 37315
rect 77484 37272 77536 37281
rect 79048 37315 79100 37324
rect 79048 37281 79057 37315
rect 79057 37281 79091 37315
rect 79091 37281 79100 37315
rect 79048 37272 79100 37281
rect 80244 37315 80296 37324
rect 80244 37281 80253 37315
rect 80253 37281 80287 37315
rect 80287 37281 80296 37315
rect 80244 37272 80296 37281
rect 81440 37272 81492 37324
rect 82912 37315 82964 37324
rect 82912 37281 82921 37315
rect 82921 37281 82955 37315
rect 82955 37281 82964 37315
rect 82912 37272 82964 37281
rect 84200 37272 84252 37324
rect 87880 37383 87932 37392
rect 87880 37349 87889 37383
rect 87889 37349 87923 37383
rect 87923 37349 87932 37383
rect 87880 37340 87932 37349
rect 88064 37383 88116 37392
rect 88064 37349 88073 37383
rect 88073 37349 88107 37383
rect 88107 37349 88116 37383
rect 88064 37340 88116 37349
rect 89444 37383 89496 37392
rect 89444 37349 89453 37383
rect 89453 37349 89487 37383
rect 89487 37349 89496 37383
rect 89444 37340 89496 37349
rect 89720 37408 89772 37460
rect 95976 37408 96028 37460
rect 97632 37451 97684 37460
rect 97632 37417 97641 37451
rect 97641 37417 97675 37451
rect 97675 37417 97684 37451
rect 97632 37408 97684 37417
rect 90548 37383 90600 37392
rect 90548 37349 90557 37383
rect 90557 37349 90591 37383
rect 90591 37349 90600 37383
rect 90548 37340 90600 37349
rect 90732 37383 90784 37392
rect 90732 37349 90741 37383
rect 90741 37349 90775 37383
rect 90775 37349 90784 37383
rect 90732 37340 90784 37349
rect 93308 37383 93360 37392
rect 93308 37349 93317 37383
rect 93317 37349 93351 37383
rect 93351 37349 93360 37383
rect 93308 37340 93360 37349
rect 96068 37383 96120 37392
rect 96068 37349 96077 37383
rect 96077 37349 96111 37383
rect 96111 37349 96120 37383
rect 96068 37340 96120 37349
rect 93492 37315 93544 37324
rect 93492 37281 93501 37315
rect 93501 37281 93535 37315
rect 93535 37281 93544 37315
rect 93492 37272 93544 37281
rect 94136 37272 94188 37324
rect 95240 37315 95292 37324
rect 95240 37281 95249 37315
rect 95249 37281 95283 37315
rect 95283 37281 95292 37315
rect 95240 37272 95292 37281
rect 98552 37340 98604 37392
rect 3148 37111 3200 37120
rect 3148 37077 3157 37111
rect 3157 37077 3191 37111
rect 3191 37077 3200 37111
rect 3148 37068 3200 37077
rect 23480 37068 23532 37120
rect 29644 37068 29696 37120
rect 32864 37068 32916 37120
rect 40868 37068 40920 37120
rect 48320 37068 48372 37120
rect 48504 37068 48556 37120
rect 50712 37068 50764 37120
rect 65064 37068 65116 37120
rect 65156 37068 65208 37120
rect 70032 37068 70084 37120
rect 71504 37068 71556 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 65686 36966 65738 37018
rect 65750 36966 65802 37018
rect 65814 36966 65866 37018
rect 65878 36966 65930 37018
rect 96406 36966 96458 37018
rect 96470 36966 96522 37018
rect 96534 36966 96586 37018
rect 96598 36966 96650 37018
rect 2596 36864 2648 36916
rect 42064 36864 42116 36916
rect 42248 36864 42300 36916
rect 46940 36864 46992 36916
rect 2136 36839 2188 36848
rect 2136 36805 2145 36839
rect 2145 36805 2179 36839
rect 2179 36805 2188 36839
rect 2136 36796 2188 36805
rect 7380 36796 7432 36848
rect 9956 36796 10008 36848
rect 12624 36796 12676 36848
rect 15292 36796 15344 36848
rect 17868 36839 17920 36848
rect 17868 36805 17877 36839
rect 17877 36805 17911 36839
rect 17911 36805 17920 36839
rect 17868 36796 17920 36805
rect 19340 36796 19392 36848
rect 19524 36796 19576 36848
rect 20352 36796 20404 36848
rect 20720 36796 20772 36848
rect 24492 36796 24544 36848
rect 3240 36771 3292 36780
rect 3240 36737 3249 36771
rect 3249 36737 3283 36771
rect 3283 36737 3292 36771
rect 3240 36728 3292 36737
rect 23480 36728 23532 36780
rect 33692 36796 33744 36848
rect 36268 36796 36320 36848
rect 36636 36796 36688 36848
rect 53564 36864 53616 36916
rect 54760 36864 54812 36916
rect 55220 36864 55272 36916
rect 57336 36864 57388 36916
rect 60004 36864 60056 36916
rect 62580 36864 62632 36916
rect 65064 36864 65116 36916
rect 70492 36864 70544 36916
rect 70584 36864 70636 36916
rect 73160 36864 73212 36916
rect 73252 36864 73304 36916
rect 86960 36864 87012 36916
rect 2320 36703 2372 36712
rect 2320 36669 2329 36703
rect 2329 36669 2363 36703
rect 2363 36669 2372 36703
rect 2320 36660 2372 36669
rect 3516 36660 3568 36712
rect 8208 36703 8260 36712
rect 8208 36669 8217 36703
rect 8217 36669 8251 36703
rect 8251 36669 8260 36703
rect 8208 36660 8260 36669
rect 15476 36660 15528 36712
rect 7472 36635 7524 36644
rect 7472 36601 7481 36635
rect 7481 36601 7515 36635
rect 7515 36601 7524 36635
rect 7472 36592 7524 36601
rect 10324 36592 10376 36644
rect 17408 36592 17460 36644
rect 19524 36703 19576 36712
rect 19524 36669 19533 36703
rect 19533 36669 19567 36703
rect 19567 36669 19576 36703
rect 26700 36703 26752 36712
rect 19524 36660 19576 36669
rect 26700 36669 26709 36703
rect 26709 36669 26743 36703
rect 26743 36669 26752 36703
rect 26700 36660 26752 36669
rect 28632 36703 28684 36712
rect 28632 36669 28641 36703
rect 28641 36669 28675 36703
rect 28675 36669 28684 36703
rect 28632 36660 28684 36669
rect 29276 36660 29328 36712
rect 31668 36703 31720 36712
rect 31668 36669 31677 36703
rect 31677 36669 31711 36703
rect 31711 36669 31720 36703
rect 31668 36660 31720 36669
rect 36636 36660 36688 36712
rect 36728 36660 36780 36712
rect 39948 36660 40000 36712
rect 42432 36703 42484 36712
rect 42432 36669 42441 36703
rect 42441 36669 42475 36703
rect 42475 36669 42484 36703
rect 42432 36660 42484 36669
rect 8392 36567 8444 36576
rect 8392 36533 8401 36567
rect 8401 36533 8435 36567
rect 8435 36533 8444 36567
rect 8392 36524 8444 36533
rect 19064 36567 19116 36576
rect 19064 36533 19073 36567
rect 19073 36533 19107 36567
rect 19107 36533 19116 36567
rect 19064 36524 19116 36533
rect 20260 36592 20312 36644
rect 28264 36592 28316 36644
rect 29000 36635 29052 36644
rect 29000 36601 29009 36635
rect 29009 36601 29043 36635
rect 29043 36601 29052 36635
rect 29000 36592 29052 36601
rect 26700 36524 26752 36576
rect 27436 36524 27488 36576
rect 30288 36524 30340 36576
rect 33968 36592 34020 36644
rect 36268 36592 36320 36644
rect 42248 36592 42300 36644
rect 38108 36524 38160 36576
rect 43536 36703 43588 36712
rect 43536 36669 43545 36703
rect 43545 36669 43579 36703
rect 43579 36669 43588 36703
rect 43536 36660 43588 36669
rect 43812 36703 43864 36712
rect 43812 36669 43821 36703
rect 43821 36669 43855 36703
rect 43855 36669 43864 36703
rect 43812 36660 43864 36669
rect 88984 36796 89036 36848
rect 94228 36839 94280 36848
rect 94228 36805 94237 36839
rect 94237 36805 94271 36839
rect 94271 36805 94280 36839
rect 94228 36796 94280 36805
rect 96804 36839 96856 36848
rect 96804 36805 96813 36839
rect 96813 36805 96847 36839
rect 96847 36805 96856 36839
rect 96804 36796 96856 36805
rect 99472 36796 99524 36848
rect 47308 36728 47360 36780
rect 53472 36728 53524 36780
rect 53564 36728 53616 36780
rect 65156 36728 65208 36780
rect 47400 36660 47452 36712
rect 48228 36592 48280 36644
rect 48320 36592 48372 36644
rect 52920 36592 52972 36644
rect 54576 36592 54628 36644
rect 55588 36660 55640 36712
rect 67732 36728 67784 36780
rect 68192 36728 68244 36780
rect 93860 36728 93912 36780
rect 65432 36703 65484 36712
rect 65432 36669 65441 36703
rect 65441 36669 65475 36703
rect 65475 36669 65484 36703
rect 65432 36660 65484 36669
rect 67824 36660 67876 36712
rect 68468 36660 68520 36712
rect 70584 36703 70636 36712
rect 70584 36669 70593 36703
rect 70593 36669 70627 36703
rect 70627 36669 70636 36703
rect 70584 36660 70636 36669
rect 57428 36635 57480 36644
rect 45100 36567 45152 36576
rect 45100 36533 45109 36567
rect 45109 36533 45143 36567
rect 45143 36533 45152 36567
rect 45100 36524 45152 36533
rect 46664 36524 46716 36576
rect 52092 36524 52144 36576
rect 52184 36524 52236 36576
rect 57428 36601 57437 36635
rect 57437 36601 57471 36635
rect 57471 36601 57480 36635
rect 57428 36592 57480 36601
rect 60096 36635 60148 36644
rect 60096 36601 60105 36635
rect 60105 36601 60139 36635
rect 60139 36601 60148 36635
rect 60096 36592 60148 36601
rect 62672 36635 62724 36644
rect 62672 36601 62681 36635
rect 62681 36601 62715 36635
rect 62715 36601 62724 36635
rect 62672 36592 62724 36601
rect 55772 36524 55824 36576
rect 56324 36567 56376 36576
rect 56324 36533 56333 36567
rect 56333 36533 56367 36567
rect 56367 36533 56376 36567
rect 56324 36524 56376 36533
rect 56508 36524 56560 36576
rect 65616 36592 65668 36644
rect 65800 36635 65852 36644
rect 65800 36601 65809 36635
rect 65809 36601 65843 36635
rect 65843 36601 65852 36635
rect 65800 36592 65852 36601
rect 68008 36635 68060 36644
rect 68008 36601 68017 36635
rect 68017 36601 68051 36635
rect 68051 36601 68060 36635
rect 68008 36592 68060 36601
rect 68284 36592 68336 36644
rect 63040 36524 63092 36576
rect 65524 36524 65576 36576
rect 68468 36567 68520 36576
rect 68468 36533 68477 36567
rect 68477 36533 68511 36567
rect 68511 36533 68520 36567
rect 68468 36524 68520 36533
rect 68560 36524 68612 36576
rect 73988 36703 74040 36712
rect 73988 36669 73997 36703
rect 73997 36669 74031 36703
rect 74031 36669 74040 36703
rect 73988 36660 74040 36669
rect 75828 36660 75880 36712
rect 76196 36660 76248 36712
rect 78680 36703 78732 36712
rect 78680 36669 78689 36703
rect 78689 36669 78723 36703
rect 78723 36669 78732 36703
rect 78680 36660 78732 36669
rect 79324 36660 79376 36712
rect 84568 36660 84620 36712
rect 87144 36703 87196 36712
rect 87144 36669 87153 36703
rect 87153 36669 87187 36703
rect 87187 36669 87196 36703
rect 87144 36660 87196 36669
rect 89812 36660 89864 36712
rect 92480 36703 92532 36712
rect 92480 36669 92489 36703
rect 92489 36669 92523 36703
rect 92523 36669 92532 36703
rect 92480 36660 92532 36669
rect 72884 36635 72936 36644
rect 72884 36601 72893 36635
rect 72893 36601 72927 36635
rect 72927 36601 72936 36635
rect 72884 36592 72936 36601
rect 75920 36635 75972 36644
rect 72056 36524 72108 36576
rect 73436 36524 73488 36576
rect 73804 36524 73856 36576
rect 75920 36601 75929 36635
rect 75929 36601 75963 36635
rect 75963 36601 75972 36635
rect 75920 36592 75972 36601
rect 97632 36635 97684 36644
rect 79416 36524 79468 36576
rect 96620 36567 96672 36576
rect 96620 36533 96629 36567
rect 96629 36533 96663 36567
rect 96663 36533 96672 36567
rect 97632 36601 97641 36635
rect 97641 36601 97675 36635
rect 97675 36601 97684 36635
rect 97632 36592 97684 36601
rect 96620 36524 96672 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 50326 36422 50378 36474
rect 50390 36422 50442 36474
rect 50454 36422 50506 36474
rect 50518 36422 50570 36474
rect 81046 36422 81098 36474
rect 81110 36422 81162 36474
rect 81174 36422 81226 36474
rect 81238 36422 81290 36474
rect 4896 36184 4948 36236
rect 8300 36320 8352 36372
rect 8392 36320 8444 36372
rect 24768 36320 24820 36372
rect 24952 36320 25004 36372
rect 26792 36320 26844 36372
rect 6184 36184 6236 36236
rect 10968 36116 11020 36168
rect 12992 36227 13044 36236
rect 12992 36193 13001 36227
rect 13001 36193 13035 36227
rect 13035 36193 13044 36227
rect 12992 36184 13044 36193
rect 18696 36227 18748 36236
rect 18696 36193 18705 36227
rect 18705 36193 18739 36227
rect 18739 36193 18748 36227
rect 18696 36184 18748 36193
rect 27436 36227 27488 36236
rect 27436 36193 27445 36227
rect 27445 36193 27479 36227
rect 27479 36193 27488 36227
rect 27436 36184 27488 36193
rect 27804 36227 27856 36236
rect 27804 36193 27813 36227
rect 27813 36193 27847 36227
rect 27847 36193 27856 36227
rect 27804 36184 27856 36193
rect 28264 36252 28316 36304
rect 33416 36252 33468 36304
rect 34152 36252 34204 36304
rect 42156 36252 42208 36304
rect 42248 36252 42300 36304
rect 46940 36252 46992 36304
rect 33692 36184 33744 36236
rect 36728 36184 36780 36236
rect 37464 36184 37516 36236
rect 43352 36184 43404 36236
rect 43536 36184 43588 36236
rect 47768 36184 47820 36236
rect 48688 36184 48740 36236
rect 49608 36184 49660 36236
rect 52184 36227 52236 36236
rect 52184 36193 52193 36227
rect 52193 36193 52227 36227
rect 52227 36193 52236 36227
rect 52184 36184 52236 36193
rect 52368 36184 52420 36236
rect 54852 36227 54904 36236
rect 54852 36193 54861 36227
rect 54861 36193 54895 36227
rect 54895 36193 54904 36227
rect 54852 36184 54904 36193
rect 14096 36116 14148 36168
rect 22100 36116 22152 36168
rect 24308 36116 24360 36168
rect 28080 36159 28132 36168
rect 28080 36125 28089 36159
rect 28089 36125 28123 36159
rect 28123 36125 28132 36159
rect 28080 36116 28132 36125
rect 28724 36159 28776 36168
rect 28724 36125 28733 36159
rect 28733 36125 28767 36159
rect 28767 36125 28776 36159
rect 28724 36116 28776 36125
rect 31668 36116 31720 36168
rect 41420 36116 41472 36168
rect 41512 36116 41564 36168
rect 46940 36116 46992 36168
rect 47400 36116 47452 36168
rect 47584 36116 47636 36168
rect 51172 36116 51224 36168
rect 52276 36116 52328 36168
rect 52736 36159 52788 36168
rect 52736 36125 52745 36159
rect 52745 36125 52779 36159
rect 52779 36125 52788 36159
rect 52736 36116 52788 36125
rect 53012 36116 53064 36168
rect 55312 36184 55364 36236
rect 55496 36252 55548 36304
rect 55772 36320 55824 36372
rect 65432 36320 65484 36372
rect 65524 36320 65576 36372
rect 70492 36320 70544 36372
rect 70584 36320 70636 36372
rect 55864 36252 55916 36304
rect 59820 36252 59872 36304
rect 56600 36184 56652 36236
rect 72884 36252 72936 36304
rect 65340 36227 65392 36236
rect 65340 36193 65349 36227
rect 65349 36193 65383 36227
rect 65383 36193 65392 36227
rect 65340 36184 65392 36193
rect 55128 36159 55180 36168
rect 55128 36125 55137 36159
rect 55137 36125 55171 36159
rect 55171 36125 55180 36159
rect 55128 36116 55180 36125
rect 55588 36116 55640 36168
rect 55956 36116 56008 36168
rect 59360 36116 59412 36168
rect 63132 36159 63184 36168
rect 63132 36125 63141 36159
rect 63141 36125 63175 36159
rect 63175 36125 63184 36159
rect 63132 36116 63184 36125
rect 63408 36159 63460 36168
rect 63408 36125 63417 36159
rect 63417 36125 63451 36159
rect 63451 36125 63460 36159
rect 63408 36116 63460 36125
rect 64972 36116 65024 36168
rect 70216 36184 70268 36236
rect 70308 36184 70360 36236
rect 65616 36116 65668 36168
rect 76012 36320 76064 36372
rect 96620 36320 96672 36372
rect 81624 36184 81676 36236
rect 93860 36184 93912 36236
rect 94596 36184 94648 36236
rect 95056 36227 95108 36236
rect 95056 36193 95065 36227
rect 95065 36193 95099 36227
rect 95099 36193 95108 36227
rect 95056 36184 95108 36193
rect 97724 36184 97776 36236
rect 94044 36159 94096 36168
rect 94044 36125 94053 36159
rect 94053 36125 94087 36159
rect 94087 36125 94096 36159
rect 94044 36116 94096 36125
rect 6460 36023 6512 36032
rect 6460 35989 6469 36023
rect 6469 35989 6503 36023
rect 6503 35989 6512 36023
rect 6460 35980 6512 35989
rect 13912 35980 13964 36032
rect 35256 36048 35308 36100
rect 47124 36091 47176 36100
rect 33324 35980 33376 36032
rect 33416 35980 33468 36032
rect 43444 35980 43496 36032
rect 47124 36057 47133 36091
rect 47133 36057 47167 36091
rect 47167 36057 47176 36091
rect 47124 36048 47176 36057
rect 48412 36048 48464 36100
rect 55864 36048 55916 36100
rect 63040 36048 63092 36100
rect 65156 36048 65208 36100
rect 48596 35980 48648 36032
rect 55312 35980 55364 36032
rect 55588 35980 55640 36032
rect 64604 35980 64656 36032
rect 75920 36048 75972 36100
rect 66168 35980 66220 36032
rect 73528 35980 73580 36032
rect 73620 35980 73672 36032
rect 74172 36023 74224 36032
rect 74172 35989 74181 36023
rect 74181 35989 74215 36023
rect 74215 35989 74224 36023
rect 74172 35980 74224 35989
rect 74540 36023 74592 36032
rect 74540 35989 74549 36023
rect 74549 35989 74583 36023
rect 74583 35989 74592 36023
rect 74540 35980 74592 35989
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 65686 35878 65738 35930
rect 65750 35878 65802 35930
rect 65814 35878 65866 35930
rect 65878 35878 65930 35930
rect 96406 35878 96458 35930
rect 96470 35878 96522 35930
rect 96534 35878 96586 35930
rect 96598 35878 96650 35930
rect 24492 35819 24544 35828
rect 24492 35785 24501 35819
rect 24501 35785 24535 35819
rect 24535 35785 24544 35819
rect 24492 35776 24544 35785
rect 28632 35776 28684 35828
rect 33508 35776 33560 35828
rect 20168 35708 20220 35760
rect 43536 35776 43588 35828
rect 44180 35776 44232 35828
rect 48136 35776 48188 35828
rect 48228 35776 48280 35828
rect 51080 35776 51132 35828
rect 51172 35776 51224 35828
rect 57152 35776 57204 35828
rect 79140 35776 79192 35828
rect 91560 35776 91612 35828
rect 95240 35776 95292 35828
rect 33876 35708 33928 35760
rect 39028 35708 39080 35760
rect 46756 35708 46808 35760
rect 55588 35708 55640 35760
rect 11888 35640 11940 35692
rect 39488 35640 39540 35692
rect 39580 35683 39632 35692
rect 39580 35649 39589 35683
rect 39589 35649 39623 35683
rect 39623 35649 39632 35683
rect 39580 35640 39632 35649
rect 40040 35640 40092 35692
rect 43628 35640 43680 35692
rect 19156 35615 19208 35624
rect 19156 35581 19165 35615
rect 19165 35581 19199 35615
rect 19199 35581 19208 35615
rect 19156 35572 19208 35581
rect 24676 35615 24728 35624
rect 24676 35581 24685 35615
rect 24685 35581 24719 35615
rect 24719 35581 24728 35615
rect 24676 35572 24728 35581
rect 24768 35572 24820 35624
rect 25228 35615 25280 35624
rect 25228 35581 25237 35615
rect 25237 35581 25271 35615
rect 25271 35581 25280 35615
rect 25228 35572 25280 35581
rect 39304 35572 39356 35624
rect 39396 35572 39448 35624
rect 41144 35572 41196 35624
rect 45100 35640 45152 35692
rect 46572 35640 46624 35692
rect 47492 35640 47544 35692
rect 48320 35640 48372 35692
rect 49884 35640 49936 35692
rect 66996 35708 67048 35760
rect 67732 35708 67784 35760
rect 72700 35708 72752 35760
rect 43812 35572 43864 35624
rect 46112 35572 46164 35624
rect 46664 35572 46716 35624
rect 56692 35640 56744 35692
rect 88340 35708 88392 35760
rect 82360 35640 82412 35692
rect 51080 35572 51132 35624
rect 55496 35572 55548 35624
rect 55772 35572 55824 35624
rect 55956 35615 56008 35624
rect 55956 35581 55965 35615
rect 55965 35581 55999 35615
rect 55999 35581 56008 35615
rect 55956 35572 56008 35581
rect 56048 35572 56100 35624
rect 57152 35572 57204 35624
rect 61844 35572 61896 35624
rect 66720 35572 66772 35624
rect 66996 35572 67048 35624
rect 81900 35615 81952 35624
rect 12992 35504 13044 35556
rect 35992 35504 36044 35556
rect 36360 35504 36412 35556
rect 39672 35504 39724 35556
rect 41052 35504 41104 35556
rect 55312 35504 55364 35556
rect 29000 35436 29052 35488
rect 36452 35436 36504 35488
rect 36544 35436 36596 35488
rect 39396 35479 39448 35488
rect 39396 35445 39405 35479
rect 39405 35445 39439 35479
rect 39439 35445 39448 35479
rect 39396 35436 39448 35445
rect 40960 35479 41012 35488
rect 40960 35445 40969 35479
rect 40969 35445 41003 35479
rect 41003 35445 41012 35479
rect 40960 35436 41012 35445
rect 41328 35436 41380 35488
rect 43904 35436 43956 35488
rect 46388 35436 46440 35488
rect 65156 35504 65208 35556
rect 76012 35504 76064 35556
rect 81900 35581 81909 35615
rect 81909 35581 81943 35615
rect 81943 35581 81952 35615
rect 81900 35572 81952 35581
rect 81992 35572 82044 35624
rect 82176 35615 82228 35624
rect 82176 35581 82185 35615
rect 82185 35581 82219 35615
rect 82219 35581 82228 35615
rect 82176 35572 82228 35581
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 50326 35334 50378 35386
rect 50390 35334 50442 35386
rect 50454 35334 50506 35386
rect 50518 35334 50570 35386
rect 81046 35334 81098 35386
rect 81110 35334 81162 35386
rect 81174 35334 81226 35386
rect 81238 35334 81290 35386
rect 19156 35232 19208 35284
rect 46572 35232 46624 35284
rect 12164 35164 12216 35216
rect 24308 35164 24360 35216
rect 19984 35096 20036 35148
rect 23664 35096 23716 35148
rect 36360 35164 36412 35216
rect 36452 35164 36504 35216
rect 43352 35164 43404 35216
rect 43536 35207 43588 35216
rect 43536 35173 43545 35207
rect 43545 35173 43579 35207
rect 43579 35173 43588 35207
rect 43536 35164 43588 35173
rect 44272 35164 44324 35216
rect 56324 35232 56376 35284
rect 59360 35232 59412 35284
rect 96712 35232 96764 35284
rect 52184 35164 52236 35216
rect 52276 35164 52328 35216
rect 56692 35164 56744 35216
rect 56784 35164 56836 35216
rect 65984 35164 66036 35216
rect 36820 35139 36872 35148
rect 36820 35105 36829 35139
rect 36829 35105 36863 35139
rect 36863 35105 36872 35139
rect 36820 35096 36872 35105
rect 36912 35096 36964 35148
rect 41328 35096 41380 35148
rect 41420 35096 41472 35148
rect 42984 35096 43036 35148
rect 43720 35139 43772 35148
rect 43720 35105 43729 35139
rect 43729 35105 43763 35139
rect 43763 35105 43772 35139
rect 43904 35139 43956 35148
rect 43720 35096 43772 35105
rect 43904 35105 43913 35139
rect 43913 35105 43947 35139
rect 43947 35105 43956 35139
rect 43904 35096 43956 35105
rect 46756 35139 46808 35148
rect 46756 35105 46765 35139
rect 46765 35105 46799 35139
rect 46799 35105 46808 35139
rect 46756 35096 46808 35105
rect 47124 35139 47176 35148
rect 47124 35105 47138 35139
rect 47138 35105 47172 35139
rect 47172 35105 47176 35139
rect 47124 35096 47176 35105
rect 47308 35139 47360 35148
rect 47308 35105 47334 35139
rect 47334 35105 47360 35139
rect 47308 35096 47360 35105
rect 47492 35096 47544 35148
rect 52368 35096 52420 35148
rect 53932 35096 53984 35148
rect 55588 35096 55640 35148
rect 61844 35096 61896 35148
rect 62028 35139 62080 35148
rect 62028 35105 62037 35139
rect 62037 35105 62071 35139
rect 62071 35105 62080 35139
rect 62028 35096 62080 35105
rect 14464 35028 14516 35080
rect 62212 35028 62264 35080
rect 62580 35096 62632 35148
rect 64604 35096 64656 35148
rect 68100 35139 68152 35148
rect 68100 35105 68109 35139
rect 68109 35105 68143 35139
rect 68143 35105 68152 35139
rect 68100 35096 68152 35105
rect 68192 35096 68244 35148
rect 68836 35139 68888 35148
rect 68836 35105 68845 35139
rect 68845 35105 68879 35139
rect 68879 35105 68888 35139
rect 68836 35096 68888 35105
rect 70032 35096 70084 35148
rect 72332 35096 72384 35148
rect 78864 35139 78916 35148
rect 78864 35105 78873 35139
rect 78873 35105 78907 35139
rect 78907 35105 78916 35139
rect 78864 35096 78916 35105
rect 68744 35071 68796 35080
rect 68744 35037 68753 35071
rect 68753 35037 68787 35071
rect 68787 35037 68796 35071
rect 68744 35028 68796 35037
rect 68928 35028 68980 35080
rect 86316 35139 86368 35148
rect 86316 35105 86324 35139
rect 86324 35105 86358 35139
rect 86358 35105 86368 35139
rect 86316 35096 86368 35105
rect 94964 35096 95016 35148
rect 86408 35071 86460 35080
rect 86408 35037 86417 35071
rect 86417 35037 86451 35071
rect 86451 35037 86460 35071
rect 86408 35028 86460 35037
rect 95424 35071 95476 35080
rect 95424 35037 95433 35071
rect 95433 35037 95467 35071
rect 95467 35037 95476 35071
rect 95424 35028 95476 35037
rect 6736 34960 6788 35012
rect 21548 34960 21600 35012
rect 54116 34960 54168 35012
rect 54392 34935 54444 34944
rect 54392 34901 54401 34935
rect 54401 34901 54435 34935
rect 54435 34901 54444 34935
rect 54392 34892 54444 34901
rect 57152 34892 57204 34944
rect 59360 34892 59412 34944
rect 61844 34935 61896 34944
rect 61844 34901 61853 34935
rect 61853 34901 61887 34935
rect 61887 34901 61896 34935
rect 61844 34892 61896 34901
rect 63500 34892 63552 34944
rect 64236 34892 64288 34944
rect 76288 34892 76340 34944
rect 77208 34892 77260 34944
rect 86684 34960 86736 35012
rect 86868 34892 86920 34944
rect 95332 34935 95384 34944
rect 95332 34901 95341 34935
rect 95341 34901 95375 34935
rect 95375 34901 95384 34935
rect 95332 34892 95384 34901
rect 95516 34935 95568 34944
rect 95516 34901 95525 34935
rect 95525 34901 95559 34935
rect 95559 34901 95568 34935
rect 95516 34892 95568 34901
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 65686 34790 65738 34842
rect 65750 34790 65802 34842
rect 65814 34790 65866 34842
rect 65878 34790 65930 34842
rect 96406 34790 96458 34842
rect 96470 34790 96522 34842
rect 96534 34790 96586 34842
rect 96598 34790 96650 34842
rect 27988 34731 28040 34740
rect 27988 34697 27997 34731
rect 27997 34697 28031 34731
rect 28031 34697 28040 34731
rect 27988 34688 28040 34697
rect 31668 34688 31720 34740
rect 7564 34620 7616 34672
rect 36452 34620 36504 34672
rect 16120 34552 16172 34604
rect 36820 34688 36872 34740
rect 92112 34688 92164 34740
rect 40868 34620 40920 34672
rect 41512 34620 41564 34672
rect 43536 34620 43588 34672
rect 43628 34620 43680 34672
rect 49700 34620 49752 34672
rect 49792 34620 49844 34672
rect 50804 34620 50856 34672
rect 50988 34620 51040 34672
rect 53104 34620 53156 34672
rect 86868 34620 86920 34672
rect 19340 34484 19392 34536
rect 24400 34484 24452 34536
rect 25320 34484 25372 34536
rect 27804 34484 27856 34536
rect 18696 34416 18748 34468
rect 29000 34416 29052 34468
rect 29828 34484 29880 34536
rect 34152 34484 34204 34536
rect 34520 34527 34572 34536
rect 34520 34493 34529 34527
rect 34529 34493 34563 34527
rect 34563 34493 34572 34527
rect 34520 34484 34572 34493
rect 36912 34484 36964 34536
rect 37280 34484 37332 34536
rect 38200 34484 38252 34536
rect 39396 34527 39448 34536
rect 39396 34493 39405 34527
rect 39405 34493 39439 34527
rect 39439 34493 39448 34527
rect 39396 34484 39448 34493
rect 39488 34484 39540 34536
rect 39672 34527 39724 34536
rect 39672 34493 39695 34527
rect 39695 34493 39724 34527
rect 39672 34484 39724 34493
rect 39948 34484 40000 34536
rect 83464 34552 83516 34604
rect 87052 34552 87104 34604
rect 88892 34552 88944 34604
rect 40500 34484 40552 34536
rect 41512 34484 41564 34536
rect 43536 34484 43588 34536
rect 46848 34484 46900 34536
rect 46940 34484 46992 34536
rect 53104 34484 53156 34536
rect 54208 34484 54260 34536
rect 54852 34416 54904 34468
rect 55128 34416 55180 34468
rect 55312 34416 55364 34468
rect 58624 34416 58676 34468
rect 59360 34527 59412 34536
rect 59360 34493 59369 34527
rect 59369 34493 59403 34527
rect 59403 34493 59412 34527
rect 59360 34484 59412 34493
rect 59636 34484 59688 34536
rect 64972 34484 65024 34536
rect 65984 34484 66036 34536
rect 67088 34484 67140 34536
rect 67456 34527 67508 34536
rect 67456 34493 67465 34527
rect 67465 34493 67499 34527
rect 67499 34493 67508 34527
rect 67456 34484 67508 34493
rect 67548 34484 67600 34536
rect 68928 34484 68980 34536
rect 75184 34484 75236 34536
rect 75552 34484 75604 34536
rect 83280 34484 83332 34536
rect 94228 34527 94280 34536
rect 94228 34493 94237 34527
rect 94237 34493 94271 34527
rect 94271 34493 94280 34527
rect 94228 34484 94280 34493
rect 9956 34348 10008 34400
rect 27988 34348 28040 34400
rect 28080 34348 28132 34400
rect 33876 34348 33928 34400
rect 33968 34348 34020 34400
rect 41328 34348 41380 34400
rect 41696 34348 41748 34400
rect 52276 34348 52328 34400
rect 52368 34348 52420 34400
rect 88800 34416 88852 34468
rect 67456 34348 67508 34400
rect 69204 34348 69256 34400
rect 69296 34348 69348 34400
rect 90640 34348 90692 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 50326 34246 50378 34298
rect 50390 34246 50442 34298
rect 50454 34246 50506 34298
rect 50518 34246 50570 34298
rect 81046 34246 81098 34298
rect 81110 34246 81162 34298
rect 81174 34246 81226 34298
rect 81238 34246 81290 34298
rect 9956 34051 10008 34060
rect 9956 34017 9965 34051
rect 9965 34017 9999 34051
rect 9999 34017 10008 34051
rect 9956 34008 10008 34017
rect 28080 34144 28132 34196
rect 30472 34144 30524 34196
rect 31484 34144 31536 34196
rect 34796 34144 34848 34196
rect 35256 34144 35308 34196
rect 36360 34144 36412 34196
rect 22836 34076 22888 34128
rect 40500 34144 40552 34196
rect 40960 34144 41012 34196
rect 41420 34144 41472 34196
rect 41512 34144 41564 34196
rect 64788 34144 64840 34196
rect 64972 34144 65024 34196
rect 84844 34144 84896 34196
rect 85488 34144 85540 34196
rect 36544 34076 36596 34128
rect 46940 34076 46992 34128
rect 47308 34076 47360 34128
rect 18696 34051 18748 34060
rect 18236 33983 18288 33992
rect 9956 33872 10008 33924
rect 18236 33949 18245 33983
rect 18245 33949 18279 33983
rect 18279 33949 18288 33983
rect 18236 33940 18288 33949
rect 18696 34017 18705 34051
rect 18705 34017 18739 34051
rect 18739 34017 18748 34051
rect 18696 34008 18748 34017
rect 21640 34008 21692 34060
rect 24860 34008 24912 34060
rect 29368 34008 29420 34060
rect 30380 34008 30432 34060
rect 36452 34008 36504 34060
rect 36636 34008 36688 34060
rect 37832 34008 37884 34060
rect 38660 34008 38712 34060
rect 39948 34008 40000 34060
rect 40408 34008 40460 34060
rect 18880 33940 18932 33992
rect 21824 33983 21876 33992
rect 21824 33949 21833 33983
rect 21833 33949 21867 33983
rect 21867 33949 21876 33983
rect 21824 33940 21876 33949
rect 18512 33872 18564 33924
rect 33968 33940 34020 33992
rect 34152 33940 34204 33992
rect 42248 34051 42300 34060
rect 42248 34017 42257 34051
rect 42257 34017 42291 34051
rect 42291 34017 42300 34051
rect 42432 34051 42484 34060
rect 42248 34008 42300 34017
rect 42432 34017 42441 34051
rect 42441 34017 42475 34051
rect 42475 34017 42484 34051
rect 42432 34008 42484 34017
rect 42616 34008 42668 34060
rect 44272 34008 44324 34060
rect 50896 34008 50948 34060
rect 51172 34076 51224 34128
rect 58164 34076 58216 34128
rect 58624 34076 58676 34128
rect 68468 34008 68520 34060
rect 70676 34008 70728 34060
rect 77760 34051 77812 34060
rect 77760 34017 77769 34051
rect 77769 34017 77803 34051
rect 77803 34017 77812 34051
rect 77760 34008 77812 34017
rect 77852 34008 77904 34060
rect 95424 34008 95476 34060
rect 24768 33872 24820 33924
rect 36544 33872 36596 33924
rect 37740 33872 37792 33924
rect 41144 33872 41196 33924
rect 44456 33940 44508 33992
rect 45468 33940 45520 33992
rect 45560 33940 45612 33992
rect 50988 33940 51040 33992
rect 52276 33940 52328 33992
rect 61660 33940 61712 33992
rect 62028 33940 62080 33992
rect 64788 33940 64840 33992
rect 24584 33804 24636 33856
rect 53104 33872 53156 33924
rect 66904 33872 66956 33924
rect 70584 33940 70636 33992
rect 72424 33940 72476 33992
rect 72976 33872 73028 33924
rect 75552 33872 75604 33924
rect 55036 33804 55088 33856
rect 58072 33804 58124 33856
rect 59360 33804 59412 33856
rect 63224 33804 63276 33856
rect 63316 33804 63368 33856
rect 70768 33804 70820 33856
rect 93216 33847 93268 33856
rect 93216 33813 93225 33847
rect 93225 33813 93259 33847
rect 93259 33813 93268 33847
rect 95148 33940 95200 33992
rect 93216 33804 93268 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 65686 33702 65738 33754
rect 65750 33702 65802 33754
rect 65814 33702 65866 33754
rect 65878 33702 65930 33754
rect 96406 33702 96458 33754
rect 96470 33702 96522 33754
rect 96534 33702 96586 33754
rect 96598 33702 96650 33754
rect 17684 33600 17736 33652
rect 34152 33600 34204 33652
rect 34244 33600 34296 33652
rect 17592 33507 17644 33516
rect 17592 33473 17601 33507
rect 17601 33473 17635 33507
rect 17635 33473 17644 33507
rect 17592 33464 17644 33473
rect 19892 33464 19944 33516
rect 18880 33396 18932 33448
rect 19156 33396 19208 33448
rect 20996 33439 21048 33448
rect 20536 33328 20588 33380
rect 20996 33405 21005 33439
rect 21005 33405 21039 33439
rect 21039 33405 21048 33439
rect 20996 33396 21048 33405
rect 27804 33532 27856 33584
rect 30196 33532 30248 33584
rect 24492 33439 24544 33448
rect 24492 33405 24501 33439
rect 24501 33405 24535 33439
rect 24535 33405 24544 33439
rect 24492 33396 24544 33405
rect 30196 33439 30248 33448
rect 30196 33405 30205 33439
rect 30205 33405 30239 33439
rect 30239 33405 30248 33439
rect 30196 33396 30248 33405
rect 30288 33396 30340 33448
rect 30472 33439 30524 33448
rect 30472 33405 30477 33439
rect 30477 33405 30511 33439
rect 30511 33405 30524 33439
rect 30472 33396 30524 33405
rect 30932 33464 30984 33516
rect 40132 33532 40184 33584
rect 41144 33600 41196 33652
rect 67824 33600 67876 33652
rect 70124 33600 70176 33652
rect 70308 33600 70360 33652
rect 72240 33532 72292 33584
rect 21364 33328 21416 33380
rect 22100 33328 22152 33380
rect 25320 33328 25372 33380
rect 27988 33328 28040 33380
rect 28816 33328 28868 33380
rect 30012 33328 30064 33380
rect 36452 33396 36504 33448
rect 32496 33328 32548 33380
rect 40040 33396 40092 33448
rect 41328 33464 41380 33516
rect 45560 33464 45612 33516
rect 45652 33464 45704 33516
rect 49148 33464 49200 33516
rect 49056 33396 49108 33448
rect 54484 33464 54536 33516
rect 56140 33464 56192 33516
rect 60372 33464 60424 33516
rect 61384 33464 61436 33516
rect 62028 33464 62080 33516
rect 69296 33464 69348 33516
rect 53104 33396 53156 33448
rect 59360 33439 59412 33448
rect 18696 33303 18748 33312
rect 18696 33269 18705 33303
rect 18705 33269 18739 33303
rect 18739 33269 18748 33303
rect 18696 33260 18748 33269
rect 30472 33260 30524 33312
rect 30748 33303 30800 33312
rect 30748 33269 30757 33303
rect 30757 33269 30791 33303
rect 30791 33269 30800 33303
rect 30748 33260 30800 33269
rect 34796 33260 34848 33312
rect 37924 33260 37976 33312
rect 38016 33260 38068 33312
rect 41696 33328 41748 33380
rect 42708 33328 42760 33380
rect 49516 33371 49568 33380
rect 49516 33337 49525 33371
rect 49525 33337 49559 33371
rect 49559 33337 49568 33371
rect 49516 33328 49568 33337
rect 49608 33328 49660 33380
rect 51080 33328 51132 33380
rect 55312 33328 55364 33380
rect 58716 33328 58768 33380
rect 59360 33405 59369 33439
rect 59369 33405 59403 33439
rect 59403 33405 59412 33439
rect 59360 33396 59412 33405
rect 60280 33396 60332 33448
rect 60740 33439 60792 33448
rect 59452 33328 59504 33380
rect 59728 33371 59780 33380
rect 59728 33337 59737 33371
rect 59737 33337 59771 33371
rect 59771 33337 59780 33371
rect 59728 33328 59780 33337
rect 60372 33328 60424 33380
rect 60740 33405 60749 33439
rect 60749 33405 60783 33439
rect 60783 33405 60792 33439
rect 60740 33396 60792 33405
rect 60924 33396 60976 33448
rect 61292 33396 61344 33448
rect 84844 33396 84896 33448
rect 61476 33328 61528 33380
rect 60740 33260 60792 33312
rect 61108 33303 61160 33312
rect 61108 33269 61117 33303
rect 61117 33269 61151 33303
rect 61151 33269 61160 33303
rect 61108 33260 61160 33269
rect 63224 33260 63276 33312
rect 65984 33260 66036 33312
rect 83832 33260 83884 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 50326 33158 50378 33210
rect 50390 33158 50442 33210
rect 50454 33158 50506 33210
rect 50518 33158 50570 33210
rect 81046 33158 81098 33210
rect 81110 33158 81162 33210
rect 81174 33158 81226 33210
rect 81238 33158 81290 33210
rect 16764 33056 16816 33108
rect 90640 33099 90692 33108
rect 22192 32988 22244 33040
rect 38936 32988 38988 33040
rect 16672 32920 16724 32972
rect 22008 32920 22060 32972
rect 22376 32920 22428 32972
rect 16856 32852 16908 32904
rect 38292 32920 38344 32972
rect 38752 32920 38804 32972
rect 42156 32988 42208 33040
rect 42432 32988 42484 33040
rect 22652 32895 22704 32904
rect 22652 32861 22661 32895
rect 22661 32861 22695 32895
rect 22695 32861 22704 32895
rect 22652 32852 22704 32861
rect 26884 32852 26936 32904
rect 35440 32852 35492 32904
rect 38844 32852 38896 32904
rect 39488 32920 39540 32972
rect 42064 32963 42116 32972
rect 42064 32929 42073 32963
rect 42073 32929 42107 32963
rect 42107 32929 42116 32963
rect 42064 32920 42116 32929
rect 49332 32988 49384 33040
rect 71780 32988 71832 33040
rect 90640 33065 90649 33099
rect 90649 33065 90683 33099
rect 90683 33065 90692 33099
rect 90640 33056 90692 33065
rect 95516 32988 95568 33040
rect 39396 32895 39448 32904
rect 39396 32861 39405 32895
rect 39405 32861 39439 32895
rect 39439 32861 39448 32895
rect 39396 32852 39448 32861
rect 40500 32852 40552 32904
rect 13636 32759 13688 32768
rect 13636 32725 13645 32759
rect 13645 32725 13679 32759
rect 13679 32725 13688 32759
rect 13636 32716 13688 32725
rect 14004 32784 14056 32836
rect 21272 32784 21324 32836
rect 22376 32784 22428 32836
rect 26056 32784 26108 32836
rect 29368 32784 29420 32836
rect 39580 32784 39632 32836
rect 32404 32716 32456 32768
rect 32588 32716 32640 32768
rect 38660 32716 38712 32768
rect 38844 32759 38896 32768
rect 38844 32725 38853 32759
rect 38853 32725 38887 32759
rect 38887 32725 38896 32759
rect 38844 32716 38896 32725
rect 39948 32716 40000 32768
rect 42340 32784 42392 32836
rect 42800 32852 42852 32904
rect 47216 32895 47268 32904
rect 47216 32861 47225 32895
rect 47225 32861 47259 32895
rect 47259 32861 47268 32895
rect 47216 32852 47268 32861
rect 47308 32852 47360 32904
rect 49700 32852 49752 32904
rect 42708 32716 42760 32768
rect 43168 32716 43220 32768
rect 46572 32784 46624 32836
rect 50620 32784 50672 32836
rect 59728 32920 59780 32972
rect 90824 32920 90876 32972
rect 56048 32852 56100 32904
rect 60924 32852 60976 32904
rect 64328 32852 64380 32904
rect 68928 32852 68980 32904
rect 58532 32784 58584 32836
rect 59268 32784 59320 32836
rect 70584 32784 70636 32836
rect 61844 32716 61896 32768
rect 68836 32716 68888 32768
rect 69664 32716 69716 32768
rect 90088 32716 90140 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 65686 32614 65738 32666
rect 65750 32614 65802 32666
rect 65814 32614 65866 32666
rect 65878 32614 65930 32666
rect 96406 32614 96458 32666
rect 96470 32614 96522 32666
rect 96534 32614 96586 32666
rect 96598 32614 96650 32666
rect 13636 32512 13688 32564
rect 26884 32512 26936 32564
rect 26976 32512 27028 32564
rect 30380 32512 30432 32564
rect 31668 32512 31720 32564
rect 43168 32512 43220 32564
rect 55036 32512 55088 32564
rect 58164 32512 58216 32564
rect 85764 32512 85816 32564
rect 14004 32444 14056 32496
rect 23020 32487 23072 32496
rect 23020 32453 23029 32487
rect 23029 32453 23063 32487
rect 23063 32453 23072 32487
rect 23020 32444 23072 32453
rect 25412 32444 25464 32496
rect 39948 32444 40000 32496
rect 12256 32376 12308 32428
rect 21916 32376 21968 32428
rect 13820 32308 13872 32360
rect 14004 32308 14056 32360
rect 11612 32240 11664 32292
rect 22100 32308 22152 32360
rect 16028 32240 16080 32292
rect 22376 32240 22428 32292
rect 22468 32240 22520 32292
rect 17316 32172 17368 32224
rect 22284 32172 22336 32224
rect 41972 32376 42024 32428
rect 53748 32376 53800 32428
rect 27896 32351 27948 32360
rect 27896 32317 27905 32351
rect 27905 32317 27939 32351
rect 27939 32317 27948 32351
rect 27896 32308 27948 32317
rect 36636 32308 36688 32360
rect 39948 32308 40000 32360
rect 40040 32308 40092 32360
rect 40408 32351 40460 32360
rect 40408 32317 40417 32351
rect 40417 32317 40451 32351
rect 40451 32317 40460 32351
rect 40408 32308 40460 32317
rect 40684 32308 40736 32360
rect 55772 32351 55824 32360
rect 55772 32317 55781 32351
rect 55781 32317 55815 32351
rect 55815 32317 55824 32351
rect 55772 32308 55824 32317
rect 55864 32308 55916 32360
rect 56140 32351 56192 32360
rect 56140 32317 56149 32351
rect 56149 32317 56183 32351
rect 56183 32317 56192 32351
rect 56140 32308 56192 32317
rect 56416 32308 56468 32360
rect 56784 32444 56836 32496
rect 77852 32444 77904 32496
rect 58072 32376 58124 32428
rect 62856 32376 62908 32428
rect 78864 32308 78916 32360
rect 79692 32308 79744 32360
rect 84752 32308 84804 32360
rect 95056 32308 95108 32360
rect 29828 32240 29880 32292
rect 29920 32172 29972 32224
rect 33692 32240 33744 32292
rect 41788 32283 41840 32292
rect 33876 32172 33928 32224
rect 37004 32172 37056 32224
rect 41788 32249 41797 32283
rect 41797 32249 41831 32283
rect 41831 32249 41840 32283
rect 41788 32240 41840 32249
rect 56048 32240 56100 32292
rect 41972 32172 42024 32224
rect 42064 32172 42116 32224
rect 46572 32172 46624 32224
rect 47032 32172 47084 32224
rect 50988 32172 51040 32224
rect 51080 32172 51132 32224
rect 52368 32172 52420 32224
rect 53748 32172 53800 32224
rect 59728 32240 59780 32292
rect 68100 32240 68152 32292
rect 89168 32240 89220 32292
rect 87328 32172 87380 32224
rect 87788 32172 87840 32224
rect 95884 32172 95936 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 50326 32070 50378 32122
rect 50390 32070 50442 32122
rect 50454 32070 50506 32122
rect 50518 32070 50570 32122
rect 81046 32070 81098 32122
rect 81110 32070 81162 32122
rect 81174 32070 81226 32122
rect 81238 32070 81290 32122
rect 16028 31968 16080 32020
rect 13084 31875 13136 31884
rect 13084 31841 13093 31875
rect 13093 31841 13127 31875
rect 13127 31841 13136 31875
rect 13084 31832 13136 31841
rect 13268 31875 13320 31884
rect 13268 31841 13277 31875
rect 13277 31841 13311 31875
rect 13311 31841 13320 31875
rect 13268 31832 13320 31841
rect 13728 31900 13780 31952
rect 16764 31943 16816 31952
rect 16764 31909 16773 31943
rect 16773 31909 16807 31943
rect 16807 31909 16816 31943
rect 16764 31900 16816 31909
rect 17040 31900 17092 31952
rect 58072 31968 58124 32020
rect 58256 31968 58308 32020
rect 61016 31968 61068 32020
rect 88984 32011 89036 32020
rect 88984 31977 88993 32011
rect 88993 31977 89027 32011
rect 89027 31977 89036 32011
rect 88984 31968 89036 31977
rect 89536 31968 89588 32020
rect 90364 32011 90416 32020
rect 90364 31977 90373 32011
rect 90373 31977 90407 32011
rect 90407 31977 90416 32011
rect 90364 31968 90416 31977
rect 92572 31968 92624 32020
rect 12440 31764 12492 31816
rect 15200 31832 15252 31884
rect 41420 31900 41472 31952
rect 16856 31764 16908 31816
rect 17132 31807 17184 31816
rect 17132 31773 17141 31807
rect 17141 31773 17175 31807
rect 17175 31773 17184 31807
rect 17132 31764 17184 31773
rect 19064 31764 19116 31816
rect 27252 31832 27304 31884
rect 27712 31832 27764 31884
rect 22284 31764 22336 31816
rect 33692 31875 33744 31884
rect 33692 31841 33720 31875
rect 33720 31841 33744 31875
rect 33876 31875 33928 31884
rect 33692 31832 33744 31841
rect 33876 31841 33885 31875
rect 33885 31841 33919 31875
rect 33919 31841 33928 31875
rect 33876 31832 33928 31841
rect 33968 31875 34020 31884
rect 33968 31841 33977 31875
rect 33977 31841 34011 31875
rect 34011 31841 34020 31875
rect 33968 31832 34020 31841
rect 41328 31832 41380 31884
rect 51080 31900 51132 31952
rect 58808 31900 58860 31952
rect 84752 31900 84804 31952
rect 37188 31764 37240 31816
rect 17040 31739 17092 31748
rect 17040 31705 17049 31739
rect 17049 31705 17083 31739
rect 17083 31705 17092 31739
rect 17040 31696 17092 31705
rect 17224 31739 17276 31748
rect 17224 31705 17233 31739
rect 17233 31705 17267 31739
rect 17267 31705 17276 31739
rect 17224 31696 17276 31705
rect 17592 31696 17644 31748
rect 19340 31696 19392 31748
rect 22560 31696 22612 31748
rect 3608 31628 3660 31680
rect 24032 31628 24084 31680
rect 27528 31696 27580 31748
rect 33968 31628 34020 31680
rect 36268 31696 36320 31748
rect 37464 31696 37516 31748
rect 38292 31764 38344 31816
rect 40868 31764 40920 31816
rect 40500 31696 40552 31748
rect 41328 31696 41380 31748
rect 57888 31832 57940 31884
rect 57980 31875 58032 31884
rect 57980 31841 57988 31875
rect 57988 31841 58022 31875
rect 58022 31841 58032 31875
rect 57980 31832 58032 31841
rect 58164 31832 58216 31884
rect 58532 31832 58584 31884
rect 66812 31832 66864 31884
rect 69664 31832 69716 31884
rect 89168 31875 89220 31884
rect 89168 31841 89177 31875
rect 89177 31841 89211 31875
rect 89211 31841 89220 31875
rect 89168 31832 89220 31841
rect 44180 31764 44232 31816
rect 52828 31807 52880 31816
rect 41788 31696 41840 31748
rect 42892 31696 42944 31748
rect 44272 31696 44324 31748
rect 45836 31696 45888 31748
rect 50160 31696 50212 31748
rect 38844 31628 38896 31680
rect 39028 31628 39080 31680
rect 41144 31628 41196 31680
rect 43536 31628 43588 31680
rect 48412 31628 48464 31680
rect 52828 31773 52837 31807
rect 52837 31773 52871 31807
rect 52871 31773 52880 31807
rect 52828 31764 52880 31773
rect 53196 31764 53248 31816
rect 56232 31764 56284 31816
rect 54208 31739 54260 31748
rect 54208 31705 54217 31739
rect 54217 31705 54251 31739
rect 54251 31705 54260 31739
rect 54208 31696 54260 31705
rect 55036 31696 55088 31748
rect 57520 31696 57572 31748
rect 55680 31628 55732 31680
rect 56140 31628 56192 31680
rect 56232 31628 56284 31680
rect 58348 31696 58400 31748
rect 84200 31696 84252 31748
rect 58072 31628 58124 31680
rect 58808 31628 58860 31680
rect 60004 31628 60056 31680
rect 60280 31628 60332 31680
rect 60556 31628 60608 31680
rect 86592 31628 86644 31680
rect 89536 31875 89588 31884
rect 89536 31841 89545 31875
rect 89545 31841 89579 31875
rect 89579 31841 89588 31875
rect 89536 31832 89588 31841
rect 89812 31807 89864 31816
rect 89812 31773 89821 31807
rect 89821 31773 89855 31807
rect 89855 31773 89864 31807
rect 89812 31764 89864 31773
rect 92480 31832 92532 31884
rect 95884 31875 95936 31884
rect 95884 31841 95893 31875
rect 95893 31841 95927 31875
rect 95927 31841 95936 31875
rect 95884 31832 95936 31841
rect 90640 31764 90692 31816
rect 96068 31807 96120 31816
rect 93860 31696 93912 31748
rect 96068 31773 96077 31807
rect 96077 31773 96111 31807
rect 96111 31773 96120 31807
rect 96068 31764 96120 31773
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 65686 31526 65738 31578
rect 65750 31526 65802 31578
rect 65814 31526 65866 31578
rect 65878 31526 65930 31578
rect 96406 31526 96458 31578
rect 96470 31526 96522 31578
rect 96534 31526 96586 31578
rect 96598 31526 96650 31578
rect 3424 31424 3476 31476
rect 40960 31424 41012 31476
rect 44088 31424 44140 31476
rect 44272 31424 44324 31476
rect 51816 31424 51868 31476
rect 51908 31424 51960 31476
rect 17592 31399 17644 31408
rect 17592 31365 17601 31399
rect 17601 31365 17635 31399
rect 17635 31365 17644 31399
rect 17592 31356 17644 31365
rect 19340 31356 19392 31408
rect 19524 31356 19576 31408
rect 21272 31356 21324 31408
rect 27620 31356 27672 31408
rect 28080 31356 28132 31408
rect 28356 31356 28408 31408
rect 43536 31356 43588 31408
rect 43628 31356 43680 31408
rect 49332 31356 49384 31408
rect 49700 31356 49752 31408
rect 52644 31356 52696 31408
rect 52828 31356 52880 31408
rect 54116 31356 54168 31408
rect 54760 31356 54812 31408
rect 84200 31424 84252 31476
rect 94504 31424 94556 31476
rect 8944 31288 8996 31340
rect 18972 31288 19024 31340
rect 19156 31288 19208 31340
rect 9312 31220 9364 31272
rect 19432 31220 19484 31272
rect 19616 31288 19668 31340
rect 59728 31288 59780 31340
rect 54760 31263 54812 31272
rect 4896 31152 4948 31204
rect 19524 31195 19576 31204
rect 16856 31084 16908 31136
rect 19524 31161 19533 31195
rect 19533 31161 19567 31195
rect 19567 31161 19576 31195
rect 19524 31152 19576 31161
rect 20076 31152 20128 31204
rect 24308 31084 24360 31136
rect 24584 31084 24636 31136
rect 26516 31084 26568 31136
rect 27528 31084 27580 31136
rect 28172 31152 28224 31204
rect 43628 31152 43680 31204
rect 54760 31229 54769 31263
rect 54769 31229 54803 31263
rect 54803 31229 54812 31263
rect 54760 31220 54812 31229
rect 55036 31263 55088 31272
rect 55036 31229 55045 31263
rect 55045 31229 55079 31263
rect 55079 31229 55088 31263
rect 55036 31220 55088 31229
rect 55312 31220 55364 31272
rect 60280 31288 60332 31340
rect 60004 31220 60056 31272
rect 60648 31288 60700 31340
rect 93860 31288 93912 31340
rect 93952 31288 94004 31340
rect 53748 31084 53800 31136
rect 57520 31152 57572 31204
rect 55312 31084 55364 31136
rect 55680 31084 55732 31136
rect 56048 31084 56100 31136
rect 56232 31084 56284 31136
rect 60004 31127 60056 31136
rect 60004 31093 60013 31127
rect 60013 31093 60047 31127
rect 60047 31093 60056 31127
rect 60004 31084 60056 31093
rect 60188 31084 60240 31136
rect 60740 31263 60792 31272
rect 60740 31229 60749 31263
rect 60749 31229 60783 31263
rect 60783 31229 60792 31263
rect 60740 31220 60792 31229
rect 62028 31220 62080 31272
rect 87236 31263 87288 31272
rect 87236 31229 87245 31263
rect 87245 31229 87279 31263
rect 87279 31229 87288 31263
rect 87236 31220 87288 31229
rect 93400 31220 93452 31272
rect 91744 31152 91796 31204
rect 91836 31152 91888 31204
rect 93860 31152 93912 31204
rect 86684 31084 86736 31136
rect 87236 31084 87288 31136
rect 93584 31084 93636 31136
rect 94320 31195 94372 31204
rect 94320 31161 94329 31195
rect 94329 31161 94363 31195
rect 94363 31161 94372 31195
rect 94320 31152 94372 31161
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 50326 30982 50378 31034
rect 50390 30982 50442 31034
rect 50454 30982 50506 31034
rect 50518 30982 50570 31034
rect 81046 30982 81098 31034
rect 81110 30982 81162 31034
rect 81174 30982 81226 31034
rect 81238 30982 81290 31034
rect 10140 30880 10192 30932
rect 57520 30880 57572 30932
rect 59360 30880 59412 30932
rect 59912 30880 59964 30932
rect 60280 30880 60332 30932
rect 86040 30923 86092 30932
rect 19432 30812 19484 30864
rect 20812 30812 20864 30864
rect 28356 30812 28408 30864
rect 36636 30812 36688 30864
rect 37004 30812 37056 30864
rect 11152 30744 11204 30796
rect 11428 30744 11480 30796
rect 36544 30744 36596 30796
rect 37188 30744 37240 30796
rect 43996 30744 44048 30796
rect 46020 30744 46072 30796
rect 46664 30744 46716 30796
rect 16948 30676 17000 30728
rect 33876 30676 33928 30728
rect 33968 30676 34020 30728
rect 35348 30676 35400 30728
rect 36728 30676 36780 30728
rect 18512 30608 18564 30660
rect 45836 30608 45888 30660
rect 46296 30676 46348 30728
rect 46756 30719 46808 30728
rect 46756 30685 46765 30719
rect 46765 30685 46799 30719
rect 46799 30685 46808 30719
rect 46756 30676 46808 30685
rect 47032 30744 47084 30796
rect 47308 30676 47360 30728
rect 53656 30744 53708 30796
rect 53748 30744 53800 30796
rect 60004 30744 60056 30796
rect 61108 30812 61160 30864
rect 67548 30812 67600 30864
rect 72056 30812 72108 30864
rect 70676 30744 70728 30796
rect 71688 30744 71740 30796
rect 72424 30787 72476 30796
rect 72424 30753 72433 30787
rect 72433 30753 72467 30787
rect 72467 30753 72476 30787
rect 72424 30744 72476 30753
rect 75460 30812 75512 30864
rect 86040 30889 86049 30923
rect 86049 30889 86083 30923
rect 86083 30889 86092 30923
rect 86040 30880 86092 30889
rect 86316 30812 86368 30864
rect 72792 30787 72844 30796
rect 72792 30753 72801 30787
rect 72801 30753 72835 30787
rect 72835 30753 72844 30787
rect 72792 30744 72844 30753
rect 73068 30744 73120 30796
rect 51080 30676 51132 30728
rect 58808 30676 58860 30728
rect 47584 30608 47636 30660
rect 55220 30608 55272 30660
rect 59360 30676 59412 30728
rect 59636 30676 59688 30728
rect 60556 30676 60608 30728
rect 63224 30676 63276 30728
rect 86592 30787 86644 30796
rect 86592 30753 86606 30787
rect 86606 30753 86640 30787
rect 86640 30753 86644 30787
rect 86592 30744 86644 30753
rect 14004 30540 14056 30592
rect 14188 30540 14240 30592
rect 17132 30540 17184 30592
rect 18788 30540 18840 30592
rect 45100 30540 45152 30592
rect 47032 30540 47084 30592
rect 47216 30540 47268 30592
rect 49148 30540 49200 30592
rect 51816 30540 51868 30592
rect 59084 30608 59136 30660
rect 72056 30608 72108 30660
rect 55496 30540 55548 30592
rect 62488 30540 62540 30592
rect 63224 30540 63276 30592
rect 66904 30540 66956 30592
rect 69480 30540 69532 30592
rect 74448 30540 74500 30592
rect 86776 30583 86828 30592
rect 86776 30549 86785 30583
rect 86785 30549 86819 30583
rect 86819 30549 86828 30583
rect 86776 30540 86828 30549
rect 88616 30583 88668 30592
rect 88616 30549 88625 30583
rect 88625 30549 88659 30583
rect 88659 30549 88668 30583
rect 88616 30540 88668 30549
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 65686 30438 65738 30490
rect 65750 30438 65802 30490
rect 65814 30438 65866 30490
rect 65878 30438 65930 30490
rect 96406 30438 96458 30490
rect 96470 30438 96522 30490
rect 96534 30438 96586 30490
rect 96598 30438 96650 30490
rect 8300 30336 8352 30388
rect 9312 30336 9364 30388
rect 10324 30336 10376 30388
rect 25228 30336 25280 30388
rect 30288 30336 30340 30388
rect 30380 30336 30432 30388
rect 69112 30336 69164 30388
rect 70216 30336 70268 30388
rect 71320 30336 71372 30388
rect 17132 30268 17184 30320
rect 54208 30268 54260 30320
rect 55128 30268 55180 30320
rect 59544 30268 59596 30320
rect 6092 30200 6144 30252
rect 10140 30243 10192 30252
rect 10140 30209 10149 30243
rect 10149 30209 10183 30243
rect 10183 30209 10192 30243
rect 10140 30200 10192 30209
rect 10784 30200 10836 30252
rect 14004 30200 14056 30252
rect 37648 30200 37700 30252
rect 43720 30200 43772 30252
rect 65616 30268 65668 30320
rect 73620 30268 73672 30320
rect 71044 30200 71096 30252
rect 10876 30132 10928 30184
rect 12072 30175 12124 30184
rect 12072 30141 12081 30175
rect 12081 30141 12115 30175
rect 12115 30141 12124 30175
rect 12072 30132 12124 30141
rect 17224 30132 17276 30184
rect 17868 30132 17920 30184
rect 33232 30132 33284 30184
rect 54668 30132 54720 30184
rect 15476 30064 15528 30116
rect 24676 30107 24728 30116
rect 24676 30073 24685 30107
rect 24685 30073 24719 30107
rect 24719 30073 24728 30107
rect 24676 30064 24728 30073
rect 25964 30064 26016 30116
rect 30380 30064 30432 30116
rect 35624 30064 35676 30116
rect 36360 30064 36412 30116
rect 40040 30064 40092 30116
rect 40684 30064 40736 30116
rect 42984 30064 43036 30116
rect 43444 30064 43496 30116
rect 55128 30132 55180 30184
rect 55220 30132 55272 30184
rect 12072 29996 12124 30048
rect 15844 29996 15896 30048
rect 17224 29996 17276 30048
rect 55036 30064 55088 30116
rect 58072 30064 58124 30116
rect 62764 30132 62816 30184
rect 68468 30132 68520 30184
rect 68560 30132 68612 30184
rect 71320 30132 71372 30184
rect 80520 30175 80572 30184
rect 45284 29996 45336 30048
rect 47216 29996 47268 30048
rect 47308 29996 47360 30048
rect 48136 29996 48188 30048
rect 49332 29996 49384 30048
rect 55680 29996 55732 30048
rect 60004 29996 60056 30048
rect 79876 30064 79928 30116
rect 62028 29996 62080 30048
rect 68284 29996 68336 30048
rect 70768 29996 70820 30048
rect 73988 29996 74040 30048
rect 80520 30141 80529 30175
rect 80529 30141 80563 30175
rect 80563 30141 80572 30175
rect 80520 30132 80572 30141
rect 86224 30132 86276 30184
rect 89628 30132 89680 30184
rect 94688 30200 94740 30252
rect 95148 30200 95200 30252
rect 93308 30132 93360 30184
rect 81624 30064 81676 30116
rect 81900 30107 81952 30116
rect 81900 30073 81909 30107
rect 81909 30073 81943 30107
rect 81943 30073 81952 30107
rect 81900 30064 81952 30073
rect 92664 30107 92716 30116
rect 92664 30073 92673 30107
rect 92673 30073 92707 30107
rect 92707 30073 92716 30107
rect 92664 30064 92716 30073
rect 80888 29996 80940 30048
rect 84476 29996 84528 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 50326 29894 50378 29946
rect 50390 29894 50442 29946
rect 50454 29894 50506 29946
rect 50518 29894 50570 29946
rect 81046 29894 81098 29946
rect 81110 29894 81162 29946
rect 81174 29894 81226 29946
rect 81238 29894 81290 29946
rect 15476 29792 15528 29844
rect 16396 29792 16448 29844
rect 43352 29792 43404 29844
rect 13452 29724 13504 29776
rect 26148 29656 26200 29708
rect 38292 29724 38344 29776
rect 39120 29767 39172 29776
rect 39120 29733 39129 29767
rect 39129 29733 39163 29767
rect 39163 29733 39172 29767
rect 39120 29724 39172 29733
rect 43168 29724 43220 29776
rect 45652 29724 45704 29776
rect 34428 29588 34480 29640
rect 35532 29588 35584 29640
rect 38292 29631 38344 29640
rect 2504 29563 2556 29572
rect 2504 29529 2513 29563
rect 2513 29529 2547 29563
rect 2547 29529 2556 29563
rect 2504 29520 2556 29529
rect 6460 29520 6512 29572
rect 35716 29520 35768 29572
rect 36360 29520 36412 29572
rect 15200 29452 15252 29504
rect 18972 29452 19024 29504
rect 22192 29452 22244 29504
rect 27712 29452 27764 29504
rect 29828 29452 29880 29504
rect 30656 29452 30708 29504
rect 37188 29495 37240 29504
rect 37188 29461 37197 29495
rect 37197 29461 37231 29495
rect 37231 29461 37240 29495
rect 37188 29452 37240 29461
rect 38292 29597 38301 29631
rect 38301 29597 38335 29631
rect 38335 29597 38344 29631
rect 38292 29588 38344 29597
rect 45744 29656 45796 29708
rect 46572 29792 46624 29844
rect 46940 29792 46992 29844
rect 55036 29792 55088 29844
rect 46664 29767 46716 29776
rect 46664 29733 46673 29767
rect 46673 29733 46707 29767
rect 46707 29733 46716 29767
rect 46664 29724 46716 29733
rect 47216 29724 47268 29776
rect 65432 29792 65484 29844
rect 61384 29724 61436 29776
rect 62028 29724 62080 29776
rect 68284 29792 68336 29844
rect 92204 29792 92256 29844
rect 70768 29724 70820 29776
rect 88340 29767 88392 29776
rect 88340 29733 88349 29767
rect 88349 29733 88383 29767
rect 88383 29733 88392 29767
rect 88340 29724 88392 29733
rect 40132 29588 40184 29640
rect 46204 29588 46256 29640
rect 46664 29588 46716 29640
rect 46940 29656 46992 29708
rect 47308 29588 47360 29640
rect 38476 29520 38528 29572
rect 38568 29520 38620 29572
rect 43352 29520 43404 29572
rect 45836 29520 45888 29572
rect 48780 29588 48832 29640
rect 55496 29588 55548 29640
rect 55680 29588 55732 29640
rect 66536 29588 66588 29640
rect 67180 29631 67232 29640
rect 67180 29597 67189 29631
rect 67189 29597 67223 29631
rect 67223 29597 67232 29631
rect 67180 29588 67232 29597
rect 67456 29631 67508 29640
rect 67456 29597 67465 29631
rect 67465 29597 67499 29631
rect 67499 29597 67508 29631
rect 67456 29588 67508 29597
rect 67548 29588 67600 29640
rect 68560 29588 68612 29640
rect 68652 29588 68704 29640
rect 61016 29520 61068 29572
rect 68928 29588 68980 29640
rect 84476 29588 84528 29640
rect 39948 29452 40000 29504
rect 41604 29452 41656 29504
rect 42616 29452 42668 29504
rect 46664 29452 46716 29504
rect 47216 29452 47268 29504
rect 68560 29495 68612 29504
rect 68560 29461 68569 29495
rect 68569 29461 68603 29495
rect 68603 29461 68612 29495
rect 68560 29452 68612 29461
rect 82912 29520 82964 29572
rect 84108 29520 84160 29572
rect 88708 29520 88760 29572
rect 89628 29452 89680 29504
rect 94044 29588 94096 29640
rect 95148 29588 95200 29640
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 65686 29350 65738 29402
rect 65750 29350 65802 29402
rect 65814 29350 65866 29402
rect 65878 29350 65930 29402
rect 96406 29350 96458 29402
rect 96470 29350 96522 29402
rect 96534 29350 96586 29402
rect 96598 29350 96650 29402
rect 17132 29248 17184 29300
rect 15844 29180 15896 29232
rect 19064 29248 19116 29300
rect 21824 29248 21876 29300
rect 71044 29248 71096 29300
rect 26148 29223 26200 29232
rect 17224 29112 17276 29164
rect 3516 29044 3568 29096
rect 9404 29044 9456 29096
rect 12072 29044 12124 29096
rect 14004 29087 14056 29096
rect 14004 29053 14013 29087
rect 14013 29053 14047 29087
rect 14047 29053 14056 29087
rect 14004 29044 14056 29053
rect 15568 29087 15620 29096
rect 15568 29053 15577 29087
rect 15577 29053 15611 29087
rect 15611 29053 15620 29087
rect 15568 29044 15620 29053
rect 26148 29189 26157 29223
rect 26157 29189 26191 29223
rect 26191 29189 26200 29223
rect 26148 29180 26200 29189
rect 26332 29180 26384 29232
rect 27160 29180 27212 29232
rect 37004 29223 37056 29232
rect 37004 29189 37013 29223
rect 37013 29189 37047 29223
rect 37047 29189 37056 29223
rect 37004 29180 37056 29189
rect 37188 29180 37240 29232
rect 42064 29180 42116 29232
rect 42800 29180 42852 29232
rect 46204 29180 46256 29232
rect 46940 29180 46992 29232
rect 53748 29180 53800 29232
rect 56508 29180 56560 29232
rect 57152 29180 57204 29232
rect 57336 29180 57388 29232
rect 57520 29180 57572 29232
rect 65432 29180 65484 29232
rect 67824 29180 67876 29232
rect 68652 29180 68704 29232
rect 68836 29180 68888 29232
rect 83924 29180 83976 29232
rect 84108 29180 84160 29232
rect 86224 29180 86276 29232
rect 95884 29248 95936 29300
rect 24308 29112 24360 29164
rect 24768 29112 24820 29164
rect 24216 29087 24268 29096
rect 24216 29053 24225 29087
rect 24225 29053 24259 29087
rect 24259 29053 24268 29087
rect 24216 29044 24268 29053
rect 26608 29044 26660 29096
rect 33416 29044 33468 29096
rect 35624 29087 35676 29096
rect 35624 29053 35633 29087
rect 35633 29053 35667 29087
rect 35667 29053 35676 29087
rect 35624 29044 35676 29053
rect 38108 29044 38160 29096
rect 38292 29044 38344 29096
rect 38476 29044 38528 29096
rect 14556 29019 14608 29028
rect 14556 28985 14565 29019
rect 14565 28985 14599 29019
rect 14599 28985 14608 29019
rect 14556 28976 14608 28985
rect 9036 28908 9088 28960
rect 36728 28976 36780 29028
rect 45836 29044 45888 29096
rect 79048 29112 79100 29164
rect 86960 29155 87012 29164
rect 86960 29121 86969 29155
rect 86969 29121 87003 29155
rect 87003 29121 87012 29155
rect 86960 29112 87012 29121
rect 88708 29112 88760 29164
rect 46112 28976 46164 29028
rect 46204 28976 46256 29028
rect 55312 28976 55364 29028
rect 55496 28976 55548 29028
rect 67916 28976 67968 29028
rect 53840 28908 53892 28960
rect 55680 28908 55732 28960
rect 59636 28908 59688 28960
rect 59728 28908 59780 28960
rect 63040 28908 63092 28960
rect 63132 28908 63184 28960
rect 67180 28908 67232 28960
rect 68468 29087 68520 29096
rect 68468 29053 68477 29087
rect 68477 29053 68511 29087
rect 68511 29053 68520 29087
rect 68468 29044 68520 29053
rect 68652 29087 68704 29096
rect 68652 29053 68662 29087
rect 68662 29053 68696 29087
rect 68696 29053 68704 29087
rect 68652 29044 68704 29053
rect 68928 29044 68980 29096
rect 71136 29044 71188 29096
rect 73988 29044 74040 29096
rect 86592 29044 86644 29096
rect 69388 28976 69440 29028
rect 79600 28976 79652 29028
rect 98092 29019 98144 29028
rect 68284 28908 68336 28960
rect 71044 28951 71096 28960
rect 71044 28917 71053 28951
rect 71053 28917 71087 28951
rect 71087 28917 71096 28951
rect 71044 28908 71096 28917
rect 74724 28908 74776 28960
rect 98092 28985 98101 29019
rect 98101 28985 98135 29019
rect 98135 28985 98144 29019
rect 98092 28976 98144 28985
rect 92664 28908 92716 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 50326 28806 50378 28858
rect 50390 28806 50442 28858
rect 50454 28806 50506 28858
rect 50518 28806 50570 28858
rect 81046 28806 81098 28858
rect 81110 28806 81162 28858
rect 81174 28806 81226 28858
rect 81238 28806 81290 28858
rect 4068 28704 4120 28756
rect 22560 28704 22612 28756
rect 26792 28704 26844 28756
rect 28080 28704 28132 28756
rect 3516 28568 3568 28620
rect 6736 28568 6788 28620
rect 15660 28611 15712 28620
rect 15660 28577 15669 28611
rect 15669 28577 15703 28611
rect 15703 28577 15712 28611
rect 15660 28568 15712 28577
rect 17040 28568 17092 28620
rect 20536 28568 20588 28620
rect 20812 28611 20864 28620
rect 20812 28577 20821 28611
rect 20821 28577 20855 28611
rect 20855 28577 20864 28611
rect 20812 28568 20864 28577
rect 5356 28364 5408 28416
rect 6000 28364 6052 28416
rect 16580 28500 16632 28552
rect 16764 28500 16816 28552
rect 20996 28500 21048 28552
rect 26240 28500 26292 28552
rect 14280 28432 14332 28484
rect 15108 28364 15160 28416
rect 22100 28432 22152 28484
rect 23388 28432 23440 28484
rect 37372 28747 37424 28756
rect 37372 28713 37381 28747
rect 37381 28713 37415 28747
rect 37415 28713 37424 28747
rect 37372 28704 37424 28713
rect 46204 28704 46256 28756
rect 47032 28704 47084 28756
rect 37740 28679 37792 28688
rect 33508 28611 33560 28620
rect 33508 28577 33517 28611
rect 33517 28577 33551 28611
rect 33551 28577 33560 28611
rect 33508 28568 33560 28577
rect 37740 28645 37749 28679
rect 37749 28645 37783 28679
rect 37783 28645 37792 28679
rect 37740 28636 37792 28645
rect 39672 28636 39724 28688
rect 48044 28636 48096 28688
rect 52368 28704 52420 28756
rect 97908 28704 97960 28756
rect 27160 28500 27212 28552
rect 37004 28568 37056 28620
rect 37280 28611 37332 28620
rect 37280 28577 37289 28611
rect 37289 28577 37323 28611
rect 37323 28577 37332 28611
rect 37280 28568 37332 28577
rect 37556 28611 37608 28620
rect 37556 28577 37565 28611
rect 37565 28577 37599 28611
rect 37599 28577 37608 28611
rect 37556 28568 37608 28577
rect 55680 28568 55732 28620
rect 37740 28500 37792 28552
rect 42432 28500 42484 28552
rect 42524 28500 42576 28552
rect 46296 28500 46348 28552
rect 31760 28432 31812 28484
rect 17224 28407 17276 28416
rect 17224 28373 17233 28407
rect 17233 28373 17267 28407
rect 17267 28373 17276 28407
rect 17224 28364 17276 28373
rect 17776 28407 17828 28416
rect 17776 28373 17785 28407
rect 17785 28373 17819 28407
rect 17819 28373 17828 28407
rect 17776 28364 17828 28373
rect 18788 28364 18840 28416
rect 19248 28364 19300 28416
rect 19892 28364 19944 28416
rect 20168 28364 20220 28416
rect 20536 28364 20588 28416
rect 27160 28364 27212 28416
rect 30288 28364 30340 28416
rect 33876 28407 33928 28416
rect 33876 28373 33885 28407
rect 33885 28373 33919 28407
rect 33919 28373 33928 28407
rect 33876 28364 33928 28373
rect 37004 28407 37056 28416
rect 37004 28373 37013 28407
rect 37013 28373 37047 28407
rect 37047 28373 37056 28407
rect 37004 28364 37056 28373
rect 38292 28364 38344 28416
rect 49424 28543 49476 28552
rect 49424 28509 49433 28543
rect 49433 28509 49467 28543
rect 49467 28509 49476 28543
rect 49424 28500 49476 28509
rect 49792 28500 49844 28552
rect 52460 28500 52512 28552
rect 53656 28500 53708 28552
rect 53840 28500 53892 28552
rect 60372 28636 60424 28688
rect 56324 28568 56376 28620
rect 61936 28568 61988 28620
rect 61844 28500 61896 28552
rect 71044 28636 71096 28688
rect 62672 28568 62724 28620
rect 78956 28611 79008 28620
rect 49516 28432 49568 28484
rect 56324 28432 56376 28484
rect 56968 28432 57020 28484
rect 59728 28432 59780 28484
rect 48044 28364 48096 28416
rect 63132 28364 63184 28416
rect 63224 28364 63276 28416
rect 69480 28364 69532 28416
rect 78956 28577 78965 28611
rect 78965 28577 78999 28611
rect 78999 28577 79008 28611
rect 78956 28568 79008 28577
rect 78404 28432 78456 28484
rect 78680 28432 78732 28484
rect 79048 28432 79100 28484
rect 94780 28432 94832 28484
rect 80888 28407 80940 28416
rect 80888 28373 80897 28407
rect 80897 28373 80931 28407
rect 80931 28373 80940 28407
rect 80888 28364 80940 28373
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 65686 28262 65738 28314
rect 65750 28262 65802 28314
rect 65814 28262 65866 28314
rect 65878 28262 65930 28314
rect 96406 28262 96458 28314
rect 96470 28262 96522 28314
rect 96534 28262 96586 28314
rect 96598 28262 96650 28314
rect 3608 28203 3660 28212
rect 3608 28169 3617 28203
rect 3617 28169 3651 28203
rect 3651 28169 3660 28203
rect 3608 28160 3660 28169
rect 3792 28160 3844 28212
rect 14280 28160 14332 28212
rect 14464 28203 14516 28212
rect 14464 28169 14473 28203
rect 14473 28169 14507 28203
rect 14507 28169 14516 28203
rect 14464 28160 14516 28169
rect 2504 28092 2556 28144
rect 5356 28092 5408 28144
rect 13820 28092 13872 28144
rect 16580 28092 16632 28144
rect 17776 28092 17828 28144
rect 19892 28092 19944 28144
rect 20076 28135 20128 28144
rect 20076 28101 20085 28135
rect 20085 28101 20119 28135
rect 20119 28101 20128 28135
rect 20076 28092 20128 28101
rect 23388 28160 23440 28212
rect 30012 28160 30064 28212
rect 30380 28160 30432 28212
rect 38292 28160 38344 28212
rect 49516 28160 49568 28212
rect 49700 28160 49752 28212
rect 88616 28160 88668 28212
rect 39304 28092 39356 28144
rect 39396 28092 39448 28144
rect 46204 28092 46256 28144
rect 46296 28092 46348 28144
rect 49792 28092 49844 28144
rect 49976 28092 50028 28144
rect 62948 28092 63000 28144
rect 63040 28092 63092 28144
rect 68376 28092 68428 28144
rect 68928 28092 68980 28144
rect 17408 28067 17460 28076
rect 3792 27999 3844 28008
rect 3792 27965 3801 27999
rect 3801 27965 3835 27999
rect 3835 27965 3844 27999
rect 3792 27956 3844 27965
rect 4068 27999 4120 28008
rect 4068 27965 4077 27999
rect 4077 27965 4111 27999
rect 4111 27965 4120 27999
rect 4068 27956 4120 27965
rect 11796 27956 11848 28008
rect 14004 27931 14056 27940
rect 14004 27897 14013 27931
rect 14013 27897 14047 27931
rect 14047 27897 14056 27931
rect 14004 27888 14056 27897
rect 3976 27863 4028 27872
rect 3976 27829 3985 27863
rect 3985 27829 4019 27863
rect 4019 27829 4028 27863
rect 3976 27820 4028 27829
rect 14096 27863 14148 27872
rect 14096 27829 14105 27863
rect 14105 27829 14139 27863
rect 14139 27829 14148 27863
rect 14096 27820 14148 27829
rect 15108 27956 15160 28008
rect 16764 27956 16816 28008
rect 17132 27999 17184 28008
rect 17132 27965 17141 27999
rect 17141 27965 17175 27999
rect 17175 27965 17184 27999
rect 17132 27956 17184 27965
rect 17408 28033 17417 28067
rect 17417 28033 17451 28067
rect 17451 28033 17460 28067
rect 17408 28024 17460 28033
rect 18604 27956 18656 28008
rect 18880 27956 18932 28008
rect 19064 27956 19116 28008
rect 20260 28024 20312 28076
rect 24216 28024 24268 28076
rect 64328 28024 64380 28076
rect 84200 28024 84252 28076
rect 92572 28092 92624 28144
rect 92480 28024 92532 28076
rect 19340 27888 19392 27940
rect 22376 27956 22428 28008
rect 23296 27956 23348 28008
rect 26240 27956 26292 28008
rect 32128 27956 32180 28008
rect 33140 27999 33192 28008
rect 33140 27965 33149 27999
rect 33149 27965 33183 27999
rect 33183 27965 33192 27999
rect 33140 27956 33192 27965
rect 33600 27931 33652 27940
rect 33600 27897 33609 27931
rect 33609 27897 33643 27931
rect 33643 27897 33652 27931
rect 34796 27956 34848 28008
rect 38936 27956 38988 28008
rect 41512 27956 41564 28008
rect 73804 27956 73856 28008
rect 74356 27956 74408 28008
rect 33600 27888 33652 27897
rect 51080 27888 51132 27940
rect 51172 27888 51224 27940
rect 69848 27888 69900 27940
rect 17960 27820 18012 27872
rect 19156 27863 19208 27872
rect 19156 27829 19165 27863
rect 19165 27829 19199 27863
rect 19199 27829 19208 27863
rect 19156 27820 19208 27829
rect 19248 27820 19300 27872
rect 20536 27820 20588 27872
rect 74724 27820 74776 27872
rect 85580 27820 85632 27872
rect 87604 27999 87656 28008
rect 87604 27965 87613 27999
rect 87613 27965 87647 27999
rect 87647 27965 87656 27999
rect 87604 27956 87656 27965
rect 87696 27956 87748 28008
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 50326 27718 50378 27770
rect 50390 27718 50442 27770
rect 50454 27718 50506 27770
rect 50518 27718 50570 27770
rect 81046 27718 81098 27770
rect 81110 27718 81162 27770
rect 81174 27718 81226 27770
rect 81238 27718 81290 27770
rect 3976 27616 4028 27668
rect 20536 27616 20588 27668
rect 21364 27616 21416 27668
rect 21548 27616 21600 27668
rect 23204 27616 23256 27668
rect 28908 27616 28960 27668
rect 29092 27659 29144 27668
rect 29092 27625 29101 27659
rect 29101 27625 29135 27659
rect 29135 27625 29144 27659
rect 29092 27616 29144 27625
rect 33508 27616 33560 27668
rect 38016 27616 38068 27668
rect 11796 27591 11848 27600
rect 11796 27557 11805 27591
rect 11805 27557 11839 27591
rect 11839 27557 11848 27591
rect 11796 27548 11848 27557
rect 11244 27523 11296 27532
rect 11244 27489 11253 27523
rect 11253 27489 11287 27523
rect 11287 27489 11296 27523
rect 11244 27480 11296 27489
rect 11520 27523 11572 27532
rect 11520 27489 11529 27523
rect 11529 27489 11563 27523
rect 11563 27489 11572 27523
rect 11520 27480 11572 27489
rect 11704 27523 11756 27532
rect 11704 27489 11713 27523
rect 11713 27489 11747 27523
rect 11747 27489 11756 27523
rect 11704 27480 11756 27489
rect 11152 27412 11204 27464
rect 15200 27548 15252 27600
rect 12808 27523 12860 27532
rect 12808 27489 12817 27523
rect 12817 27489 12851 27523
rect 12851 27489 12860 27523
rect 12808 27480 12860 27489
rect 26148 27548 26200 27600
rect 23664 27523 23716 27532
rect 23664 27489 23673 27523
rect 23673 27489 23707 27523
rect 23707 27489 23716 27523
rect 23664 27480 23716 27489
rect 27804 27523 27856 27532
rect 27804 27489 27813 27523
rect 27813 27489 27847 27523
rect 27847 27489 27856 27523
rect 27804 27480 27856 27489
rect 27896 27480 27948 27532
rect 33324 27548 33376 27600
rect 34336 27548 34388 27600
rect 35900 27548 35952 27600
rect 35992 27548 36044 27600
rect 38568 27548 38620 27600
rect 28908 27480 28960 27532
rect 30380 27480 30432 27532
rect 30472 27480 30524 27532
rect 38752 27548 38804 27600
rect 40040 27616 40092 27668
rect 41236 27616 41288 27668
rect 41420 27616 41472 27668
rect 46204 27616 46256 27668
rect 51080 27616 51132 27668
rect 51172 27616 51224 27668
rect 53932 27616 53984 27668
rect 59360 27616 59412 27668
rect 61844 27616 61896 27668
rect 69756 27616 69808 27668
rect 74264 27616 74316 27668
rect 39028 27480 39080 27532
rect 13912 27412 13964 27464
rect 14372 27412 14424 27464
rect 15844 27455 15896 27464
rect 15844 27421 15853 27455
rect 15853 27421 15887 27455
rect 15887 27421 15896 27455
rect 15844 27412 15896 27421
rect 16028 27412 16080 27464
rect 22008 27412 22060 27464
rect 27528 27455 27580 27464
rect 27528 27421 27537 27455
rect 27537 27421 27571 27455
rect 27571 27421 27580 27455
rect 27528 27412 27580 27421
rect 15476 27344 15528 27396
rect 12716 27276 12768 27328
rect 12992 27319 13044 27328
rect 12992 27285 13001 27319
rect 13001 27285 13035 27319
rect 13035 27285 13044 27319
rect 12992 27276 13044 27285
rect 17592 27276 17644 27328
rect 21916 27276 21968 27328
rect 23020 27344 23072 27396
rect 27160 27344 27212 27396
rect 32680 27412 32732 27464
rect 35256 27412 35308 27464
rect 38016 27412 38068 27464
rect 38844 27412 38896 27464
rect 39580 27480 39632 27532
rect 39304 27455 39356 27464
rect 39304 27421 39313 27455
rect 39313 27421 39347 27455
rect 39347 27421 39356 27455
rect 39304 27412 39356 27421
rect 39672 27455 39724 27464
rect 39672 27421 39681 27455
rect 39681 27421 39715 27455
rect 39715 27421 39724 27455
rect 39672 27412 39724 27421
rect 28632 27344 28684 27396
rect 40500 27344 40552 27396
rect 41512 27523 41564 27532
rect 41512 27489 41521 27523
rect 41521 27489 41555 27523
rect 41555 27489 41564 27523
rect 41512 27480 41564 27489
rect 50620 27548 50672 27600
rect 50712 27548 50764 27600
rect 52828 27548 52880 27600
rect 42064 27523 42116 27532
rect 41696 27455 41748 27464
rect 41696 27421 41705 27455
rect 41705 27421 41739 27455
rect 41739 27421 41748 27455
rect 41696 27412 41748 27421
rect 42064 27489 42073 27523
rect 42073 27489 42107 27523
rect 42107 27489 42116 27523
rect 42064 27480 42116 27489
rect 29000 27276 29052 27328
rect 31024 27276 31076 27328
rect 33876 27276 33928 27328
rect 37648 27276 37700 27328
rect 38016 27276 38068 27328
rect 40960 27276 41012 27328
rect 41328 27319 41380 27328
rect 41328 27285 41337 27319
rect 41337 27285 41371 27319
rect 41371 27285 41380 27319
rect 41328 27276 41380 27285
rect 41788 27344 41840 27396
rect 53288 27480 53340 27532
rect 53380 27523 53432 27532
rect 53380 27489 53388 27523
rect 53388 27489 53422 27523
rect 53422 27489 53432 27523
rect 53380 27480 53432 27489
rect 53748 27523 53800 27532
rect 53748 27489 53757 27523
rect 53757 27489 53791 27523
rect 53791 27489 53800 27523
rect 53748 27480 53800 27489
rect 53932 27480 53984 27532
rect 72056 27548 72108 27600
rect 76748 27548 76800 27600
rect 46204 27412 46256 27464
rect 42524 27344 42576 27396
rect 50712 27344 50764 27396
rect 42800 27276 42852 27328
rect 53104 27344 53156 27396
rect 52368 27276 52420 27328
rect 53840 27412 53892 27464
rect 60464 27412 60516 27464
rect 91652 27480 91704 27532
rect 72148 27412 72200 27464
rect 78312 27412 78364 27464
rect 79324 27455 79376 27464
rect 79324 27421 79333 27455
rect 79333 27421 79367 27455
rect 79367 27421 79376 27455
rect 79324 27412 79376 27421
rect 79600 27455 79652 27464
rect 79600 27421 79609 27455
rect 79609 27421 79643 27455
rect 79643 27421 79652 27455
rect 79600 27412 79652 27421
rect 83556 27412 83608 27464
rect 86868 27412 86920 27464
rect 53656 27344 53708 27396
rect 72608 27344 72660 27396
rect 83280 27344 83332 27396
rect 87052 27344 87104 27396
rect 53932 27276 53984 27328
rect 55680 27276 55732 27328
rect 60648 27276 60700 27328
rect 60924 27276 60976 27328
rect 68100 27276 68152 27328
rect 74356 27276 74408 27328
rect 84844 27276 84896 27328
rect 94412 27276 94464 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 65686 27174 65738 27226
rect 65750 27174 65802 27226
rect 65814 27174 65866 27226
rect 65878 27174 65930 27226
rect 96406 27174 96458 27226
rect 96470 27174 96522 27226
rect 96534 27174 96586 27226
rect 96598 27174 96650 27226
rect 12716 27072 12768 27124
rect 14188 27072 14240 27124
rect 15936 27072 15988 27124
rect 17592 27072 17644 27124
rect 18144 27072 18196 27124
rect 19892 27072 19944 27124
rect 21640 27072 21692 27124
rect 21824 27072 21876 27124
rect 28632 27072 28684 27124
rect 28908 27072 28960 27124
rect 35256 27072 35308 27124
rect 37648 27072 37700 27124
rect 46204 27072 46256 27124
rect 46296 27072 46348 27124
rect 55680 27072 55732 27124
rect 7288 27004 7340 27056
rect 21548 27004 21600 27056
rect 22284 27004 22336 27056
rect 41420 27004 41472 27056
rect 43352 27004 43404 27056
rect 56048 27004 56100 27056
rect 60648 27072 60700 27124
rect 84844 27072 84896 27124
rect 14096 26936 14148 26988
rect 21824 26936 21876 26988
rect 22008 26936 22060 26988
rect 29000 26936 29052 26988
rect 29920 26936 29972 26988
rect 30288 26936 30340 26988
rect 36176 26936 36228 26988
rect 36636 26936 36688 26988
rect 38936 26936 38988 26988
rect 39672 26936 39724 26988
rect 40408 26936 40460 26988
rect 40868 26936 40920 26988
rect 40960 26936 41012 26988
rect 59176 26936 59228 26988
rect 75092 27004 75144 27056
rect 77668 27004 77720 27056
rect 78220 27004 78272 27056
rect 79324 27004 79376 27056
rect 80888 27004 80940 27056
rect 61200 26979 61252 26988
rect 17316 26868 17368 26920
rect 17868 26868 17920 26920
rect 21088 26868 21140 26920
rect 35992 26868 36044 26920
rect 5356 26800 5408 26852
rect 23204 26800 23256 26852
rect 27528 26800 27580 26852
rect 30840 26800 30892 26852
rect 30932 26800 30984 26852
rect 37188 26868 37240 26920
rect 37280 26868 37332 26920
rect 37924 26868 37976 26920
rect 38660 26868 38712 26920
rect 39396 26868 39448 26920
rect 41604 26868 41656 26920
rect 41880 26868 41932 26920
rect 48228 26868 48280 26920
rect 48412 26868 48464 26920
rect 49240 26868 49292 26920
rect 49884 26868 49936 26920
rect 50712 26868 50764 26920
rect 36360 26800 36412 26852
rect 52552 26868 52604 26920
rect 52644 26868 52696 26920
rect 53472 26868 53524 26920
rect 54208 26868 54260 26920
rect 54944 26868 54996 26920
rect 55036 26868 55088 26920
rect 59912 26911 59964 26920
rect 59912 26877 59921 26911
rect 59921 26877 59955 26911
rect 59955 26877 59964 26911
rect 61200 26945 61209 26979
rect 61209 26945 61243 26979
rect 61243 26945 61252 26979
rect 61200 26936 61252 26945
rect 87512 27004 87564 27056
rect 94320 27004 94372 27056
rect 94780 27047 94832 27056
rect 94780 27013 94789 27047
rect 94789 27013 94823 27047
rect 94823 27013 94832 27047
rect 94780 27004 94832 27013
rect 59912 26868 59964 26877
rect 75552 26868 75604 26920
rect 77392 26868 77444 26920
rect 52828 26800 52880 26852
rect 59268 26800 59320 26852
rect 17960 26732 18012 26784
rect 63040 26800 63092 26852
rect 68836 26800 68888 26852
rect 69020 26800 69072 26852
rect 77024 26800 77076 26852
rect 78220 26911 78272 26920
rect 78220 26877 78229 26911
rect 78229 26877 78263 26911
rect 78263 26877 78272 26911
rect 78220 26868 78272 26877
rect 80888 26868 80940 26920
rect 86224 26936 86276 26988
rect 86500 26936 86552 26988
rect 87420 26936 87472 26988
rect 78496 26800 78548 26852
rect 86684 26868 86736 26920
rect 86868 26868 86920 26920
rect 94504 26911 94556 26920
rect 94504 26877 94513 26911
rect 94513 26877 94547 26911
rect 94547 26877 94556 26911
rect 94504 26868 94556 26877
rect 78128 26775 78180 26784
rect 78128 26741 78137 26775
rect 78137 26741 78171 26775
rect 78171 26741 78180 26775
rect 78128 26732 78180 26741
rect 79416 26732 79468 26784
rect 87512 26732 87564 26784
rect 87788 26732 87840 26784
rect 95148 26868 95200 26920
rect 96896 26911 96948 26920
rect 96896 26877 96905 26911
rect 96905 26877 96939 26911
rect 96939 26877 96948 26911
rect 96896 26868 96948 26877
rect 97448 26911 97500 26920
rect 97448 26877 97457 26911
rect 97457 26877 97491 26911
rect 97491 26877 97500 26911
rect 97448 26868 97500 26877
rect 97816 26732 97868 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 50326 26630 50378 26682
rect 50390 26630 50442 26682
rect 50454 26630 50506 26682
rect 50518 26630 50570 26682
rect 81046 26630 81098 26682
rect 81110 26630 81162 26682
rect 81174 26630 81226 26682
rect 81238 26630 81290 26682
rect 5356 26571 5408 26580
rect 5356 26537 5365 26571
rect 5365 26537 5399 26571
rect 5399 26537 5408 26571
rect 5356 26528 5408 26537
rect 13544 26528 13596 26580
rect 21548 26528 21600 26580
rect 30380 26528 30432 26580
rect 30564 26571 30616 26580
rect 30564 26537 30573 26571
rect 30573 26537 30607 26571
rect 30607 26537 30616 26571
rect 30564 26528 30616 26537
rect 30840 26528 30892 26580
rect 33416 26528 33468 26580
rect 35256 26528 35308 26580
rect 37096 26528 37148 26580
rect 37188 26528 37240 26580
rect 40960 26528 41012 26580
rect 41512 26528 41564 26580
rect 87512 26528 87564 26580
rect 90456 26571 90508 26580
rect 90456 26537 90465 26571
rect 90465 26537 90499 26571
rect 90499 26537 90508 26571
rect 90456 26528 90508 26537
rect 4712 26435 4764 26444
rect 4712 26401 4721 26435
rect 4721 26401 4755 26435
rect 4755 26401 4764 26435
rect 4712 26392 4764 26401
rect 4620 26299 4672 26308
rect 4620 26265 4629 26299
rect 4629 26265 4663 26299
rect 4663 26265 4672 26299
rect 5172 26392 5224 26444
rect 10324 26460 10376 26512
rect 6736 26392 6788 26444
rect 14004 26392 14056 26444
rect 5080 26367 5132 26376
rect 5080 26333 5089 26367
rect 5089 26333 5123 26367
rect 5123 26333 5132 26367
rect 15108 26367 15160 26376
rect 5080 26324 5132 26333
rect 15108 26333 15117 26367
rect 15117 26333 15151 26367
rect 15151 26333 15160 26367
rect 15108 26324 15160 26333
rect 19064 26392 19116 26444
rect 20720 26460 20772 26512
rect 21640 26460 21692 26512
rect 33692 26460 33744 26512
rect 36728 26460 36780 26512
rect 40500 26460 40552 26512
rect 46664 26460 46716 26512
rect 21088 26392 21140 26444
rect 21272 26392 21324 26444
rect 21916 26392 21968 26444
rect 26332 26392 26384 26444
rect 26884 26392 26936 26444
rect 27160 26392 27212 26444
rect 30472 26435 30524 26444
rect 30472 26401 30481 26435
rect 30481 26401 30515 26435
rect 30515 26401 30524 26435
rect 30472 26392 30524 26401
rect 30656 26392 30708 26444
rect 30932 26435 30984 26444
rect 30932 26401 30941 26435
rect 30941 26401 30975 26435
rect 30975 26401 30984 26435
rect 30932 26392 30984 26401
rect 31024 26392 31076 26444
rect 33324 26392 33376 26444
rect 34336 26392 34388 26444
rect 35808 26392 35860 26444
rect 35992 26435 36044 26444
rect 35992 26401 36001 26435
rect 36001 26401 36035 26435
rect 36035 26401 36044 26435
rect 35992 26392 36044 26401
rect 36360 26392 36412 26444
rect 36452 26392 36504 26444
rect 41052 26392 41104 26444
rect 47584 26392 47636 26444
rect 48228 26435 48280 26444
rect 48228 26401 48237 26435
rect 48237 26401 48271 26435
rect 48271 26401 48280 26435
rect 48228 26392 48280 26401
rect 48596 26435 48648 26444
rect 48596 26401 48605 26435
rect 48605 26401 48639 26435
rect 48639 26401 48648 26435
rect 48596 26392 48648 26401
rect 4620 26256 4672 26265
rect 13452 26256 13504 26308
rect 11520 26188 11572 26240
rect 17592 26256 17644 26308
rect 21272 26256 21324 26308
rect 33692 26324 33744 26376
rect 36084 26367 36136 26376
rect 36084 26333 36093 26367
rect 36093 26333 36127 26367
rect 36127 26333 36136 26367
rect 36084 26324 36136 26333
rect 36728 26324 36780 26376
rect 42892 26324 42944 26376
rect 45376 26324 45428 26376
rect 45836 26324 45888 26376
rect 48044 26367 48096 26376
rect 48044 26333 48053 26367
rect 48053 26333 48087 26367
rect 48087 26333 48096 26367
rect 48044 26324 48096 26333
rect 48320 26324 48372 26376
rect 50068 26460 50120 26512
rect 60556 26460 60608 26512
rect 60648 26460 60700 26512
rect 87788 26460 87840 26512
rect 49884 26392 49936 26444
rect 50252 26435 50304 26444
rect 50252 26401 50261 26435
rect 50261 26401 50295 26435
rect 50295 26401 50304 26435
rect 50252 26392 50304 26401
rect 50344 26435 50396 26444
rect 50344 26401 50353 26435
rect 50353 26401 50387 26435
rect 50387 26401 50396 26435
rect 50344 26392 50396 26401
rect 52552 26392 52604 26444
rect 53840 26392 53892 26444
rect 57888 26392 57940 26444
rect 59268 26392 59320 26444
rect 59452 26392 59504 26444
rect 60280 26392 60332 26444
rect 60372 26392 60424 26444
rect 64604 26392 64656 26444
rect 64696 26392 64748 26444
rect 70584 26392 70636 26444
rect 72884 26392 72936 26444
rect 72516 26324 72568 26376
rect 48688 26256 48740 26308
rect 48872 26256 48924 26308
rect 53104 26256 53156 26308
rect 60372 26256 60424 26308
rect 60464 26256 60516 26308
rect 64696 26256 64748 26308
rect 73344 26256 73396 26308
rect 73804 26392 73856 26444
rect 74080 26435 74132 26444
rect 73620 26367 73672 26376
rect 73620 26333 73629 26367
rect 73629 26333 73663 26367
rect 73663 26333 73672 26367
rect 73620 26324 73672 26333
rect 74080 26401 74089 26435
rect 74089 26401 74123 26435
rect 74123 26401 74132 26435
rect 74080 26392 74132 26401
rect 75092 26392 75144 26444
rect 86316 26392 86368 26444
rect 86408 26435 86460 26444
rect 86408 26401 86417 26435
rect 86417 26401 86451 26435
rect 86451 26401 86460 26435
rect 86408 26392 86460 26401
rect 86684 26435 86736 26444
rect 73988 26324 74040 26376
rect 74356 26324 74408 26376
rect 86132 26324 86184 26376
rect 74632 26256 74684 26308
rect 83556 26256 83608 26308
rect 83648 26256 83700 26308
rect 43260 26188 43312 26240
rect 43352 26188 43404 26240
rect 49884 26188 49936 26240
rect 50068 26188 50120 26240
rect 52828 26188 52880 26240
rect 60188 26188 60240 26240
rect 61292 26188 61344 26240
rect 63500 26188 63552 26240
rect 65432 26188 65484 26240
rect 73436 26188 73488 26240
rect 74264 26188 74316 26240
rect 81808 26188 81860 26240
rect 86316 26256 86368 26308
rect 86684 26401 86693 26435
rect 86693 26401 86727 26435
rect 86727 26401 86736 26435
rect 86684 26392 86736 26401
rect 86868 26392 86920 26444
rect 87052 26392 87104 26444
rect 91652 26435 91704 26444
rect 91652 26401 91661 26435
rect 91661 26401 91695 26435
rect 91695 26401 91704 26435
rect 91652 26392 91704 26401
rect 91836 26435 91888 26444
rect 91836 26401 91845 26435
rect 91845 26401 91879 26435
rect 91879 26401 91888 26435
rect 91836 26392 91888 26401
rect 87972 26367 88024 26376
rect 87972 26333 87981 26367
rect 87981 26333 88015 26367
rect 88015 26333 88024 26367
rect 87972 26324 88024 26333
rect 88248 26324 88300 26376
rect 91560 26324 91612 26376
rect 91928 26256 91980 26308
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 65686 26086 65738 26138
rect 65750 26086 65802 26138
rect 65814 26086 65866 26138
rect 65878 26086 65930 26138
rect 96406 26086 96458 26138
rect 96470 26086 96522 26138
rect 96534 26086 96586 26138
rect 96598 26086 96650 26138
rect 11704 25984 11756 26036
rect 15108 25916 15160 25968
rect 15936 25916 15988 25968
rect 20352 25984 20404 26036
rect 26884 25984 26936 26036
rect 41420 25984 41472 26036
rect 41512 25984 41564 26036
rect 31852 25916 31904 25968
rect 37004 25916 37056 25968
rect 37464 25916 37516 25968
rect 38200 25916 38252 25968
rect 38292 25916 38344 25968
rect 45560 25916 45612 25968
rect 45652 25916 45704 25968
rect 50436 25916 50488 25968
rect 53748 25984 53800 26036
rect 65432 25984 65484 26036
rect 77484 25984 77536 26036
rect 69112 25916 69164 25968
rect 73436 25916 73488 25968
rect 75920 25916 75972 25968
rect 91560 25916 91612 25968
rect 17224 25848 17276 25900
rect 18880 25780 18932 25832
rect 19064 25823 19116 25832
rect 19064 25789 19073 25823
rect 19073 25789 19107 25823
rect 19107 25789 19116 25823
rect 19064 25780 19116 25789
rect 20352 25780 20404 25832
rect 19892 25712 19944 25764
rect 22928 25823 22980 25832
rect 22928 25789 22937 25823
rect 22937 25789 22971 25823
rect 22971 25789 22980 25823
rect 22928 25780 22980 25789
rect 24492 25848 24544 25900
rect 15476 25644 15528 25696
rect 20904 25712 20956 25764
rect 39212 25823 39264 25832
rect 39212 25789 39228 25823
rect 39228 25789 39262 25823
rect 39262 25789 39264 25823
rect 39396 25823 39448 25832
rect 39212 25780 39264 25789
rect 39396 25789 39405 25823
rect 39405 25789 39439 25823
rect 39439 25789 39448 25823
rect 39396 25780 39448 25789
rect 39580 25823 39632 25832
rect 39580 25789 39589 25823
rect 39589 25789 39623 25823
rect 39623 25789 39632 25823
rect 39856 25823 39908 25832
rect 39580 25780 39632 25789
rect 39856 25789 39865 25823
rect 39865 25789 39899 25823
rect 39899 25789 39908 25823
rect 39856 25780 39908 25789
rect 20260 25644 20312 25696
rect 26884 25644 26936 25696
rect 34612 25644 34664 25696
rect 35808 25644 35860 25696
rect 35992 25644 36044 25696
rect 38016 25644 38068 25696
rect 39580 25644 39632 25696
rect 43352 25712 43404 25764
rect 43536 25780 43588 25832
rect 52828 25780 52880 25832
rect 49792 25712 49844 25764
rect 50436 25712 50488 25764
rect 52368 25712 52420 25764
rect 56232 25848 56284 25900
rect 65432 25848 65484 25900
rect 56048 25780 56100 25832
rect 61200 25780 61252 25832
rect 61660 25823 61712 25832
rect 61660 25789 61669 25823
rect 61669 25789 61703 25823
rect 61703 25789 61712 25823
rect 61660 25780 61712 25789
rect 61752 25780 61804 25832
rect 65248 25780 65300 25832
rect 86592 25848 86644 25900
rect 87420 25848 87472 25900
rect 66352 25823 66404 25832
rect 66352 25789 66361 25823
rect 66361 25789 66395 25823
rect 66395 25789 66404 25823
rect 66352 25780 66404 25789
rect 67180 25823 67232 25832
rect 67180 25789 67189 25823
rect 67189 25789 67223 25823
rect 67223 25789 67232 25823
rect 67180 25780 67232 25789
rect 67548 25780 67600 25832
rect 73252 25780 73304 25832
rect 73988 25780 74040 25832
rect 80428 25823 80480 25832
rect 80428 25789 80437 25823
rect 80437 25789 80471 25823
rect 80471 25789 80480 25823
rect 80428 25780 80480 25789
rect 70124 25712 70176 25764
rect 82176 25712 82228 25764
rect 82728 25712 82780 25764
rect 93216 25644 93268 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 50326 25542 50378 25594
rect 50390 25542 50442 25594
rect 50454 25542 50506 25594
rect 50518 25542 50570 25594
rect 81046 25542 81098 25594
rect 81110 25542 81162 25594
rect 81174 25542 81226 25594
rect 81238 25542 81290 25594
rect 15200 25440 15252 25492
rect 20904 25440 20956 25492
rect 21824 25440 21876 25492
rect 21916 25440 21968 25492
rect 37372 25440 37424 25492
rect 38568 25440 38620 25492
rect 39396 25440 39448 25492
rect 3056 25372 3108 25424
rect 21180 25372 21232 25424
rect 21732 25304 21784 25356
rect 22100 25304 22152 25356
rect 22468 25304 22520 25356
rect 19892 25236 19944 25288
rect 30932 25304 30984 25356
rect 32128 25372 32180 25424
rect 42340 25372 42392 25424
rect 42616 25415 42668 25424
rect 42616 25381 42625 25415
rect 42625 25381 42659 25415
rect 42659 25381 42668 25415
rect 42616 25372 42668 25381
rect 52092 25440 52144 25492
rect 53196 25440 53248 25492
rect 54576 25440 54628 25492
rect 56324 25440 56376 25492
rect 56508 25440 56560 25492
rect 60740 25440 60792 25492
rect 61384 25440 61436 25492
rect 65248 25440 65300 25492
rect 70124 25440 70176 25492
rect 70216 25440 70268 25492
rect 82360 25440 82412 25492
rect 38660 25304 38712 25356
rect 40500 25304 40552 25356
rect 25872 25236 25924 25288
rect 39028 25236 39080 25288
rect 41328 25304 41380 25356
rect 41512 25304 41564 25356
rect 41880 25304 41932 25356
rect 43720 25372 43772 25424
rect 43628 25347 43680 25356
rect 43628 25313 43637 25347
rect 43637 25313 43671 25347
rect 43671 25313 43680 25347
rect 43628 25304 43680 25313
rect 17776 25168 17828 25220
rect 15200 25100 15252 25152
rect 15384 25100 15436 25152
rect 21824 25100 21876 25152
rect 21916 25100 21968 25152
rect 27712 25143 27764 25152
rect 27712 25109 27721 25143
rect 27721 25109 27755 25143
rect 27755 25109 27764 25143
rect 27712 25100 27764 25109
rect 30472 25168 30524 25220
rect 39856 25168 39908 25220
rect 40684 25168 40736 25220
rect 43352 25236 43404 25288
rect 44088 25304 44140 25356
rect 44548 25304 44600 25356
rect 47584 25372 47636 25424
rect 44272 25236 44324 25288
rect 45652 25236 45704 25288
rect 48504 25304 48556 25356
rect 50988 25304 51040 25356
rect 63132 25372 63184 25424
rect 65432 25372 65484 25424
rect 76472 25372 76524 25424
rect 82728 25372 82780 25424
rect 51816 25347 51868 25356
rect 51816 25313 51825 25347
rect 51825 25313 51859 25347
rect 51859 25313 51868 25347
rect 51816 25304 51868 25313
rect 52184 25347 52236 25356
rect 52184 25313 52193 25347
rect 52193 25313 52227 25347
rect 52227 25313 52236 25347
rect 52184 25304 52236 25313
rect 53196 25347 53248 25356
rect 48412 25236 48464 25288
rect 48596 25236 48648 25288
rect 49516 25236 49568 25288
rect 51908 25279 51960 25288
rect 51264 25168 51316 25220
rect 51908 25245 51917 25279
rect 51917 25245 51951 25279
rect 51951 25245 51960 25279
rect 51908 25236 51960 25245
rect 53196 25313 53205 25347
rect 53205 25313 53239 25347
rect 53239 25313 53248 25347
rect 53196 25304 53248 25313
rect 53564 25304 53616 25356
rect 53656 25304 53708 25356
rect 56048 25236 56100 25288
rect 56232 25304 56284 25356
rect 61292 25304 61344 25356
rect 61384 25304 61436 25356
rect 64972 25304 65024 25356
rect 66444 25304 66496 25356
rect 81808 25304 81860 25356
rect 89536 25304 89588 25356
rect 74356 25279 74408 25288
rect 74356 25245 74365 25279
rect 74365 25245 74399 25279
rect 74399 25245 74408 25279
rect 74356 25236 74408 25245
rect 90456 25236 90508 25288
rect 91284 25279 91336 25288
rect 91284 25245 91293 25279
rect 91293 25245 91327 25279
rect 91327 25245 91336 25279
rect 91284 25236 91336 25245
rect 43628 25100 43680 25152
rect 43720 25100 43772 25152
rect 47492 25100 47544 25152
rect 50436 25100 50488 25152
rect 53748 25168 53800 25220
rect 56784 25168 56836 25220
rect 57520 25168 57572 25220
rect 60004 25168 60056 25220
rect 60188 25168 60240 25220
rect 65616 25168 65668 25220
rect 70216 25168 70268 25220
rect 73160 25168 73212 25220
rect 97448 25168 97500 25220
rect 52828 25143 52880 25152
rect 52828 25109 52837 25143
rect 52837 25109 52871 25143
rect 52871 25109 52880 25143
rect 52828 25100 52880 25109
rect 53196 25100 53248 25152
rect 54760 25100 54812 25152
rect 56508 25100 56560 25152
rect 56876 25100 56928 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 65686 24998 65738 25050
rect 65750 24998 65802 25050
rect 65814 24998 65866 25050
rect 65878 24998 65930 25050
rect 96406 24998 96458 25050
rect 96470 24998 96522 25050
rect 96534 24998 96586 25050
rect 96598 24998 96650 25050
rect 9128 24896 9180 24948
rect 14004 24896 14056 24948
rect 4712 24828 4764 24880
rect 25872 24896 25924 24948
rect 27712 24896 27764 24948
rect 38292 24896 38344 24948
rect 38568 24896 38620 24948
rect 39488 24896 39540 24948
rect 1492 24735 1544 24744
rect 1492 24701 1501 24735
rect 1501 24701 1535 24735
rect 1535 24701 1544 24735
rect 1492 24692 1544 24701
rect 1768 24735 1820 24744
rect 1768 24701 1777 24735
rect 1777 24701 1811 24735
rect 1811 24701 1820 24735
rect 1768 24692 1820 24701
rect 2136 24692 2188 24744
rect 3240 24760 3292 24812
rect 2872 24692 2924 24744
rect 3056 24692 3108 24744
rect 3332 24735 3384 24744
rect 3332 24701 3341 24735
rect 3341 24701 3375 24735
rect 3375 24701 3384 24735
rect 3332 24692 3384 24701
rect 2688 24556 2740 24608
rect 2964 24599 3016 24608
rect 2964 24565 2973 24599
rect 2973 24565 3007 24599
rect 3007 24565 3016 24599
rect 2964 24556 3016 24565
rect 3700 24735 3752 24744
rect 3700 24701 3709 24735
rect 3709 24701 3743 24735
rect 3743 24701 3752 24735
rect 3700 24692 3752 24701
rect 12716 24760 12768 24812
rect 12808 24760 12860 24812
rect 16488 24760 16540 24812
rect 17132 24760 17184 24812
rect 18420 24760 18472 24812
rect 24492 24760 24544 24812
rect 13452 24692 13504 24744
rect 36912 24828 36964 24880
rect 37096 24828 37148 24880
rect 43536 24828 43588 24880
rect 44640 24828 44692 24880
rect 50436 24828 50488 24880
rect 52828 24896 52880 24948
rect 66260 24896 66312 24948
rect 69296 24896 69348 24948
rect 91284 24896 91336 24948
rect 56232 24828 56284 24880
rect 56324 24828 56376 24880
rect 69940 24828 69992 24880
rect 71412 24871 71464 24880
rect 71412 24837 71421 24871
rect 71421 24837 71455 24871
rect 71455 24837 71464 24871
rect 71412 24828 71464 24837
rect 72700 24828 72752 24880
rect 75828 24828 75880 24880
rect 35992 24760 36044 24812
rect 50528 24760 50580 24812
rect 51356 24760 51408 24812
rect 87972 24760 88024 24812
rect 5080 24624 5132 24676
rect 5356 24624 5408 24676
rect 36912 24692 36964 24744
rect 39304 24692 39356 24744
rect 40500 24692 40552 24744
rect 40684 24692 40736 24744
rect 41420 24692 41472 24744
rect 43812 24735 43864 24744
rect 43812 24701 43821 24735
rect 43821 24701 43855 24735
rect 43855 24701 43864 24735
rect 43812 24692 43864 24701
rect 44732 24692 44784 24744
rect 44916 24692 44968 24744
rect 45468 24692 45520 24744
rect 47308 24692 47360 24744
rect 48780 24692 48832 24744
rect 50988 24692 51040 24744
rect 51172 24735 51224 24744
rect 51172 24701 51181 24735
rect 51181 24701 51215 24735
rect 51215 24701 51224 24735
rect 51172 24692 51224 24701
rect 51540 24692 51592 24744
rect 22744 24624 22796 24676
rect 28080 24624 28132 24676
rect 34244 24624 34296 24676
rect 37004 24624 37056 24676
rect 43628 24624 43680 24676
rect 14740 24556 14792 24608
rect 18052 24556 18104 24608
rect 22560 24556 22612 24608
rect 23112 24556 23164 24608
rect 30380 24556 30432 24608
rect 30840 24556 30892 24608
rect 46112 24624 46164 24676
rect 50528 24624 50580 24676
rect 52460 24599 52512 24608
rect 52460 24565 52469 24599
rect 52469 24565 52503 24599
rect 52503 24565 52512 24599
rect 52460 24556 52512 24565
rect 55680 24624 55732 24676
rect 63408 24624 63460 24676
rect 65524 24692 65576 24744
rect 72792 24692 72844 24744
rect 66904 24624 66956 24676
rect 67272 24624 67324 24676
rect 74632 24624 74684 24676
rect 75644 24624 75696 24676
rect 78312 24735 78364 24744
rect 78312 24701 78321 24735
rect 78321 24701 78355 24735
rect 78355 24701 78364 24735
rect 78312 24692 78364 24701
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 50326 24454 50378 24506
rect 50390 24454 50442 24506
rect 50454 24454 50506 24506
rect 50518 24454 50570 24506
rect 81046 24454 81098 24506
rect 81110 24454 81162 24506
rect 81174 24454 81226 24506
rect 81238 24454 81290 24506
rect 3700 24352 3752 24404
rect 12624 24352 12676 24404
rect 13360 24352 13412 24404
rect 15108 24284 15160 24336
rect 21824 24395 21876 24404
rect 4712 24216 4764 24268
rect 10600 24148 10652 24200
rect 10876 24148 10928 24200
rect 16948 24216 17000 24268
rect 17132 24259 17184 24268
rect 17132 24225 17141 24259
rect 17141 24225 17175 24259
rect 17175 24225 17184 24259
rect 17132 24216 17184 24225
rect 19064 24284 19116 24336
rect 21824 24361 21833 24395
rect 21833 24361 21867 24395
rect 21867 24361 21876 24395
rect 21824 24352 21876 24361
rect 25136 24352 25188 24404
rect 43536 24352 43588 24404
rect 43996 24352 44048 24404
rect 25320 24284 25372 24336
rect 42800 24284 42852 24336
rect 43628 24284 43680 24336
rect 46112 24284 46164 24336
rect 46388 24327 46440 24336
rect 46388 24293 46397 24327
rect 46397 24293 46431 24327
rect 46431 24293 46440 24327
rect 46388 24284 46440 24293
rect 46480 24327 46532 24336
rect 46480 24293 46489 24327
rect 46489 24293 46523 24327
rect 46523 24293 46532 24327
rect 46480 24284 46532 24293
rect 46664 24284 46716 24336
rect 22560 24259 22612 24268
rect 19616 24148 19668 24200
rect 20720 24191 20772 24200
rect 20720 24157 20729 24191
rect 20729 24157 20763 24191
rect 20763 24157 20772 24191
rect 20720 24148 20772 24157
rect 22560 24225 22569 24259
rect 22569 24225 22603 24259
rect 22603 24225 22612 24259
rect 22560 24216 22612 24225
rect 42248 24216 42300 24268
rect 44364 24216 44416 24268
rect 44732 24216 44784 24268
rect 46296 24216 46348 24268
rect 23020 24148 23072 24200
rect 23296 24191 23348 24200
rect 23296 24157 23305 24191
rect 23305 24157 23339 24191
rect 23339 24157 23348 24191
rect 23296 24148 23348 24157
rect 24216 24148 24268 24200
rect 24768 24148 24820 24200
rect 25228 24148 25280 24200
rect 25320 24148 25372 24200
rect 43996 24148 44048 24200
rect 45376 24148 45428 24200
rect 45836 24148 45888 24200
rect 11152 24012 11204 24064
rect 19524 24012 19576 24064
rect 20168 24012 20220 24064
rect 40960 24080 41012 24132
rect 41052 24080 41104 24132
rect 46388 24080 46440 24132
rect 46940 24352 46992 24404
rect 65524 24352 65576 24404
rect 48136 24284 48188 24336
rect 63500 24284 63552 24336
rect 75000 24352 75052 24404
rect 66260 24284 66312 24336
rect 72700 24284 72752 24336
rect 72792 24284 72844 24336
rect 75828 24327 75880 24336
rect 75828 24293 75837 24327
rect 75837 24293 75871 24327
rect 75871 24293 75880 24327
rect 75828 24284 75880 24293
rect 86868 24352 86920 24404
rect 91928 24352 91980 24404
rect 47308 24216 47360 24268
rect 75092 24216 75144 24268
rect 75736 24259 75788 24268
rect 75736 24225 75745 24259
rect 75745 24225 75779 24259
rect 75779 24225 75788 24259
rect 75736 24216 75788 24225
rect 75920 24259 75972 24268
rect 75920 24225 75929 24259
rect 75929 24225 75963 24259
rect 75963 24225 75972 24259
rect 75920 24216 75972 24225
rect 72792 24148 72844 24200
rect 46940 24080 46992 24132
rect 55680 24080 55732 24132
rect 23020 24012 23072 24064
rect 26884 24012 26936 24064
rect 28540 24012 28592 24064
rect 35992 24012 36044 24064
rect 36452 24012 36504 24064
rect 43260 24012 43312 24064
rect 44088 24012 44140 24064
rect 61200 24012 61252 24064
rect 63224 24012 63276 24064
rect 63408 24012 63460 24064
rect 65432 24012 65484 24064
rect 71688 24080 71740 24132
rect 74724 24080 74776 24132
rect 75092 24080 75144 24132
rect 78312 24216 78364 24268
rect 78496 24216 78548 24268
rect 76288 24191 76340 24200
rect 76288 24157 76297 24191
rect 76297 24157 76331 24191
rect 76331 24157 76340 24191
rect 76288 24148 76340 24157
rect 76380 24148 76432 24200
rect 90180 24284 90232 24336
rect 90824 24284 90876 24336
rect 83188 24259 83240 24268
rect 83188 24225 83196 24259
rect 83196 24225 83230 24259
rect 83230 24225 83240 24259
rect 83556 24259 83608 24268
rect 83188 24216 83240 24225
rect 83556 24225 83565 24259
rect 83565 24225 83599 24259
rect 83599 24225 83608 24259
rect 83556 24216 83608 24225
rect 95332 24216 95384 24268
rect 84016 24148 84068 24200
rect 76012 24012 76064 24064
rect 76288 24012 76340 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 65686 23910 65738 23962
rect 65750 23910 65802 23962
rect 65814 23910 65866 23962
rect 65878 23910 65930 23962
rect 96406 23910 96458 23962
rect 96470 23910 96522 23962
rect 96534 23910 96586 23962
rect 96598 23910 96650 23962
rect 1768 23808 1820 23860
rect 9496 23808 9548 23860
rect 19524 23808 19576 23860
rect 19616 23808 19668 23860
rect 20536 23808 20588 23860
rect 35532 23808 35584 23860
rect 35808 23808 35860 23860
rect 2688 23740 2740 23792
rect 20628 23740 20680 23792
rect 25136 23740 25188 23792
rect 25228 23783 25280 23792
rect 25228 23749 25237 23783
rect 25237 23749 25271 23783
rect 25271 23749 25280 23783
rect 25228 23740 25280 23749
rect 13360 23672 13412 23724
rect 23940 23672 23992 23724
rect 24308 23672 24360 23724
rect 25136 23647 25188 23656
rect 25136 23613 25142 23647
rect 25142 23613 25188 23647
rect 25136 23604 25188 23613
rect 25688 23672 25740 23724
rect 34428 23672 34480 23724
rect 36452 23672 36504 23724
rect 43260 23808 43312 23860
rect 45192 23808 45244 23860
rect 37740 23740 37792 23792
rect 45008 23740 45060 23792
rect 42984 23672 43036 23724
rect 43260 23672 43312 23724
rect 43812 23672 43864 23724
rect 50344 23808 50396 23860
rect 45376 23740 45428 23792
rect 48688 23740 48740 23792
rect 50620 23740 50672 23792
rect 53564 23740 53616 23792
rect 63408 23740 63460 23792
rect 63500 23740 63552 23792
rect 69940 23783 69992 23792
rect 69940 23749 69949 23783
rect 69949 23749 69983 23783
rect 69983 23749 69992 23783
rect 69940 23740 69992 23749
rect 46204 23672 46256 23724
rect 46664 23672 46716 23724
rect 48780 23715 48832 23724
rect 48780 23681 48789 23715
rect 48789 23681 48823 23715
rect 48823 23681 48832 23715
rect 48780 23672 48832 23681
rect 71872 23672 71924 23724
rect 47032 23604 47084 23656
rect 48688 23604 48740 23656
rect 22100 23536 22152 23588
rect 24952 23579 25004 23588
rect 24952 23545 24961 23579
rect 24961 23545 24995 23579
rect 24995 23545 25004 23579
rect 24952 23536 25004 23545
rect 18236 23468 18288 23520
rect 25596 23511 25648 23520
rect 25596 23477 25605 23511
rect 25605 23477 25639 23511
rect 25639 23477 25648 23511
rect 25596 23468 25648 23477
rect 26884 23536 26936 23588
rect 34336 23536 34388 23588
rect 65616 23604 65668 23656
rect 65892 23604 65944 23656
rect 69020 23604 69072 23656
rect 50344 23536 50396 23588
rect 61384 23536 61436 23588
rect 61752 23536 61804 23588
rect 65432 23536 65484 23588
rect 73160 23740 73212 23792
rect 76104 23808 76156 23860
rect 80060 23851 80112 23860
rect 80060 23817 80069 23851
rect 80069 23817 80103 23851
rect 80103 23817 80112 23851
rect 80060 23808 80112 23817
rect 76380 23740 76432 23792
rect 84016 23808 84068 23860
rect 83832 23740 83884 23792
rect 83556 23672 83608 23724
rect 73068 23604 73120 23656
rect 75092 23604 75144 23656
rect 74448 23536 74500 23588
rect 65892 23511 65944 23520
rect 65892 23477 65901 23511
rect 65901 23477 65935 23511
rect 65935 23477 65944 23511
rect 65892 23468 65944 23477
rect 75000 23468 75052 23520
rect 75460 23468 75512 23520
rect 76012 23468 76064 23520
rect 77116 23647 77168 23656
rect 77116 23613 77125 23647
rect 77125 23613 77159 23647
rect 77159 23613 77168 23647
rect 77116 23604 77168 23613
rect 77208 23604 77260 23656
rect 76564 23536 76616 23588
rect 78772 23604 78824 23656
rect 84936 23604 84988 23656
rect 90180 23536 90232 23588
rect 94688 23604 94740 23656
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 50326 23366 50378 23418
rect 50390 23366 50442 23418
rect 50454 23366 50506 23418
rect 50518 23366 50570 23418
rect 81046 23366 81098 23418
rect 81110 23366 81162 23418
rect 81174 23366 81226 23418
rect 81238 23366 81290 23418
rect 1860 23264 1912 23316
rect 6920 23264 6972 23316
rect 2320 23196 2372 23248
rect 17224 23264 17276 23316
rect 25872 23264 25924 23316
rect 26148 23264 26200 23316
rect 29092 23264 29144 23316
rect 29920 23264 29972 23316
rect 35992 23264 36044 23316
rect 36544 23264 36596 23316
rect 37924 23264 37976 23316
rect 48136 23264 48188 23316
rect 48504 23307 48556 23316
rect 48504 23273 48513 23307
rect 48513 23273 48547 23307
rect 48547 23273 48556 23307
rect 48504 23264 48556 23273
rect 48872 23264 48924 23316
rect 49516 23264 49568 23316
rect 56048 23264 56100 23316
rect 56232 23264 56284 23316
rect 11428 23196 11480 23248
rect 14188 23196 14240 23248
rect 39212 23196 39264 23248
rect 6920 23128 6972 23180
rect 7564 23128 7616 23180
rect 9220 23128 9272 23180
rect 14740 23171 14792 23180
rect 9404 23060 9456 23112
rect 9772 23103 9824 23112
rect 9772 23069 9781 23103
rect 9781 23069 9815 23103
rect 9815 23069 9824 23103
rect 9772 23060 9824 23069
rect 14740 23137 14749 23171
rect 14749 23137 14783 23171
rect 14783 23137 14792 23171
rect 14740 23128 14792 23137
rect 14924 23171 14976 23180
rect 14924 23137 14933 23171
rect 14933 23137 14967 23171
rect 14967 23137 14976 23171
rect 14924 23128 14976 23137
rect 15660 23128 15712 23180
rect 17040 23128 17092 23180
rect 4712 22924 4764 22976
rect 15200 22992 15252 23044
rect 19892 23060 19944 23112
rect 25228 23060 25280 23112
rect 26056 23103 26108 23112
rect 26056 23069 26065 23103
rect 26065 23069 26099 23103
rect 26099 23069 26108 23103
rect 26332 23171 26384 23180
rect 26332 23137 26341 23171
rect 26341 23137 26375 23171
rect 26375 23137 26384 23171
rect 26332 23128 26384 23137
rect 26516 23128 26568 23180
rect 33140 23128 33192 23180
rect 35624 23128 35676 23180
rect 44180 23128 44232 23180
rect 44548 23128 44600 23180
rect 47492 23171 47544 23180
rect 47492 23137 47501 23171
rect 47501 23137 47535 23171
rect 47535 23137 47544 23171
rect 48412 23171 48464 23180
rect 47492 23128 47544 23137
rect 48412 23137 48421 23171
rect 48421 23137 48455 23171
rect 48455 23137 48464 23171
rect 48412 23128 48464 23137
rect 48688 23128 48740 23180
rect 49056 23128 49108 23180
rect 49148 23128 49200 23180
rect 53748 23128 53800 23180
rect 53840 23128 53892 23180
rect 56140 23128 56192 23180
rect 66168 23196 66220 23248
rect 62120 23171 62172 23180
rect 62120 23137 62129 23171
rect 62129 23137 62163 23171
rect 62163 23137 62172 23171
rect 62120 23128 62172 23137
rect 62488 23171 62540 23180
rect 62488 23137 62497 23171
rect 62497 23137 62531 23171
rect 62531 23137 62540 23171
rect 62488 23128 62540 23137
rect 64696 23128 64748 23180
rect 72240 23264 72292 23316
rect 75460 23264 75512 23316
rect 76380 23264 76432 23316
rect 76748 23264 76800 23316
rect 88248 23264 88300 23316
rect 72148 23196 72200 23248
rect 72056 23128 72108 23180
rect 72608 23171 72660 23180
rect 72608 23137 72617 23171
rect 72617 23137 72651 23171
rect 72651 23137 72660 23171
rect 72608 23128 72660 23137
rect 72700 23128 72752 23180
rect 76656 23196 76708 23248
rect 90088 23196 90140 23248
rect 26056 23060 26108 23069
rect 26884 23060 26936 23112
rect 46848 23060 46900 23112
rect 47676 23103 47728 23112
rect 47676 23069 47685 23103
rect 47685 23069 47719 23103
rect 47719 23069 47728 23103
rect 47676 23060 47728 23069
rect 48044 23103 48096 23112
rect 48044 23069 48053 23103
rect 48053 23069 48087 23103
rect 48087 23069 48096 23103
rect 48044 23060 48096 23069
rect 48136 23060 48188 23112
rect 55496 23060 55548 23112
rect 55680 23060 55732 23112
rect 61016 23060 61068 23112
rect 62212 23103 62264 23112
rect 62212 23069 62221 23103
rect 62221 23069 62255 23103
rect 62255 23069 62264 23103
rect 62212 23060 62264 23069
rect 17316 22992 17368 23044
rect 25320 22992 25372 23044
rect 26148 22992 26200 23044
rect 47308 23035 47360 23044
rect 47308 23001 47317 23035
rect 47317 23001 47351 23035
rect 47351 23001 47360 23035
rect 47308 22992 47360 23001
rect 26884 22924 26936 22976
rect 33140 22924 33192 22976
rect 37740 22924 37792 22976
rect 46020 22924 46072 22976
rect 46388 22924 46440 22976
rect 46848 22924 46900 22976
rect 49332 22992 49384 23044
rect 49792 22992 49844 23044
rect 62580 23060 62632 23112
rect 67180 23060 67232 23112
rect 67456 23103 67508 23112
rect 67456 23069 67465 23103
rect 67465 23069 67499 23103
rect 67499 23069 67508 23103
rect 67456 23060 67508 23069
rect 67640 23060 67692 23112
rect 71964 23060 72016 23112
rect 62856 22992 62908 23044
rect 63684 22992 63736 23044
rect 64420 22992 64472 23044
rect 66536 22992 66588 23044
rect 48504 22924 48556 22976
rect 48780 22924 48832 22976
rect 53840 22924 53892 22976
rect 53932 22924 53984 22976
rect 55128 22924 55180 22976
rect 55496 22924 55548 22976
rect 56232 22924 56284 22976
rect 62764 22924 62816 22976
rect 65248 22924 65300 22976
rect 71044 22992 71096 23044
rect 71688 22992 71740 23044
rect 72240 22992 72292 23044
rect 72424 22992 72476 23044
rect 69112 22924 69164 22976
rect 70492 22924 70544 22976
rect 81900 23128 81952 23180
rect 89352 23128 89404 23180
rect 73436 23060 73488 23112
rect 74356 23060 74408 23112
rect 91100 23060 91152 23112
rect 93400 22992 93452 23044
rect 74448 22924 74500 22976
rect 78772 22924 78824 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 65686 22822 65738 22874
rect 65750 22822 65802 22874
rect 65814 22822 65866 22874
rect 65878 22822 65930 22874
rect 96406 22822 96458 22874
rect 96470 22822 96522 22874
rect 96534 22822 96586 22874
rect 96598 22822 96650 22874
rect 15016 22720 15068 22772
rect 17224 22720 17276 22772
rect 26332 22720 26384 22772
rect 37740 22720 37792 22772
rect 47676 22720 47728 22772
rect 48320 22720 48372 22772
rect 48504 22720 48556 22772
rect 49884 22720 49936 22772
rect 55680 22720 55732 22772
rect 56048 22720 56100 22772
rect 2044 22652 2096 22704
rect 15108 22652 15160 22704
rect 15200 22652 15252 22704
rect 27160 22652 27212 22704
rect 33416 22652 33468 22704
rect 11244 22584 11296 22636
rect 11704 22584 11756 22636
rect 17316 22584 17368 22636
rect 23756 22584 23808 22636
rect 33600 22584 33652 22636
rect 36452 22652 36504 22704
rect 64788 22652 64840 22704
rect 65432 22652 65484 22704
rect 33876 22584 33928 22636
rect 64420 22584 64472 22636
rect 64972 22627 65024 22636
rect 64972 22593 64981 22627
rect 64981 22593 65015 22627
rect 65015 22593 65024 22627
rect 64972 22584 65024 22593
rect 65064 22584 65116 22636
rect 71412 22720 71464 22772
rect 95792 22720 95844 22772
rect 73804 22652 73856 22704
rect 12992 22516 13044 22568
rect 43996 22516 44048 22568
rect 55312 22516 55364 22568
rect 58808 22516 58860 22568
rect 62672 22516 62724 22568
rect 63132 22516 63184 22568
rect 65248 22516 65300 22568
rect 65432 22559 65484 22568
rect 65432 22525 65441 22559
rect 65441 22525 65475 22559
rect 65475 22525 65484 22559
rect 65708 22559 65760 22568
rect 65432 22516 65484 22525
rect 65708 22525 65717 22559
rect 65717 22525 65751 22559
rect 65751 22525 65760 22559
rect 65708 22516 65760 22525
rect 66536 22584 66588 22636
rect 74448 22584 74500 22636
rect 75460 22584 75512 22636
rect 74632 22516 74684 22568
rect 75552 22516 75604 22568
rect 76104 22559 76156 22568
rect 76104 22525 76113 22559
rect 76113 22525 76147 22559
rect 76147 22525 76156 22559
rect 76104 22516 76156 22525
rect 12716 22448 12768 22500
rect 15108 22448 15160 22500
rect 15660 22448 15712 22500
rect 19248 22448 19300 22500
rect 25228 22448 25280 22500
rect 16488 22380 16540 22432
rect 33416 22380 33468 22432
rect 35256 22423 35308 22432
rect 35256 22389 35265 22423
rect 35265 22389 35299 22423
rect 35299 22389 35308 22423
rect 35256 22380 35308 22389
rect 48780 22380 48832 22432
rect 50712 22380 50764 22432
rect 54668 22380 54720 22432
rect 55128 22380 55180 22432
rect 64696 22380 64748 22432
rect 65064 22448 65116 22500
rect 96896 22448 96948 22500
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 50326 22278 50378 22330
rect 50390 22278 50442 22330
rect 50454 22278 50506 22330
rect 50518 22278 50570 22330
rect 81046 22278 81098 22330
rect 81110 22278 81162 22330
rect 81174 22278 81226 22330
rect 81238 22278 81290 22330
rect 20444 22176 20496 22228
rect 26884 22176 26936 22228
rect 29920 22176 29972 22228
rect 11428 22108 11480 22160
rect 13544 22108 13596 22160
rect 21088 22108 21140 22160
rect 25596 22108 25648 22160
rect 26240 22108 26292 22160
rect 33048 22108 33100 22160
rect 33416 22176 33468 22228
rect 35256 22176 35308 22228
rect 38568 22176 38620 22228
rect 95884 22176 95936 22228
rect 36452 22108 36504 22160
rect 37648 22108 37700 22160
rect 9864 22083 9916 22092
rect 9864 22049 9873 22083
rect 9873 22049 9907 22083
rect 9907 22049 9916 22083
rect 9864 22040 9916 22049
rect 17316 22040 17368 22092
rect 30196 22040 30248 22092
rect 38200 22040 38252 22092
rect 38476 22083 38528 22092
rect 17132 21972 17184 22024
rect 24124 21972 24176 22024
rect 38476 22049 38485 22083
rect 38485 22049 38519 22083
rect 38519 22049 38528 22083
rect 46848 22108 46900 22160
rect 52368 22108 52420 22160
rect 54668 22108 54720 22160
rect 64604 22108 64656 22160
rect 64788 22108 64840 22160
rect 70492 22108 70544 22160
rect 38476 22040 38528 22049
rect 40040 22040 40092 22092
rect 40500 22040 40552 22092
rect 43812 22083 43864 22092
rect 25596 21904 25648 21956
rect 29000 21904 29052 21956
rect 38384 21904 38436 21956
rect 42156 21972 42208 22024
rect 6184 21836 6236 21888
rect 37924 21836 37976 21888
rect 38200 21836 38252 21888
rect 41512 21836 41564 21888
rect 43812 22049 43821 22083
rect 43821 22049 43855 22083
rect 43855 22049 43864 22083
rect 43812 22040 43864 22049
rect 46756 22040 46808 22092
rect 52644 22040 52696 22092
rect 55496 22040 55548 22092
rect 55772 22040 55824 22092
rect 46204 21972 46256 22024
rect 46296 21972 46348 22024
rect 51724 21972 51776 22024
rect 53104 21972 53156 22024
rect 73436 22040 73488 22092
rect 75368 22083 75420 22092
rect 75368 22049 75377 22083
rect 75377 22049 75411 22083
rect 75411 22049 75420 22083
rect 75368 22040 75420 22049
rect 75920 22040 75972 22092
rect 76012 21972 76064 22024
rect 85488 22040 85540 22092
rect 85304 22015 85356 22024
rect 85304 21981 85313 22015
rect 85313 21981 85347 22015
rect 85347 21981 85356 22015
rect 85304 21972 85356 21981
rect 56140 21904 56192 21956
rect 46296 21836 46348 21888
rect 51724 21836 51776 21888
rect 53104 21836 53156 21888
rect 53196 21836 53248 21888
rect 56968 21836 57020 21888
rect 58624 21879 58676 21888
rect 58624 21845 58633 21879
rect 58633 21845 58667 21879
rect 58667 21845 58676 21879
rect 58624 21836 58676 21845
rect 58900 21904 58952 21956
rect 60832 21904 60884 21956
rect 62672 21904 62724 21956
rect 88248 21904 88300 21956
rect 92848 21904 92900 21956
rect 85120 21836 85172 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 65686 21734 65738 21786
rect 65750 21734 65802 21786
rect 65814 21734 65866 21786
rect 65878 21734 65930 21786
rect 96406 21734 96458 21786
rect 96470 21734 96522 21786
rect 96534 21734 96586 21786
rect 96598 21734 96650 21786
rect 17408 21632 17460 21684
rect 17776 21632 17828 21684
rect 5448 21564 5500 21616
rect 17316 21564 17368 21616
rect 2412 21496 2464 21548
rect 25872 21564 25924 21616
rect 28908 21564 28960 21616
rect 32864 21607 32916 21616
rect 32864 21573 32873 21607
rect 32873 21573 32907 21607
rect 32907 21573 32916 21607
rect 32864 21564 32916 21573
rect 34060 21564 34112 21616
rect 37096 21564 37148 21616
rect 37372 21564 37424 21616
rect 40040 21564 40092 21616
rect 42248 21564 42300 21616
rect 50896 21632 50948 21684
rect 43996 21607 44048 21616
rect 43996 21573 44005 21607
rect 44005 21573 44039 21607
rect 44039 21573 44048 21607
rect 43996 21564 44048 21573
rect 44548 21564 44600 21616
rect 51356 21632 51408 21684
rect 25412 21496 25464 21548
rect 12072 21471 12124 21480
rect 12072 21437 12081 21471
rect 12081 21437 12115 21471
rect 12115 21437 12124 21471
rect 12072 21428 12124 21437
rect 12164 21428 12216 21480
rect 12624 21471 12676 21480
rect 12624 21437 12633 21471
rect 12633 21437 12667 21471
rect 12667 21437 12676 21471
rect 12624 21428 12676 21437
rect 12808 21471 12860 21480
rect 12808 21437 12817 21471
rect 12817 21437 12851 21471
rect 12851 21437 12860 21471
rect 12808 21428 12860 21437
rect 17132 21428 17184 21480
rect 25872 21471 25924 21480
rect 25872 21437 25881 21471
rect 25881 21437 25915 21471
rect 25915 21437 25924 21471
rect 25872 21428 25924 21437
rect 32220 21496 32272 21548
rect 34796 21496 34848 21548
rect 35348 21496 35400 21548
rect 55036 21632 55088 21684
rect 62672 21632 62724 21684
rect 66260 21632 66312 21684
rect 85488 21632 85540 21684
rect 60832 21564 60884 21616
rect 52276 21539 52328 21548
rect 26148 21471 26200 21480
rect 26148 21437 26157 21471
rect 26157 21437 26191 21471
rect 26191 21437 26200 21471
rect 26148 21428 26200 21437
rect 17224 21360 17276 21412
rect 17500 21360 17552 21412
rect 25596 21360 25648 21412
rect 26332 21428 26384 21480
rect 38568 21428 38620 21480
rect 26884 21360 26936 21412
rect 27804 21360 27856 21412
rect 33784 21360 33836 21412
rect 38752 21428 38804 21480
rect 39396 21428 39448 21480
rect 16304 21292 16356 21344
rect 26240 21292 26292 21344
rect 35256 21292 35308 21344
rect 35716 21292 35768 21344
rect 37924 21292 37976 21344
rect 38476 21292 38528 21344
rect 41420 21471 41472 21480
rect 41420 21437 41429 21471
rect 41429 21437 41463 21471
rect 41463 21437 41472 21471
rect 41420 21428 41472 21437
rect 46204 21428 46256 21480
rect 52276 21505 52285 21539
rect 52285 21505 52319 21539
rect 52319 21505 52328 21539
rect 52276 21496 52328 21505
rect 41512 21360 41564 21412
rect 44088 21360 44140 21412
rect 49240 21360 49292 21412
rect 50160 21360 50212 21412
rect 52184 21471 52236 21480
rect 52184 21437 52193 21471
rect 52193 21437 52227 21471
rect 52227 21437 52236 21471
rect 52552 21496 52604 21548
rect 54024 21539 54076 21548
rect 54024 21505 54033 21539
rect 54033 21505 54067 21539
rect 54067 21505 54076 21539
rect 54024 21496 54076 21505
rect 54392 21496 54444 21548
rect 58624 21496 58676 21548
rect 58992 21496 59044 21548
rect 52184 21428 52236 21437
rect 53748 21428 53800 21480
rect 55680 21471 55732 21480
rect 55680 21437 55689 21471
rect 55689 21437 55723 21471
rect 55723 21437 55732 21471
rect 55680 21428 55732 21437
rect 59360 21428 59412 21480
rect 60464 21428 60516 21480
rect 60832 21471 60884 21480
rect 60832 21437 60841 21471
rect 60841 21437 60875 21471
rect 60875 21437 60884 21471
rect 60832 21428 60884 21437
rect 61016 21564 61068 21616
rect 61108 21564 61160 21616
rect 77944 21564 77996 21616
rect 80704 21564 80756 21616
rect 86316 21564 86368 21616
rect 61844 21496 61896 21548
rect 64420 21496 64472 21548
rect 65156 21539 65208 21548
rect 65156 21505 65165 21539
rect 65165 21505 65199 21539
rect 65199 21505 65208 21539
rect 65156 21496 65208 21505
rect 65248 21496 65300 21548
rect 78036 21496 78088 21548
rect 78128 21496 78180 21548
rect 93860 21496 93912 21548
rect 53196 21360 53248 21412
rect 55036 21360 55088 21412
rect 61568 21428 61620 21480
rect 80704 21428 80756 21480
rect 82452 21428 82504 21480
rect 62580 21360 62632 21412
rect 62672 21360 62724 21412
rect 90640 21360 90692 21412
rect 38752 21292 38804 21344
rect 40408 21292 40460 21344
rect 42892 21292 42944 21344
rect 48688 21292 48740 21344
rect 50620 21292 50672 21344
rect 52276 21292 52328 21344
rect 52736 21292 52788 21344
rect 55864 21292 55916 21344
rect 61292 21292 61344 21344
rect 62948 21292 63000 21344
rect 63592 21292 63644 21344
rect 66260 21292 66312 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 50326 21190 50378 21242
rect 50390 21190 50442 21242
rect 50454 21190 50506 21242
rect 50518 21190 50570 21242
rect 81046 21190 81098 21242
rect 81110 21190 81162 21242
rect 81174 21190 81226 21242
rect 81238 21190 81290 21242
rect 1860 21131 1912 21140
rect 1860 21097 1869 21131
rect 1869 21097 1903 21131
rect 1903 21097 1912 21131
rect 1860 21088 1912 21097
rect 17500 21131 17552 21140
rect 6184 21063 6236 21072
rect 2412 20952 2464 21004
rect 4896 20952 4948 21004
rect 5448 20995 5500 21004
rect 5448 20961 5457 20995
rect 5457 20961 5491 20995
rect 5491 20961 5500 20995
rect 5448 20952 5500 20961
rect 5908 20952 5960 21004
rect 6184 21029 6193 21063
rect 6193 21029 6227 21063
rect 6227 21029 6236 21063
rect 6184 21020 6236 21029
rect 17500 21097 17509 21131
rect 17509 21097 17543 21131
rect 17543 21097 17552 21131
rect 17500 21088 17552 21097
rect 26148 21088 26200 21140
rect 42800 21088 42852 21140
rect 42892 21088 42944 21140
rect 47676 21088 47728 21140
rect 51356 21088 51408 21140
rect 55864 21088 55916 21140
rect 18788 21020 18840 21072
rect 58900 21088 58952 21140
rect 58992 21088 59044 21140
rect 81532 21088 81584 21140
rect 57428 21020 57480 21072
rect 61844 21020 61896 21072
rect 14556 20952 14608 21004
rect 15936 20995 15988 21004
rect 15936 20961 15945 20995
rect 15945 20961 15979 20995
rect 15979 20961 15988 20995
rect 15936 20952 15988 20961
rect 17960 20952 18012 21004
rect 26056 20952 26108 21004
rect 45928 20952 45980 21004
rect 46112 20952 46164 21004
rect 51080 20952 51132 21004
rect 51172 20952 51224 21004
rect 63224 20995 63276 21004
rect 63224 20961 63233 20995
rect 63233 20961 63267 20995
rect 63267 20961 63276 20995
rect 63224 20952 63276 20961
rect 63684 20952 63736 21004
rect 67364 20995 67416 21004
rect 67364 20961 67373 20995
rect 67373 20961 67407 20995
rect 67407 20961 67416 20995
rect 67364 20952 67416 20961
rect 72148 21020 72200 21072
rect 73712 21020 73764 21072
rect 75644 20952 75696 21004
rect 84200 21088 84252 21140
rect 3424 20816 3476 20868
rect 5632 20927 5684 20936
rect 5632 20893 5641 20927
rect 5641 20893 5675 20927
rect 5675 20893 5684 20927
rect 5632 20884 5684 20893
rect 6184 20884 6236 20936
rect 15752 20884 15804 20936
rect 5540 20816 5592 20868
rect 5908 20816 5960 20868
rect 8116 20816 8168 20868
rect 6644 20748 6696 20800
rect 11060 20748 11112 20800
rect 12164 20748 12216 20800
rect 14740 20748 14792 20800
rect 26792 20884 26844 20936
rect 29000 20884 29052 20936
rect 30104 20884 30156 20936
rect 35256 20884 35308 20936
rect 17132 20816 17184 20868
rect 17500 20816 17552 20868
rect 21732 20816 21784 20868
rect 38384 20816 38436 20868
rect 42800 20884 42852 20936
rect 44088 20884 44140 20936
rect 44548 20927 44600 20936
rect 44548 20893 44557 20927
rect 44557 20893 44591 20927
rect 44591 20893 44600 20927
rect 44548 20884 44600 20893
rect 78036 20884 78088 20936
rect 80060 20927 80112 20936
rect 80060 20893 80069 20927
rect 80069 20893 80103 20927
rect 80103 20893 80112 20927
rect 80060 20884 80112 20893
rect 45928 20816 45980 20868
rect 46940 20816 46992 20868
rect 47952 20816 48004 20868
rect 50896 20816 50948 20868
rect 51080 20816 51132 20868
rect 55680 20816 55732 20868
rect 55864 20816 55916 20868
rect 60556 20816 60608 20868
rect 17224 20748 17276 20800
rect 29092 20748 29144 20800
rect 35900 20748 35952 20800
rect 37004 20748 37056 20800
rect 37924 20748 37976 20800
rect 38292 20748 38344 20800
rect 38752 20748 38804 20800
rect 62856 20748 62908 20800
rect 64144 20791 64196 20800
rect 64144 20757 64153 20791
rect 64153 20757 64187 20791
rect 64187 20757 64196 20791
rect 64144 20748 64196 20757
rect 64420 20748 64472 20800
rect 65064 20748 65116 20800
rect 65156 20748 65208 20800
rect 67456 20748 67508 20800
rect 72700 20816 72752 20868
rect 76656 20816 76708 20868
rect 85580 21020 85632 21072
rect 95884 21020 95936 21072
rect 93584 20952 93636 21004
rect 92940 20884 92992 20936
rect 92756 20791 92808 20800
rect 92756 20757 92765 20791
rect 92765 20757 92799 20791
rect 92799 20757 92808 20791
rect 92756 20748 92808 20757
rect 93584 20748 93636 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 65686 20646 65738 20698
rect 65750 20646 65802 20698
rect 65814 20646 65866 20698
rect 65878 20646 65930 20698
rect 96406 20646 96458 20698
rect 96470 20646 96522 20698
rect 96534 20646 96586 20698
rect 96598 20646 96650 20698
rect 2964 20544 3016 20596
rect 22468 20544 22520 20596
rect 22744 20587 22796 20596
rect 22744 20553 22753 20587
rect 22753 20553 22787 20587
rect 22787 20553 22796 20587
rect 22744 20544 22796 20553
rect 23020 20544 23072 20596
rect 44088 20544 44140 20596
rect 44640 20544 44692 20596
rect 46112 20544 46164 20596
rect 16856 20476 16908 20528
rect 51908 20544 51960 20596
rect 53932 20544 53984 20596
rect 54024 20544 54076 20596
rect 81624 20544 81676 20596
rect 93308 20544 93360 20596
rect 64512 20476 64564 20528
rect 70584 20519 70636 20528
rect 5540 20408 5592 20460
rect 6276 20408 6328 20460
rect 22468 20408 22520 20460
rect 23020 20408 23072 20460
rect 33692 20408 33744 20460
rect 15844 20272 15896 20324
rect 34060 20272 34112 20324
rect 12808 20204 12860 20256
rect 23204 20204 23256 20256
rect 26608 20204 26660 20256
rect 27160 20204 27212 20256
rect 27252 20204 27304 20256
rect 34152 20204 34204 20256
rect 38844 20340 38896 20392
rect 39028 20340 39080 20392
rect 34704 20272 34756 20324
rect 45284 20340 45336 20392
rect 46940 20408 46992 20460
rect 52276 20408 52328 20460
rect 53104 20408 53156 20460
rect 45468 20340 45520 20392
rect 51908 20340 51960 20392
rect 54116 20340 54168 20392
rect 54484 20408 54536 20460
rect 58900 20408 58952 20460
rect 59728 20408 59780 20460
rect 62764 20408 62816 20460
rect 63684 20408 63736 20460
rect 63960 20340 64012 20392
rect 65156 20340 65208 20392
rect 65248 20340 65300 20392
rect 70216 20451 70268 20460
rect 70216 20417 70225 20451
rect 70225 20417 70259 20451
rect 70259 20417 70268 20451
rect 70216 20408 70268 20417
rect 70584 20485 70593 20519
rect 70593 20485 70627 20519
rect 70627 20485 70636 20519
rect 70584 20476 70636 20485
rect 71780 20519 71832 20528
rect 71780 20485 71789 20519
rect 71789 20485 71823 20519
rect 71823 20485 71832 20519
rect 71780 20476 71832 20485
rect 73160 20476 73212 20528
rect 72700 20451 72752 20460
rect 72700 20417 72709 20451
rect 72709 20417 72743 20451
rect 72743 20417 72752 20451
rect 72700 20408 72752 20417
rect 73068 20408 73120 20460
rect 81716 20476 81768 20528
rect 81900 20476 81952 20528
rect 93952 20476 94004 20528
rect 94596 20476 94648 20528
rect 95148 20476 95200 20528
rect 69756 20340 69808 20392
rect 69940 20340 69992 20392
rect 70124 20383 70176 20392
rect 70124 20349 70133 20383
rect 70133 20349 70167 20383
rect 70167 20349 70176 20383
rect 70124 20340 70176 20349
rect 70768 20340 70820 20392
rect 71136 20340 71188 20392
rect 72148 20383 72200 20392
rect 72148 20349 72157 20383
rect 72157 20349 72191 20383
rect 72191 20349 72200 20383
rect 72148 20340 72200 20349
rect 72608 20340 72660 20392
rect 72884 20383 72936 20392
rect 72884 20349 72893 20383
rect 72893 20349 72927 20383
rect 72927 20349 72936 20383
rect 72884 20340 72936 20349
rect 72976 20340 73028 20392
rect 80980 20408 81032 20460
rect 82268 20408 82320 20460
rect 81532 20340 81584 20392
rect 81716 20340 81768 20392
rect 81900 20340 81952 20392
rect 82084 20383 82136 20392
rect 82084 20349 82093 20383
rect 82093 20349 82127 20383
rect 82127 20349 82136 20383
rect 82084 20340 82136 20349
rect 82176 20383 82228 20392
rect 82176 20349 82186 20383
rect 82186 20349 82220 20383
rect 82220 20349 82228 20383
rect 82360 20383 82412 20392
rect 82176 20340 82228 20349
rect 82360 20349 82369 20383
rect 82369 20349 82403 20383
rect 82403 20349 82412 20383
rect 82360 20340 82412 20349
rect 89536 20340 89588 20392
rect 93676 20383 93728 20392
rect 93676 20349 93685 20383
rect 93685 20349 93719 20383
rect 93719 20349 93728 20383
rect 93676 20340 93728 20349
rect 52276 20315 52328 20324
rect 52276 20281 52285 20315
rect 52285 20281 52319 20315
rect 52319 20281 52328 20315
rect 52276 20272 52328 20281
rect 52460 20272 52512 20324
rect 53932 20272 53984 20324
rect 64788 20315 64840 20324
rect 44640 20204 44692 20256
rect 45100 20204 45152 20256
rect 45284 20204 45336 20256
rect 46211 20204 46263 20256
rect 54116 20204 54168 20256
rect 64052 20204 64104 20256
rect 64788 20281 64822 20315
rect 64822 20281 64840 20315
rect 64788 20272 64840 20281
rect 79048 20272 79100 20324
rect 65064 20204 65116 20256
rect 65984 20204 66036 20256
rect 70860 20204 70912 20256
rect 71136 20204 71188 20256
rect 71780 20204 71832 20256
rect 73160 20204 73212 20256
rect 81808 20204 81860 20256
rect 92848 20272 92900 20324
rect 93952 20340 94004 20392
rect 92296 20204 92348 20256
rect 92664 20204 92716 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 50326 20102 50378 20154
rect 50390 20102 50442 20154
rect 50454 20102 50506 20154
rect 50518 20102 50570 20154
rect 81046 20102 81098 20154
rect 81110 20102 81162 20154
rect 81174 20102 81226 20154
rect 81238 20102 81290 20154
rect 3240 20000 3292 20052
rect 34060 20000 34112 20052
rect 34152 20000 34204 20052
rect 3792 19932 3844 19984
rect 19248 19932 19300 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 9404 19864 9456 19916
rect 18144 19864 18196 19916
rect 20168 19796 20220 19848
rect 33692 19932 33744 19984
rect 26424 19864 26476 19916
rect 26884 19864 26936 19916
rect 27252 19864 27304 19916
rect 27528 19864 27580 19916
rect 26976 19796 27028 19848
rect 29092 19839 29144 19848
rect 29092 19805 29101 19839
rect 29101 19805 29135 19839
rect 29135 19805 29144 19839
rect 29092 19796 29144 19805
rect 38568 20000 38620 20052
rect 44088 20000 44140 20052
rect 48320 20000 48372 20052
rect 48596 20000 48648 20052
rect 78680 20000 78732 20052
rect 91836 20000 91888 20052
rect 97632 20043 97684 20052
rect 97632 20009 97641 20043
rect 97641 20009 97675 20043
rect 97675 20009 97684 20043
rect 97632 20000 97684 20009
rect 38752 19864 38804 19916
rect 45468 19864 45520 19916
rect 46940 19864 46992 19916
rect 48320 19864 48372 19916
rect 48780 19907 48832 19916
rect 48780 19873 48789 19907
rect 48789 19873 48823 19907
rect 48823 19873 48832 19907
rect 48780 19864 48832 19873
rect 54208 19932 54260 19984
rect 56600 19932 56652 19984
rect 54484 19864 54536 19916
rect 54668 19907 54720 19916
rect 54668 19873 54677 19907
rect 54677 19873 54711 19907
rect 54711 19873 54720 19907
rect 54668 19864 54720 19873
rect 55128 19864 55180 19916
rect 55680 19864 55732 19916
rect 59728 19932 59780 19984
rect 43444 19796 43496 19848
rect 12072 19728 12124 19780
rect 36268 19728 36320 19780
rect 27160 19660 27212 19712
rect 34796 19660 34848 19712
rect 38660 19728 38712 19780
rect 39028 19728 39080 19780
rect 46204 19728 46256 19780
rect 46296 19728 46348 19780
rect 47768 19728 47820 19780
rect 61752 19864 61804 19916
rect 53472 19728 53524 19780
rect 62948 19796 63000 19848
rect 63224 19796 63276 19848
rect 73068 19932 73120 19984
rect 73988 19907 74040 19916
rect 73988 19873 73997 19907
rect 73997 19873 74031 19907
rect 74031 19873 74040 19907
rect 73988 19864 74040 19873
rect 74632 19864 74684 19916
rect 75644 19907 75696 19916
rect 75644 19873 75653 19907
rect 75653 19873 75687 19907
rect 75687 19873 75696 19907
rect 75644 19864 75696 19873
rect 75828 19907 75880 19916
rect 75828 19873 75837 19907
rect 75837 19873 75871 19907
rect 75871 19873 75880 19907
rect 75828 19864 75880 19873
rect 97540 19975 97592 19984
rect 97540 19941 97549 19975
rect 97549 19941 97583 19975
rect 97583 19941 97592 19975
rect 97540 19932 97592 19941
rect 86960 19864 87012 19916
rect 76288 19796 76340 19848
rect 63960 19728 64012 19780
rect 87696 19728 87748 19780
rect 43904 19660 43956 19712
rect 43996 19660 44048 19712
rect 50160 19660 50212 19712
rect 55036 19660 55088 19712
rect 57520 19660 57572 19712
rect 59360 19660 59412 19712
rect 60924 19660 60976 19712
rect 61108 19660 61160 19712
rect 63776 19660 63828 19712
rect 71228 19660 71280 19712
rect 71688 19660 71740 19712
rect 71780 19660 71832 19712
rect 75736 19660 75788 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 65686 19558 65738 19610
rect 65750 19558 65802 19610
rect 65814 19558 65866 19610
rect 65878 19558 65930 19610
rect 96406 19558 96458 19610
rect 96470 19558 96522 19610
rect 96534 19558 96586 19610
rect 96598 19558 96650 19610
rect 21916 19456 21968 19508
rect 50436 19456 50488 19508
rect 52276 19456 52328 19508
rect 73988 19456 74040 19508
rect 18052 19388 18104 19440
rect 34796 19388 34848 19440
rect 34888 19388 34940 19440
rect 6736 19320 6788 19372
rect 33692 19320 33744 19372
rect 4988 19252 5040 19304
rect 27344 19252 27396 19304
rect 35900 19295 35952 19304
rect 35900 19261 35909 19295
rect 35909 19261 35943 19295
rect 35943 19261 35952 19295
rect 35900 19252 35952 19261
rect 36084 19295 36136 19304
rect 36084 19261 36092 19295
rect 36092 19261 36126 19295
rect 36126 19261 36136 19295
rect 36084 19252 36136 19261
rect 36268 19388 36320 19440
rect 44088 19388 44140 19440
rect 36636 19320 36688 19372
rect 45100 19388 45152 19440
rect 46112 19388 46164 19440
rect 47860 19388 47912 19440
rect 36360 19252 36412 19304
rect 36544 19252 36596 19304
rect 36912 19252 36964 19304
rect 45468 19320 45520 19372
rect 48596 19320 48648 19372
rect 50068 19320 50120 19372
rect 52644 19388 52696 19440
rect 56508 19388 56560 19440
rect 56600 19388 56652 19440
rect 57428 19388 57480 19440
rect 57520 19388 57572 19440
rect 61936 19388 61988 19440
rect 64604 19388 64656 19440
rect 67272 19388 67324 19440
rect 69480 19388 69532 19440
rect 72976 19388 73028 19440
rect 60740 19320 60792 19372
rect 60832 19320 60884 19372
rect 45836 19295 45888 19304
rect 5540 19184 5592 19236
rect 21640 19184 21692 19236
rect 23020 19184 23072 19236
rect 34704 19184 34756 19236
rect 35808 19184 35860 19236
rect 10140 19116 10192 19168
rect 22468 19116 22520 19168
rect 22744 19116 22796 19168
rect 30840 19116 30892 19168
rect 36728 19184 36780 19236
rect 43444 19184 43496 19236
rect 36636 19116 36688 19168
rect 44088 19116 44140 19168
rect 44640 19116 44692 19168
rect 45836 19261 45845 19295
rect 45845 19261 45879 19295
rect 45879 19261 45888 19295
rect 45836 19252 45888 19261
rect 46204 19252 46256 19304
rect 46940 19252 46992 19304
rect 47952 19252 48004 19304
rect 50252 19295 50304 19304
rect 50252 19261 50261 19295
rect 50261 19261 50295 19295
rect 50295 19261 50304 19295
rect 50252 19252 50304 19261
rect 50436 19295 50488 19304
rect 50436 19261 50445 19295
rect 50445 19261 50479 19295
rect 50479 19261 50488 19295
rect 50436 19252 50488 19261
rect 50620 19295 50672 19304
rect 50620 19261 50629 19295
rect 50629 19261 50663 19295
rect 50663 19261 50672 19295
rect 50620 19252 50672 19261
rect 50804 19295 50856 19304
rect 50804 19261 50813 19295
rect 50813 19261 50847 19295
rect 50847 19261 50856 19295
rect 50804 19252 50856 19261
rect 58440 19252 58492 19304
rect 58624 19252 58676 19304
rect 60372 19252 60424 19304
rect 50804 19116 50856 19168
rect 51264 19184 51316 19236
rect 52644 19227 52696 19236
rect 52644 19193 52653 19227
rect 52653 19193 52687 19227
rect 52687 19193 52696 19227
rect 52644 19184 52696 19193
rect 60648 19184 60700 19236
rect 51080 19116 51132 19168
rect 51172 19116 51224 19168
rect 54760 19116 54812 19168
rect 55864 19116 55916 19168
rect 60740 19116 60792 19168
rect 61108 19252 61160 19304
rect 71872 19320 71924 19372
rect 72608 19320 72660 19372
rect 98368 19320 98420 19372
rect 73252 19252 73304 19304
rect 63224 19184 63276 19236
rect 69020 19116 69072 19168
rect 75920 19116 75972 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 50326 19014 50378 19066
rect 50390 19014 50442 19066
rect 50454 19014 50506 19066
rect 50518 19014 50570 19066
rect 81046 19014 81098 19066
rect 81110 19014 81162 19066
rect 81174 19014 81226 19066
rect 81238 19014 81290 19066
rect 5632 18912 5684 18964
rect 6828 18844 6880 18896
rect 13544 18912 13596 18964
rect 17316 18912 17368 18964
rect 35808 18912 35860 18964
rect 36728 18912 36780 18964
rect 39028 18912 39080 18964
rect 44548 18912 44600 18964
rect 45468 18912 45520 18964
rect 46296 18912 46348 18964
rect 55864 18912 55916 18964
rect 56416 18912 56468 18964
rect 59360 18912 59412 18964
rect 59452 18912 59504 18964
rect 62120 18912 62172 18964
rect 62396 18912 62448 18964
rect 76104 18912 76156 18964
rect 8208 18776 8260 18828
rect 60832 18844 60884 18896
rect 63408 18844 63460 18896
rect 63500 18844 63552 18896
rect 69296 18844 69348 18896
rect 72424 18844 72476 18896
rect 82084 18844 82136 18896
rect 33600 18776 33652 18828
rect 33692 18776 33744 18828
rect 35256 18776 35308 18828
rect 35808 18776 35860 18828
rect 13820 18708 13872 18760
rect 16304 18708 16356 18760
rect 17960 18708 18012 18760
rect 22652 18708 22704 18760
rect 25228 18708 25280 18760
rect 25320 18708 25372 18760
rect 25688 18708 25740 18760
rect 26516 18708 26568 18760
rect 26884 18708 26936 18760
rect 36452 18708 36504 18760
rect 36728 18776 36780 18828
rect 40040 18708 40092 18760
rect 41328 18776 41380 18828
rect 47308 18776 47360 18828
rect 50804 18776 50856 18828
rect 53012 18776 53064 18828
rect 53104 18819 53156 18828
rect 53104 18785 53113 18819
rect 53113 18785 53147 18819
rect 53147 18785 53156 18819
rect 53104 18776 53156 18785
rect 56048 18776 56100 18828
rect 59360 18776 59412 18828
rect 59728 18776 59780 18828
rect 59820 18776 59872 18828
rect 69480 18776 69532 18828
rect 69756 18776 69808 18828
rect 70676 18776 70728 18828
rect 70768 18819 70820 18828
rect 70768 18785 70777 18819
rect 70777 18785 70811 18819
rect 70811 18785 70820 18819
rect 70768 18776 70820 18785
rect 70952 18776 71004 18828
rect 71136 18776 71188 18828
rect 72884 18776 72936 18828
rect 78128 18776 78180 18828
rect 1952 18640 2004 18692
rect 5264 18572 5316 18624
rect 8576 18640 8628 18692
rect 17224 18640 17276 18692
rect 40960 18640 41012 18692
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 17132 18572 17184 18624
rect 92480 18708 92532 18760
rect 47124 18572 47176 18624
rect 51724 18572 51776 18624
rect 52276 18615 52328 18624
rect 52276 18581 52285 18615
rect 52285 18581 52319 18615
rect 52319 18581 52328 18615
rect 60832 18640 60884 18692
rect 60924 18640 60976 18692
rect 64512 18640 64564 18692
rect 65524 18640 65576 18692
rect 78220 18640 78272 18692
rect 78312 18640 78364 18692
rect 82728 18640 82780 18692
rect 52276 18572 52328 18581
rect 54852 18572 54904 18624
rect 59820 18572 59872 18624
rect 61936 18572 61988 18624
rect 76288 18572 76340 18624
rect 93952 18572 94004 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 65686 18470 65738 18522
rect 65750 18470 65802 18522
rect 65814 18470 65866 18522
rect 65878 18470 65930 18522
rect 96406 18470 96458 18522
rect 96470 18470 96522 18522
rect 96534 18470 96586 18522
rect 96598 18470 96650 18522
rect 5540 18411 5592 18420
rect 5540 18377 5549 18411
rect 5549 18377 5583 18411
rect 5583 18377 5592 18411
rect 5540 18368 5592 18377
rect 12164 18368 12216 18420
rect 17224 18368 17276 18420
rect 22100 18368 22152 18420
rect 33600 18368 33652 18420
rect 6092 18300 6144 18352
rect 7932 18300 7984 18352
rect 4988 18207 5040 18216
rect 4988 18173 4997 18207
rect 4997 18173 5031 18207
rect 5031 18173 5040 18207
rect 4988 18164 5040 18173
rect 8300 18232 8352 18284
rect 9312 18232 9364 18284
rect 10508 18300 10560 18352
rect 26240 18300 26292 18352
rect 26516 18300 26568 18352
rect 33692 18300 33744 18352
rect 17132 18232 17184 18284
rect 17960 18232 18012 18284
rect 33508 18232 33560 18284
rect 35348 18368 35400 18420
rect 35900 18368 35952 18420
rect 38292 18368 38344 18420
rect 39856 18368 39908 18420
rect 50712 18368 50764 18420
rect 56508 18368 56560 18420
rect 65524 18368 65576 18420
rect 66260 18368 66312 18420
rect 35256 18300 35308 18352
rect 35808 18300 35860 18352
rect 36084 18300 36136 18352
rect 36452 18300 36504 18352
rect 41420 18300 41472 18352
rect 43444 18300 43496 18352
rect 50620 18300 50672 18352
rect 51264 18300 51316 18352
rect 63592 18300 63644 18352
rect 63684 18300 63736 18352
rect 65616 18300 65668 18352
rect 65800 18300 65852 18352
rect 67824 18300 67876 18352
rect 69756 18300 69808 18352
rect 70860 18368 70912 18420
rect 92664 18368 92716 18420
rect 73160 18300 73212 18352
rect 73344 18343 73396 18352
rect 73344 18309 73353 18343
rect 73353 18309 73387 18343
rect 73387 18309 73396 18343
rect 73344 18300 73396 18309
rect 34152 18232 34204 18284
rect 26884 18164 26936 18216
rect 30380 18164 30432 18216
rect 34428 18164 34480 18216
rect 36912 18164 36964 18216
rect 37280 18164 37332 18216
rect 38108 18164 38160 18216
rect 38568 18164 38620 18216
rect 39304 18207 39356 18216
rect 39304 18173 39313 18207
rect 39313 18173 39347 18207
rect 39347 18173 39356 18207
rect 39304 18164 39356 18173
rect 39764 18232 39816 18284
rect 41788 18232 41840 18284
rect 56048 18232 56100 18284
rect 56140 18232 56192 18284
rect 62396 18232 62448 18284
rect 62580 18232 62632 18284
rect 65524 18232 65576 18284
rect 8300 18028 8352 18080
rect 8576 18096 8628 18148
rect 13360 18028 13412 18080
rect 13544 18028 13596 18080
rect 22928 18096 22980 18148
rect 31116 18096 31168 18148
rect 31484 18096 31536 18148
rect 32496 18096 32548 18148
rect 33048 18096 33100 18148
rect 33416 18028 33468 18080
rect 43628 18164 43680 18216
rect 45836 18164 45888 18216
rect 46020 18164 46072 18216
rect 46112 18164 46164 18216
rect 56416 18164 56468 18216
rect 59360 18164 59412 18216
rect 60556 18164 60608 18216
rect 62672 18207 62724 18216
rect 62672 18173 62681 18207
rect 62681 18173 62715 18207
rect 62715 18173 62724 18207
rect 69756 18207 69808 18216
rect 62672 18164 62724 18173
rect 69756 18173 69765 18207
rect 69765 18173 69799 18207
rect 69799 18173 69808 18207
rect 69756 18164 69808 18173
rect 70032 18207 70084 18216
rect 70032 18173 70041 18207
rect 70041 18173 70075 18207
rect 70075 18173 70084 18207
rect 70032 18164 70084 18173
rect 70216 18232 70268 18284
rect 73712 18275 73764 18284
rect 73712 18241 73721 18275
rect 73721 18241 73755 18275
rect 73755 18241 73764 18275
rect 73712 18232 73764 18241
rect 89536 18275 89588 18284
rect 89536 18241 89545 18275
rect 89545 18241 89579 18275
rect 89579 18241 89588 18275
rect 89536 18232 89588 18241
rect 92480 18232 92532 18284
rect 92940 18275 92992 18284
rect 92940 18241 92949 18275
rect 92949 18241 92983 18275
rect 92983 18241 92992 18275
rect 92940 18232 92992 18241
rect 70768 18164 70820 18216
rect 63224 18139 63276 18148
rect 35164 18028 35216 18080
rect 39212 18028 39264 18080
rect 41236 18028 41288 18080
rect 41420 18028 41472 18080
rect 60464 18028 60516 18080
rect 63224 18105 63233 18139
rect 63233 18105 63267 18139
rect 63267 18105 63276 18139
rect 63224 18096 63276 18105
rect 71780 18096 71832 18148
rect 72424 18096 72476 18148
rect 73068 18139 73120 18148
rect 73068 18105 73077 18139
rect 73077 18105 73111 18139
rect 73111 18105 73120 18139
rect 73068 18096 73120 18105
rect 77576 18164 77628 18216
rect 82728 18164 82780 18216
rect 78404 18028 78456 18080
rect 91192 18071 91244 18080
rect 91192 18037 91201 18071
rect 91201 18037 91235 18071
rect 91235 18037 91244 18071
rect 91192 18028 91244 18037
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 50326 17926 50378 17978
rect 50390 17926 50442 17978
rect 50454 17926 50506 17978
rect 50518 17926 50570 17978
rect 81046 17926 81098 17978
rect 81110 17926 81162 17978
rect 81174 17926 81226 17978
rect 81238 17926 81290 17978
rect 16304 17824 16356 17876
rect 19340 17824 19392 17876
rect 23020 17756 23072 17808
rect 40132 17756 40184 17808
rect 42800 17756 42852 17808
rect 43812 17756 43864 17808
rect 45468 17756 45520 17808
rect 45560 17756 45612 17808
rect 46296 17756 46348 17808
rect 46388 17756 46440 17808
rect 49148 17756 49200 17808
rect 2596 17688 2648 17740
rect 2964 17688 3016 17740
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 2412 17663 2464 17672
rect 2412 17629 2421 17663
rect 2421 17629 2455 17663
rect 2455 17629 2464 17663
rect 2412 17620 2464 17629
rect 20352 17688 20404 17740
rect 21824 17620 21876 17672
rect 22652 17688 22704 17740
rect 26884 17688 26936 17740
rect 53656 17688 53708 17740
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 28632 17620 28684 17672
rect 30472 17620 30524 17672
rect 31760 17620 31812 17672
rect 40776 17620 40828 17672
rect 40960 17620 41012 17672
rect 46572 17620 46624 17672
rect 48412 17620 48464 17672
rect 1124 17552 1176 17604
rect 48780 17552 48832 17604
rect 49148 17552 49200 17604
rect 6644 17484 6696 17536
rect 31760 17484 31812 17536
rect 31944 17484 31996 17536
rect 42616 17484 42668 17536
rect 43628 17484 43680 17536
rect 56416 17484 56468 17536
rect 56600 17484 56652 17536
rect 59728 17688 59780 17740
rect 64788 17688 64840 17740
rect 72148 17688 72200 17740
rect 64972 17620 65024 17672
rect 66260 17620 66312 17672
rect 74264 17620 74316 17672
rect 78772 17620 78824 17672
rect 75184 17552 75236 17604
rect 83096 17552 83148 17604
rect 83648 17552 83700 17604
rect 61292 17484 61344 17536
rect 90732 17484 90784 17536
rect 94320 17484 94372 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 65686 17382 65738 17434
rect 65750 17382 65802 17434
rect 65814 17382 65866 17434
rect 65878 17382 65930 17434
rect 96406 17382 96458 17434
rect 96470 17382 96522 17434
rect 96534 17382 96586 17434
rect 96598 17382 96650 17434
rect 2044 17280 2096 17332
rect 2320 17280 2372 17332
rect 8024 17280 8076 17332
rect 28908 17280 28960 17332
rect 2412 17144 2464 17196
rect 23296 17212 23348 17264
rect 25596 17212 25648 17264
rect 25688 17212 25740 17264
rect 29092 17212 29144 17264
rect 33968 17212 34020 17264
rect 17040 17144 17092 17196
rect 22652 17144 22704 17196
rect 31944 17144 31996 17196
rect 32036 17144 32088 17196
rect 25596 17076 25648 17128
rect 34428 17076 34480 17128
rect 34796 17076 34848 17128
rect 36360 17280 36412 17332
rect 40408 17280 40460 17332
rect 75184 17280 75236 17332
rect 77944 17323 77996 17332
rect 77944 17289 77953 17323
rect 77953 17289 77987 17323
rect 77987 17289 77996 17323
rect 77944 17280 77996 17289
rect 78036 17280 78088 17332
rect 93952 17323 94004 17332
rect 93952 17289 93961 17323
rect 93961 17289 93995 17323
rect 93995 17289 94004 17323
rect 93952 17280 94004 17289
rect 94320 17280 94372 17332
rect 35164 17212 35216 17264
rect 40960 17212 41012 17264
rect 41328 17212 41380 17264
rect 43536 17212 43588 17264
rect 45284 17212 45336 17264
rect 48136 17212 48188 17264
rect 35900 17144 35952 17196
rect 46388 17144 46440 17196
rect 46572 17144 46624 17196
rect 72148 17212 72200 17264
rect 72976 17212 73028 17264
rect 78772 17212 78824 17264
rect 50712 17144 50764 17196
rect 57152 17144 57204 17196
rect 64788 17144 64840 17196
rect 69296 17144 69348 17196
rect 69848 17144 69900 17196
rect 35256 17119 35308 17128
rect 35256 17085 35265 17119
rect 35265 17085 35299 17119
rect 35299 17085 35308 17119
rect 35256 17076 35308 17085
rect 7840 17008 7892 17060
rect 8116 17008 8168 17060
rect 32036 17008 32088 17060
rect 45560 17076 45612 17128
rect 46296 17076 46348 17128
rect 51356 17076 51408 17128
rect 56416 17076 56468 17128
rect 57520 17076 57572 17128
rect 58716 17076 58768 17128
rect 78036 17119 78088 17128
rect 78036 17085 78045 17119
rect 78045 17085 78079 17119
rect 78079 17085 78088 17119
rect 78036 17076 78088 17085
rect 78220 17119 78272 17128
rect 78220 17085 78229 17119
rect 78229 17085 78263 17119
rect 78263 17085 78272 17119
rect 78220 17076 78272 17085
rect 78312 17119 78364 17128
rect 78312 17085 78321 17119
rect 78321 17085 78355 17119
rect 78355 17085 78364 17119
rect 78312 17076 78364 17085
rect 78496 17076 78548 17128
rect 83280 17076 83332 17128
rect 87512 17119 87564 17128
rect 87512 17085 87521 17119
rect 87521 17085 87555 17119
rect 87555 17085 87564 17119
rect 87512 17076 87564 17085
rect 11152 16940 11204 16992
rect 34244 16983 34296 16992
rect 34244 16949 34253 16983
rect 34253 16949 34287 16983
rect 34287 16949 34296 16983
rect 34244 16940 34296 16949
rect 35072 16940 35124 16992
rect 45100 17008 45152 17060
rect 49332 17008 49384 17060
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 50326 16838 50378 16890
rect 50390 16838 50442 16890
rect 50454 16838 50506 16890
rect 50518 16838 50570 16890
rect 81046 16838 81098 16890
rect 81110 16838 81162 16890
rect 81174 16838 81226 16890
rect 81238 16838 81290 16890
rect 11612 16736 11664 16788
rect 17132 16736 17184 16788
rect 10324 16668 10376 16720
rect 40224 16736 40276 16788
rect 2964 16600 3016 16652
rect 17040 16600 17092 16652
rect 17132 16600 17184 16652
rect 25596 16668 25648 16720
rect 26976 16668 27028 16720
rect 28816 16711 28868 16720
rect 16396 16464 16448 16516
rect 20996 16600 21048 16652
rect 25688 16600 25740 16652
rect 27988 16643 28040 16652
rect 27988 16609 27997 16643
rect 27997 16609 28031 16643
rect 28031 16609 28040 16643
rect 27988 16600 28040 16609
rect 28816 16677 28825 16711
rect 28825 16677 28859 16711
rect 28859 16677 28868 16711
rect 28816 16668 28868 16677
rect 28908 16668 28960 16720
rect 35808 16668 35860 16720
rect 35900 16668 35952 16720
rect 40040 16668 40092 16720
rect 40960 16668 41012 16720
rect 41144 16668 41196 16720
rect 57980 16736 58032 16788
rect 58532 16736 58584 16788
rect 58716 16736 58768 16788
rect 30472 16600 30524 16652
rect 30564 16600 30616 16652
rect 34244 16600 34296 16652
rect 35624 16600 35676 16652
rect 40408 16600 40460 16652
rect 41052 16643 41104 16652
rect 41052 16609 41061 16643
rect 41061 16609 41095 16643
rect 41095 16609 41104 16643
rect 41052 16600 41104 16609
rect 17224 16396 17276 16448
rect 24124 16532 24176 16584
rect 26128 16575 26180 16584
rect 26128 16541 26151 16575
rect 26151 16541 26180 16575
rect 26128 16532 26180 16541
rect 26516 16532 26568 16584
rect 46388 16668 46440 16720
rect 52828 16668 52880 16720
rect 57152 16711 57204 16720
rect 42432 16600 42484 16652
rect 18328 16464 18380 16516
rect 25688 16464 25740 16516
rect 17776 16396 17828 16448
rect 36268 16464 36320 16516
rect 44824 16532 44876 16584
rect 45284 16532 45336 16584
rect 46940 16600 46992 16652
rect 56508 16600 56560 16652
rect 57152 16677 57161 16711
rect 57161 16677 57195 16711
rect 57195 16677 57204 16711
rect 57152 16668 57204 16677
rect 57520 16668 57572 16720
rect 60096 16668 60148 16720
rect 69388 16736 69440 16788
rect 69848 16736 69900 16788
rect 61292 16668 61344 16720
rect 61844 16668 61896 16720
rect 71964 16668 72016 16720
rect 78496 16668 78548 16720
rect 67732 16643 67784 16652
rect 67732 16609 67741 16643
rect 67741 16609 67775 16643
rect 67775 16609 67784 16643
rect 67732 16600 67784 16609
rect 69756 16600 69808 16652
rect 72976 16600 73028 16652
rect 46572 16532 46624 16584
rect 49148 16532 49200 16584
rect 53748 16532 53800 16584
rect 53840 16532 53892 16584
rect 56048 16464 56100 16516
rect 58072 16532 58124 16584
rect 59084 16532 59136 16584
rect 59176 16532 59228 16584
rect 65064 16532 65116 16584
rect 65248 16532 65300 16584
rect 66168 16532 66220 16584
rect 27344 16396 27396 16448
rect 31760 16396 31812 16448
rect 31944 16396 31996 16448
rect 65524 16396 65576 16448
rect 94044 16464 94096 16516
rect 70768 16396 70820 16448
rect 72700 16396 72752 16448
rect 85488 16396 85540 16448
rect 92020 16396 92072 16448
rect 92388 16396 92440 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 65686 16294 65738 16346
rect 65750 16294 65802 16346
rect 65814 16294 65866 16346
rect 65878 16294 65930 16346
rect 96406 16294 96458 16346
rect 96470 16294 96522 16346
rect 96534 16294 96586 16346
rect 96598 16294 96650 16346
rect 6736 16235 6788 16244
rect 6736 16201 6745 16235
rect 6745 16201 6779 16235
rect 6779 16201 6788 16235
rect 6736 16192 6788 16201
rect 9864 16192 9916 16244
rect 17224 16192 17276 16244
rect 14556 16124 14608 16176
rect 5540 16056 5592 16108
rect 10600 16056 10652 16108
rect 18328 16124 18380 16176
rect 23480 16192 23532 16244
rect 24400 16192 24452 16244
rect 25780 16192 25832 16244
rect 26700 16192 26752 16244
rect 27344 16124 27396 16176
rect 29644 16192 29696 16244
rect 31392 16235 31444 16244
rect 31392 16201 31401 16235
rect 31401 16201 31435 16235
rect 31435 16201 31444 16235
rect 31392 16192 31444 16201
rect 17776 16099 17828 16108
rect 17776 16065 17785 16099
rect 17785 16065 17819 16099
rect 17819 16065 17828 16099
rect 17776 16056 17828 16065
rect 31392 16056 31444 16108
rect 31576 16056 31628 16108
rect 32772 16192 32824 16244
rect 39304 16192 39356 16244
rect 40224 16192 40276 16244
rect 41144 16192 41196 16244
rect 31760 16124 31812 16176
rect 17868 16031 17920 16040
rect 17868 15997 17878 16031
rect 17878 15997 17912 16031
rect 17912 15997 17920 16031
rect 17868 15988 17920 15997
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 19248 15988 19300 16040
rect 25688 15988 25740 16040
rect 31024 15988 31076 16040
rect 32496 16124 32548 16176
rect 34060 16167 34112 16176
rect 34060 16133 34069 16167
rect 34069 16133 34103 16167
rect 34103 16133 34112 16167
rect 34060 16124 34112 16133
rect 35808 16124 35860 16176
rect 38200 16124 38252 16176
rect 32036 16056 32088 16108
rect 48872 16192 48924 16244
rect 53748 16192 53800 16244
rect 58992 16192 59044 16244
rect 62396 16192 62448 16244
rect 64144 16192 64196 16244
rect 65432 16192 65484 16244
rect 66168 16192 66220 16244
rect 66260 16192 66312 16244
rect 44272 16124 44324 16176
rect 44088 16056 44140 16108
rect 32128 16031 32180 16040
rect 32128 15997 32137 16031
rect 32137 15997 32171 16031
rect 32171 15997 32180 16031
rect 32128 15988 32180 15997
rect 34704 15988 34756 16040
rect 37280 15988 37332 16040
rect 53288 15988 53340 16040
rect 53748 16056 53800 16108
rect 53932 16056 53984 16108
rect 54024 16056 54076 16108
rect 55772 16056 55824 16108
rect 56048 16124 56100 16176
rect 62672 16124 62724 16176
rect 65524 16124 65576 16176
rect 70860 16124 70912 16176
rect 63224 16056 63276 16108
rect 65340 16056 65392 16108
rect 73344 16056 73396 16108
rect 80060 16056 80112 16108
rect 85488 16056 85540 16108
rect 56048 15988 56100 16040
rect 56324 16031 56376 16040
rect 56324 15997 56333 16031
rect 56333 15997 56367 16031
rect 56367 15997 56376 16031
rect 56324 15988 56376 15997
rect 56508 15988 56560 16040
rect 59176 15988 59228 16040
rect 59360 15988 59412 16040
rect 69756 15988 69808 16040
rect 17224 15895 17276 15904
rect 17224 15861 17233 15895
rect 17233 15861 17267 15895
rect 17267 15861 17276 15895
rect 17224 15852 17276 15861
rect 18144 15920 18196 15972
rect 31208 15920 31260 15972
rect 31392 15920 31444 15972
rect 21456 15852 21508 15904
rect 26884 15852 26936 15904
rect 32036 15920 32088 15972
rect 73804 15988 73856 16040
rect 93124 15920 93176 15972
rect 97172 15920 97224 15972
rect 31760 15852 31812 15904
rect 65340 15852 65392 15904
rect 65432 15852 65484 15904
rect 70768 15852 70820 15904
rect 70860 15852 70912 15904
rect 72608 15852 72660 15904
rect 75920 15852 75972 15904
rect 77116 15852 77168 15904
rect 84752 15852 84804 15904
rect 91744 15852 91796 15904
rect 97356 15852 97408 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 50326 15750 50378 15802
rect 50390 15750 50442 15802
rect 50454 15750 50506 15802
rect 50518 15750 50570 15802
rect 81046 15750 81098 15802
rect 81110 15750 81162 15802
rect 81174 15750 81226 15802
rect 81238 15750 81290 15802
rect 17500 15648 17552 15700
rect 17868 15648 17920 15700
rect 24400 15648 24452 15700
rect 36084 15648 36136 15700
rect 36268 15648 36320 15700
rect 41052 15648 41104 15700
rect 41328 15648 41380 15700
rect 2964 15580 3016 15632
rect 40224 15580 40276 15632
rect 40316 15580 40368 15632
rect 17316 15555 17368 15564
rect 17316 15521 17325 15555
rect 17325 15521 17359 15555
rect 17359 15521 17368 15555
rect 17316 15512 17368 15521
rect 17592 15555 17644 15564
rect 17592 15521 17601 15555
rect 17601 15521 17635 15555
rect 17635 15521 17644 15555
rect 17592 15512 17644 15521
rect 17684 15555 17736 15564
rect 17684 15521 17693 15555
rect 17693 15521 17727 15555
rect 17727 15521 17736 15555
rect 17868 15555 17920 15564
rect 17684 15512 17736 15521
rect 17868 15521 17877 15555
rect 17877 15521 17911 15555
rect 17911 15521 17920 15555
rect 17868 15512 17920 15521
rect 18420 15555 18472 15564
rect 18420 15521 18429 15555
rect 18429 15521 18463 15555
rect 18463 15521 18472 15555
rect 18420 15512 18472 15521
rect 18788 15555 18840 15564
rect 18788 15521 18797 15555
rect 18797 15521 18831 15555
rect 18831 15521 18840 15555
rect 18788 15512 18840 15521
rect 19340 15512 19392 15564
rect 24032 15512 24084 15564
rect 24124 15512 24176 15564
rect 30196 15512 30248 15564
rect 32128 15512 32180 15564
rect 7196 15444 7248 15496
rect 16396 15444 16448 15496
rect 8116 15376 8168 15428
rect 16304 15376 16356 15428
rect 19432 15444 19484 15496
rect 20444 15444 20496 15496
rect 22928 15444 22980 15496
rect 38660 15512 38712 15564
rect 41788 15648 41840 15700
rect 47492 15580 47544 15632
rect 54024 15648 54076 15700
rect 55864 15648 55916 15700
rect 36084 15444 36136 15496
rect 40408 15444 40460 15496
rect 41512 15555 41564 15564
rect 41512 15521 41521 15555
rect 41521 15521 41555 15555
rect 41555 15521 41564 15555
rect 41512 15512 41564 15521
rect 45376 15512 45428 15564
rect 48780 15555 48832 15564
rect 48780 15521 48789 15555
rect 48789 15521 48823 15555
rect 48823 15521 48832 15555
rect 48780 15512 48832 15521
rect 53932 15580 53984 15632
rect 54300 15580 54352 15632
rect 55772 15580 55824 15632
rect 58072 15580 58124 15632
rect 26424 15376 26476 15428
rect 26884 15376 26936 15428
rect 49608 15512 49660 15564
rect 54484 15555 54536 15564
rect 54484 15521 54493 15555
rect 54493 15521 54527 15555
rect 54527 15521 54536 15555
rect 54484 15512 54536 15521
rect 54760 15555 54812 15564
rect 54760 15521 54769 15555
rect 54769 15521 54803 15555
rect 54803 15521 54812 15555
rect 54760 15512 54812 15521
rect 55128 15512 55180 15564
rect 55404 15512 55456 15564
rect 56508 15512 56560 15564
rect 58532 15555 58584 15564
rect 58532 15521 58541 15555
rect 58541 15521 58575 15555
rect 58575 15521 58584 15555
rect 58532 15512 58584 15521
rect 58808 15648 58860 15700
rect 58992 15648 59044 15700
rect 65432 15648 65484 15700
rect 72240 15648 72292 15700
rect 77300 15648 77352 15700
rect 78220 15648 78272 15700
rect 65616 15580 65668 15632
rect 68468 15580 68520 15632
rect 69664 15623 69716 15632
rect 17132 15351 17184 15360
rect 17132 15317 17141 15351
rect 17141 15317 17175 15351
rect 17175 15317 17184 15351
rect 17132 15308 17184 15317
rect 17224 15308 17276 15360
rect 18144 15308 18196 15360
rect 31484 15308 31536 15360
rect 32036 15308 32088 15360
rect 35348 15308 35400 15360
rect 38016 15308 38068 15360
rect 41788 15308 41840 15360
rect 47952 15308 48004 15360
rect 48044 15308 48096 15360
rect 55864 15444 55916 15496
rect 58808 15444 58860 15496
rect 58992 15487 59044 15496
rect 58992 15453 59001 15487
rect 59001 15453 59035 15487
rect 59035 15453 59044 15487
rect 58992 15444 59044 15453
rect 59176 15444 59228 15496
rect 62396 15444 62448 15496
rect 62948 15512 63000 15564
rect 65432 15512 65484 15564
rect 69388 15512 69440 15564
rect 69664 15589 69673 15623
rect 69673 15589 69707 15623
rect 69707 15589 69716 15623
rect 69664 15580 69716 15589
rect 84752 15648 84804 15700
rect 75920 15512 75972 15564
rect 83924 15555 83976 15564
rect 83924 15521 83933 15555
rect 83933 15521 83967 15555
rect 83967 15521 83976 15555
rect 83924 15512 83976 15521
rect 89260 15487 89312 15496
rect 89260 15453 89269 15487
rect 89269 15453 89303 15487
rect 89303 15453 89312 15487
rect 89260 15444 89312 15453
rect 55772 15376 55824 15428
rect 62672 15376 62724 15428
rect 49424 15351 49476 15360
rect 49424 15317 49433 15351
rect 49433 15317 49467 15351
rect 49467 15317 49476 15351
rect 49424 15308 49476 15317
rect 50160 15308 50212 15360
rect 51080 15308 51132 15360
rect 54024 15351 54076 15360
rect 54024 15317 54033 15351
rect 54033 15317 54067 15351
rect 54067 15317 54076 15351
rect 54024 15308 54076 15317
rect 54300 15351 54352 15360
rect 54300 15317 54309 15351
rect 54309 15317 54343 15351
rect 54343 15317 54352 15351
rect 54300 15308 54352 15317
rect 73620 15376 73672 15428
rect 83740 15419 83792 15428
rect 83740 15385 83749 15419
rect 83749 15385 83783 15419
rect 83783 15385 83792 15419
rect 83740 15376 83792 15385
rect 90180 15555 90232 15564
rect 90180 15521 90189 15555
rect 90189 15521 90223 15555
rect 90223 15521 90232 15555
rect 90180 15512 90232 15521
rect 65064 15308 65116 15360
rect 89812 15308 89864 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 65686 15206 65738 15258
rect 65750 15206 65802 15258
rect 65814 15206 65866 15258
rect 65878 15206 65930 15258
rect 96406 15206 96458 15258
rect 96470 15206 96522 15258
rect 96534 15206 96586 15258
rect 96598 15206 96650 15258
rect 12256 15147 12308 15156
rect 12256 15113 12265 15147
rect 12265 15113 12299 15147
rect 12299 15113 12308 15147
rect 12256 15104 12308 15113
rect 7472 15036 7524 15088
rect 19340 15104 19392 15156
rect 20260 15104 20312 15156
rect 24032 15104 24084 15156
rect 52460 15104 52512 15156
rect 53840 15104 53892 15156
rect 55864 15104 55916 15156
rect 62304 15104 62356 15156
rect 63408 15104 63460 15156
rect 68008 15104 68060 15156
rect 68560 15104 68612 15156
rect 19524 15036 19576 15088
rect 19616 15036 19668 15088
rect 6736 14968 6788 15020
rect 31484 15036 31536 15088
rect 31944 15036 31996 15088
rect 32588 15036 32640 15088
rect 20260 14968 20312 15020
rect 20536 14968 20588 15020
rect 33692 14968 33744 15020
rect 37924 15036 37976 15088
rect 41052 15036 41104 15088
rect 41144 15036 41196 15088
rect 42892 15036 42944 15088
rect 45836 15036 45888 15088
rect 51172 15036 51224 15088
rect 51264 15036 51316 15088
rect 55680 15036 55732 15088
rect 36268 14968 36320 15020
rect 51080 14968 51132 15020
rect 54760 14968 54812 15020
rect 9864 14900 9916 14952
rect 17960 14900 18012 14952
rect 13084 14832 13136 14884
rect 19708 14943 19760 14952
rect 19708 14909 19717 14943
rect 19717 14909 19751 14943
rect 19751 14909 19760 14943
rect 19708 14900 19760 14909
rect 18972 14875 19024 14884
rect 18972 14841 18981 14875
rect 18981 14841 19015 14875
rect 19015 14841 19024 14875
rect 18972 14832 19024 14841
rect 9772 14764 9824 14816
rect 19340 14832 19392 14884
rect 19432 14832 19484 14884
rect 19616 14832 19668 14884
rect 19156 14764 19208 14816
rect 22836 14900 22888 14952
rect 33140 14943 33192 14952
rect 33140 14909 33149 14943
rect 33149 14909 33183 14943
rect 33183 14909 33192 14943
rect 33140 14900 33192 14909
rect 33232 14900 33284 14952
rect 35532 14943 35584 14952
rect 35532 14909 35541 14943
rect 35541 14909 35575 14943
rect 35575 14909 35584 14943
rect 35532 14900 35584 14909
rect 26516 14832 26568 14884
rect 26884 14832 26936 14884
rect 35808 14943 35860 14952
rect 35808 14909 35817 14943
rect 35817 14909 35851 14943
rect 35851 14909 35860 14943
rect 35808 14900 35860 14909
rect 35992 14900 36044 14952
rect 36544 14900 36596 14952
rect 20536 14764 20588 14816
rect 20720 14764 20772 14816
rect 43812 14900 43864 14952
rect 46112 14900 46164 14952
rect 48044 14900 48096 14952
rect 51172 14900 51224 14952
rect 54300 14900 54352 14952
rect 57796 14900 57848 14952
rect 58348 14900 58400 14952
rect 58440 14900 58492 14952
rect 59268 14900 59320 14952
rect 59452 14900 59504 14952
rect 60464 14943 60516 14952
rect 60464 14909 60473 14943
rect 60473 14909 60507 14943
rect 60507 14909 60516 14943
rect 60464 14900 60516 14909
rect 53656 14832 53708 14884
rect 61292 14900 61344 14952
rect 62120 15036 62172 15088
rect 62764 15036 62816 15088
rect 70032 15036 70084 15088
rect 75092 15104 75144 15156
rect 78496 15104 78548 15156
rect 92204 15147 92256 15156
rect 92204 15113 92213 15147
rect 92213 15113 92247 15147
rect 92247 15113 92256 15147
rect 92204 15104 92256 15113
rect 92388 15104 92440 15156
rect 93860 15104 93912 15156
rect 77300 15036 77352 15088
rect 62396 14968 62448 15020
rect 97448 14968 97500 15020
rect 68008 14900 68060 14952
rect 69756 14900 69808 14952
rect 70308 14943 70360 14952
rect 70308 14909 70317 14943
rect 70317 14909 70351 14943
rect 70351 14909 70360 14943
rect 70308 14900 70360 14909
rect 71780 14900 71832 14952
rect 62120 14832 62172 14884
rect 71044 14832 71096 14884
rect 73436 14832 73488 14884
rect 69664 14764 69716 14816
rect 92020 14832 92072 14884
rect 92480 14900 92532 14952
rect 94964 14764 95016 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 50326 14662 50378 14714
rect 50390 14662 50442 14714
rect 50454 14662 50506 14714
rect 50518 14662 50570 14714
rect 81046 14662 81098 14714
rect 81110 14662 81162 14714
rect 81174 14662 81226 14714
rect 81238 14662 81290 14714
rect 17316 14560 17368 14612
rect 24584 14560 24636 14612
rect 31852 14603 31904 14612
rect 17684 14492 17736 14544
rect 26884 14492 26936 14544
rect 5448 14356 5500 14408
rect 8208 14356 8260 14408
rect 18972 14424 19024 14476
rect 20260 14424 20312 14476
rect 30472 14467 30524 14476
rect 30472 14433 30481 14467
rect 30481 14433 30515 14467
rect 30515 14433 30524 14467
rect 30472 14424 30524 14433
rect 31852 14569 31861 14603
rect 31861 14569 31895 14603
rect 31895 14569 31904 14603
rect 31852 14560 31904 14569
rect 34704 14560 34756 14612
rect 35808 14560 35860 14612
rect 37648 14560 37700 14612
rect 41144 14560 41196 14612
rect 55864 14560 55916 14612
rect 56232 14560 56284 14612
rect 60280 14603 60332 14612
rect 38016 14424 38068 14476
rect 6644 14263 6696 14272
rect 6644 14229 6653 14263
rect 6653 14229 6687 14263
rect 6687 14229 6696 14263
rect 6644 14220 6696 14229
rect 11152 14220 11204 14272
rect 23664 14356 23716 14408
rect 43904 14492 43956 14544
rect 46388 14492 46440 14544
rect 51080 14492 51132 14544
rect 40776 14467 40828 14476
rect 40776 14433 40785 14467
rect 40785 14433 40819 14467
rect 40819 14433 40828 14467
rect 40776 14424 40828 14433
rect 43168 14424 43220 14476
rect 52552 14492 52604 14544
rect 53288 14492 53340 14544
rect 51264 14424 51316 14476
rect 54760 14424 54812 14476
rect 54944 14424 54996 14476
rect 57244 14492 57296 14544
rect 57796 14492 57848 14544
rect 60280 14569 60289 14603
rect 60289 14569 60323 14603
rect 60323 14569 60332 14603
rect 60280 14560 60332 14569
rect 63408 14560 63460 14612
rect 81900 14560 81952 14612
rect 13084 14263 13136 14272
rect 13084 14229 13093 14263
rect 13093 14229 13127 14263
rect 13127 14229 13136 14263
rect 13084 14220 13136 14229
rect 43536 14356 43588 14408
rect 49056 14356 49108 14408
rect 55128 14356 55180 14408
rect 55496 14424 55548 14476
rect 58716 14424 58768 14476
rect 59636 14467 59688 14476
rect 59636 14433 59645 14467
rect 59645 14433 59679 14467
rect 59679 14433 59688 14467
rect 59636 14424 59688 14433
rect 59728 14424 59780 14476
rect 60188 14467 60240 14476
rect 60188 14433 60197 14467
rect 60197 14433 60231 14467
rect 60231 14433 60240 14467
rect 60188 14424 60240 14433
rect 60740 14424 60792 14476
rect 63500 14424 63552 14476
rect 63684 14424 63736 14476
rect 35256 14288 35308 14340
rect 43076 14220 43128 14272
rect 43720 14220 43772 14272
rect 43904 14220 43956 14272
rect 51264 14220 51316 14272
rect 52460 14288 52512 14340
rect 55588 14288 55640 14340
rect 60280 14288 60332 14340
rect 60464 14288 60516 14340
rect 67456 14356 67508 14408
rect 69848 14424 69900 14476
rect 70400 14535 70452 14544
rect 70400 14501 70409 14535
rect 70409 14501 70443 14535
rect 70443 14501 70452 14535
rect 70400 14492 70452 14501
rect 70768 14424 70820 14476
rect 75368 14492 75420 14544
rect 91928 14492 91980 14544
rect 61108 14288 61160 14340
rect 75368 14356 75420 14408
rect 96252 14356 96304 14408
rect 96712 14399 96764 14408
rect 96712 14365 96721 14399
rect 96721 14365 96755 14399
rect 96755 14365 96764 14399
rect 96712 14356 96764 14365
rect 97172 14467 97224 14476
rect 97172 14433 97181 14467
rect 97181 14433 97215 14467
rect 97215 14433 97224 14467
rect 97172 14424 97224 14433
rect 81716 14288 81768 14340
rect 60740 14220 60792 14272
rect 60832 14220 60884 14272
rect 70584 14220 70636 14272
rect 70676 14220 70728 14272
rect 72700 14220 72752 14272
rect 81900 14220 81952 14272
rect 89812 14220 89864 14272
rect 97264 14220 97316 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 65686 14118 65738 14170
rect 65750 14118 65802 14170
rect 65814 14118 65866 14170
rect 65878 14118 65930 14170
rect 96406 14118 96458 14170
rect 96470 14118 96522 14170
rect 96534 14118 96586 14170
rect 96598 14118 96650 14170
rect 13084 14016 13136 14068
rect 31208 14016 31260 14068
rect 33968 14016 34020 14068
rect 40408 14016 40460 14068
rect 40868 14059 40920 14068
rect 40868 14025 40877 14059
rect 40877 14025 40911 14059
rect 40911 14025 40920 14059
rect 40868 14016 40920 14025
rect 66904 14016 66956 14068
rect 70584 14016 70636 14068
rect 72700 14016 72752 14068
rect 76196 14016 76248 14068
rect 86224 14016 86276 14068
rect 6644 13948 6696 14000
rect 13544 13948 13596 14000
rect 32496 13948 32548 14000
rect 41144 13948 41196 14000
rect 10324 13923 10376 13932
rect 10324 13889 10333 13923
rect 10333 13889 10367 13923
rect 10367 13889 10376 13923
rect 10324 13880 10376 13889
rect 10600 13880 10652 13932
rect 24124 13880 24176 13932
rect 40408 13880 40460 13932
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 9772 13812 9824 13821
rect 9864 13812 9916 13864
rect 5080 13744 5132 13796
rect 17224 13744 17276 13796
rect 22100 13744 22152 13796
rect 22744 13744 22796 13796
rect 27344 13744 27396 13796
rect 31392 13744 31444 13796
rect 36912 13744 36964 13796
rect 40408 13744 40460 13796
rect 42984 13812 43036 13864
rect 43812 13880 43864 13932
rect 43720 13855 43772 13864
rect 42524 13744 42576 13796
rect 43720 13821 43729 13855
rect 43729 13821 43763 13855
rect 43763 13821 43772 13855
rect 43720 13812 43772 13821
rect 47032 13948 47084 14000
rect 50804 13948 50856 14000
rect 58716 13948 58768 14000
rect 60832 13948 60884 14000
rect 44088 13880 44140 13932
rect 53104 13880 53156 13932
rect 46020 13812 46072 13864
rect 46388 13812 46440 13864
rect 49516 13855 49568 13864
rect 49516 13821 49525 13855
rect 49525 13821 49559 13855
rect 49559 13821 49568 13855
rect 49516 13812 49568 13821
rect 43628 13744 43680 13796
rect 45192 13744 45244 13796
rect 48320 13744 48372 13796
rect 49332 13744 49384 13796
rect 49608 13744 49660 13796
rect 54852 13744 54904 13796
rect 55680 13812 55732 13864
rect 56048 13812 56100 13864
rect 56876 13880 56928 13932
rect 65984 13923 66036 13932
rect 65984 13889 65993 13923
rect 65993 13889 66027 13923
rect 66027 13889 66036 13923
rect 65984 13880 66036 13889
rect 66260 13880 66312 13932
rect 66536 13812 66588 13864
rect 66904 13880 66956 13932
rect 71872 13880 71924 13932
rect 72056 13880 72108 13932
rect 96252 13948 96304 14000
rect 55772 13744 55824 13796
rect 56508 13744 56560 13796
rect 57980 13744 58032 13796
rect 65524 13744 65576 13796
rect 10232 13676 10284 13728
rect 62120 13676 62172 13728
rect 63684 13676 63736 13728
rect 69020 13812 69072 13864
rect 69756 13744 69808 13796
rect 70032 13812 70084 13864
rect 72700 13855 72752 13864
rect 72700 13821 72709 13855
rect 72709 13821 72743 13855
rect 72743 13821 72752 13855
rect 72700 13812 72752 13821
rect 72884 13855 72936 13864
rect 72884 13821 72893 13855
rect 72893 13821 72927 13855
rect 72927 13821 72936 13855
rect 72884 13812 72936 13821
rect 79876 13880 79928 13932
rect 82728 13812 82780 13864
rect 97448 14016 97500 14068
rect 97264 13923 97316 13932
rect 97264 13889 97273 13923
rect 97273 13889 97307 13923
rect 97307 13889 97316 13923
rect 97264 13880 97316 13889
rect 97356 13855 97408 13864
rect 97356 13821 97365 13855
rect 97365 13821 97399 13855
rect 97399 13821 97408 13855
rect 97356 13812 97408 13821
rect 65984 13676 66036 13728
rect 81348 13676 81400 13728
rect 88524 13676 88576 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 50326 13574 50378 13626
rect 50390 13574 50442 13626
rect 50454 13574 50506 13626
rect 50518 13574 50570 13626
rect 81046 13574 81098 13626
rect 81110 13574 81162 13626
rect 81174 13574 81226 13626
rect 81238 13574 81290 13626
rect 13268 13472 13320 13524
rect 13544 13472 13596 13524
rect 45192 13472 45244 13524
rect 48228 13472 48280 13524
rect 49792 13472 49844 13524
rect 96712 13472 96764 13524
rect 3608 13404 3660 13456
rect 20444 13404 20496 13456
rect 22468 13404 22520 13456
rect 26792 13336 26844 13388
rect 27068 13379 27120 13388
rect 27068 13345 27077 13379
rect 27077 13345 27111 13379
rect 27111 13345 27120 13379
rect 27068 13336 27120 13345
rect 27252 13379 27304 13388
rect 27252 13345 27261 13379
rect 27261 13345 27295 13379
rect 27295 13345 27304 13379
rect 27252 13336 27304 13345
rect 27712 13404 27764 13456
rect 39028 13404 39080 13456
rect 33784 13336 33836 13388
rect 36728 13336 36780 13388
rect 39396 13336 39448 13388
rect 39764 13336 39816 13388
rect 45928 13404 45980 13456
rect 62580 13404 62632 13456
rect 65984 13404 66036 13456
rect 66168 13404 66220 13456
rect 12992 13268 13044 13320
rect 16948 13268 17000 13320
rect 42800 13268 42852 13320
rect 64972 13268 65024 13320
rect 65524 13336 65576 13388
rect 71780 13336 71832 13388
rect 72792 13379 72844 13388
rect 72792 13345 72801 13379
rect 72801 13345 72835 13379
rect 72835 13345 72844 13379
rect 72792 13336 72844 13345
rect 72976 13336 73028 13388
rect 75368 13404 75420 13456
rect 85672 13404 85724 13456
rect 69112 13268 69164 13320
rect 70124 13268 70176 13320
rect 75736 13268 75788 13320
rect 83096 13336 83148 13388
rect 83372 13268 83424 13320
rect 13084 13200 13136 13252
rect 44640 13200 44692 13252
rect 49240 13200 49292 13252
rect 49792 13200 49844 13252
rect 54300 13200 54352 13252
rect 81348 13200 81400 13252
rect 12900 13132 12952 13184
rect 16028 13132 16080 13184
rect 20536 13132 20588 13184
rect 28632 13132 28684 13184
rect 36728 13132 36780 13184
rect 37004 13132 37056 13184
rect 46388 13132 46440 13184
rect 82084 13132 82136 13184
rect 93952 13132 94004 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 65686 13030 65738 13082
rect 65750 13030 65802 13082
rect 65814 13030 65866 13082
rect 65878 13030 65930 13082
rect 96406 13030 96458 13082
rect 96470 13030 96522 13082
rect 96534 13030 96586 13082
rect 96598 13030 96650 13082
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 22100 12928 22152 12980
rect 22376 12971 22428 12980
rect 22376 12937 22385 12971
rect 22385 12937 22419 12971
rect 22419 12937 22428 12971
rect 22376 12928 22428 12937
rect 23020 12928 23072 12980
rect 30380 12928 30432 12980
rect 40408 12928 40460 12980
rect 17224 12860 17276 12912
rect 28632 12860 28684 12912
rect 31392 12860 31444 12912
rect 52828 12928 52880 12980
rect 54852 12928 54904 12980
rect 55128 12928 55180 12980
rect 75368 12928 75420 12980
rect 75460 12928 75512 12980
rect 60464 12860 60516 12912
rect 65064 12860 65116 12912
rect 65248 12860 65300 12912
rect 66444 12860 66496 12912
rect 67180 12860 67232 12912
rect 69756 12860 69808 12912
rect 79692 12928 79744 12980
rect 7656 12767 7708 12776
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 8208 12724 8260 12776
rect 12716 12724 12768 12776
rect 12992 12724 13044 12776
rect 17408 12792 17460 12844
rect 39120 12792 39172 12844
rect 39672 12792 39724 12844
rect 43168 12792 43220 12844
rect 43812 12835 43864 12844
rect 43812 12801 43821 12835
rect 43821 12801 43855 12835
rect 43855 12801 43864 12835
rect 43812 12792 43864 12801
rect 46388 12792 46440 12844
rect 63684 12792 63736 12844
rect 85580 12860 85632 12912
rect 13084 12656 13136 12708
rect 22560 12724 22612 12776
rect 23020 12767 23072 12776
rect 23020 12733 23029 12767
rect 23029 12733 23063 12767
rect 23063 12733 23072 12767
rect 23020 12724 23072 12733
rect 39580 12724 39632 12776
rect 39764 12724 39816 12776
rect 31024 12656 31076 12708
rect 40316 12656 40368 12708
rect 42432 12724 42484 12776
rect 43536 12767 43588 12776
rect 43536 12733 43545 12767
rect 43545 12733 43579 12767
rect 43579 12733 43588 12767
rect 43536 12724 43588 12733
rect 13820 12588 13872 12640
rect 16856 12588 16908 12640
rect 17224 12588 17276 12640
rect 21548 12588 21600 12640
rect 24216 12588 24268 12640
rect 39120 12588 39172 12640
rect 42248 12588 42300 12640
rect 44640 12588 44692 12640
rect 48228 12724 48280 12776
rect 46572 12656 46624 12708
rect 54300 12656 54352 12708
rect 55772 12724 55824 12776
rect 58624 12656 58676 12708
rect 60556 12656 60608 12708
rect 61752 12656 61804 12708
rect 61844 12656 61896 12708
rect 65432 12656 65484 12708
rect 66168 12724 66220 12776
rect 66444 12767 66496 12776
rect 66444 12733 66453 12767
rect 66453 12733 66487 12767
rect 66487 12733 66496 12767
rect 66444 12724 66496 12733
rect 65984 12656 66036 12708
rect 69848 12656 69900 12708
rect 70216 12588 70268 12640
rect 71596 12767 71648 12776
rect 71596 12733 71605 12767
rect 71605 12733 71639 12767
rect 71639 12733 71648 12767
rect 71596 12724 71648 12733
rect 71688 12724 71740 12776
rect 72424 12724 72476 12776
rect 75460 12724 75512 12776
rect 81900 12724 81952 12776
rect 85580 12724 85632 12776
rect 85856 12767 85908 12776
rect 85856 12733 85865 12767
rect 85865 12733 85899 12767
rect 85899 12733 85908 12767
rect 85856 12724 85908 12733
rect 86040 12767 86092 12776
rect 86040 12733 86049 12767
rect 86049 12733 86083 12767
rect 86083 12733 86092 12767
rect 86040 12724 86092 12733
rect 75736 12656 75788 12708
rect 75460 12631 75512 12640
rect 75460 12597 75469 12631
rect 75469 12597 75503 12631
rect 75503 12597 75512 12631
rect 75460 12588 75512 12597
rect 75920 12588 75972 12640
rect 85396 12631 85448 12640
rect 85396 12597 85405 12631
rect 85405 12597 85439 12631
rect 85439 12597 85448 12631
rect 85396 12588 85448 12597
rect 85672 12588 85724 12640
rect 85856 12588 85908 12640
rect 90640 12588 90692 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 50326 12486 50378 12538
rect 50390 12486 50442 12538
rect 50454 12486 50506 12538
rect 50518 12486 50570 12538
rect 81046 12486 81098 12538
rect 81110 12486 81162 12538
rect 81174 12486 81226 12538
rect 81238 12486 81290 12538
rect 7012 12384 7064 12436
rect 38200 12384 38252 12436
rect 38568 12384 38620 12436
rect 10784 12316 10836 12368
rect 20444 12316 20496 12368
rect 10876 12291 10928 12300
rect 10876 12257 10885 12291
rect 10885 12257 10919 12291
rect 10919 12257 10928 12291
rect 10876 12248 10928 12257
rect 17960 12248 18012 12300
rect 35348 12316 35400 12368
rect 37924 12316 37976 12368
rect 38016 12316 38068 12368
rect 42708 12359 42760 12368
rect 42708 12325 42717 12359
rect 42717 12325 42751 12359
rect 42751 12325 42760 12359
rect 42708 12316 42760 12325
rect 42800 12359 42852 12368
rect 42800 12325 42809 12359
rect 42809 12325 42843 12359
rect 42843 12325 42852 12359
rect 42800 12316 42852 12325
rect 47216 12316 47268 12368
rect 54668 12316 54720 12368
rect 30748 12248 30800 12300
rect 35900 12248 35952 12300
rect 36452 12248 36504 12300
rect 42064 12248 42116 12300
rect 42248 12248 42300 12300
rect 42524 12291 42576 12300
rect 42524 12257 42533 12291
rect 42533 12257 42567 12291
rect 42567 12257 42576 12291
rect 42524 12248 42576 12257
rect 42892 12291 42944 12300
rect 42892 12257 42901 12291
rect 42901 12257 42935 12291
rect 42935 12257 42944 12291
rect 42892 12248 42944 12257
rect 44640 12248 44692 12300
rect 44824 12248 44876 12300
rect 45652 12248 45704 12300
rect 47124 12248 47176 12300
rect 56048 12384 56100 12436
rect 57428 12316 57480 12368
rect 59544 12384 59596 12436
rect 65432 12384 65484 12436
rect 65892 12384 65944 12436
rect 91008 12384 91060 12436
rect 26424 12180 26476 12232
rect 30472 12180 30524 12232
rect 32036 12180 32088 12232
rect 37556 12180 37608 12232
rect 42432 12180 42484 12232
rect 46204 12223 46256 12232
rect 46204 12189 46213 12223
rect 46213 12189 46247 12223
rect 46247 12189 46256 12223
rect 46204 12180 46256 12189
rect 46664 12180 46716 12232
rect 48044 12180 48096 12232
rect 50068 12180 50120 12232
rect 58808 12291 58860 12300
rect 58808 12257 58817 12291
rect 58817 12257 58851 12291
rect 58851 12257 58860 12291
rect 58808 12248 58860 12257
rect 70768 12316 70820 12368
rect 55864 12180 55916 12232
rect 55956 12180 56008 12232
rect 58072 12180 58124 12232
rect 58532 12180 58584 12232
rect 58992 12180 59044 12232
rect 3424 12112 3476 12164
rect 30656 12112 30708 12164
rect 36544 12112 36596 12164
rect 41696 12112 41748 12164
rect 42708 12112 42760 12164
rect 46020 12112 46072 12164
rect 47308 12112 47360 12164
rect 59268 12248 59320 12300
rect 64972 12248 65024 12300
rect 62672 12180 62724 12232
rect 63960 12180 64012 12232
rect 65892 12248 65944 12300
rect 75460 12316 75512 12368
rect 85396 12316 85448 12368
rect 85672 12316 85724 12368
rect 72608 12291 72660 12300
rect 72608 12257 72617 12291
rect 72617 12257 72651 12291
rect 72651 12257 72660 12291
rect 72608 12248 72660 12257
rect 65524 12180 65576 12232
rect 93676 12180 93728 12232
rect 59268 12112 59320 12164
rect 31024 12044 31076 12096
rect 32496 12044 32548 12096
rect 39580 12044 39632 12096
rect 40500 12044 40552 12096
rect 42984 12044 43036 12096
rect 45468 12044 45520 12096
rect 45652 12044 45704 12096
rect 46664 12044 46716 12096
rect 46848 12044 46900 12096
rect 49056 12044 49108 12096
rect 50068 12044 50120 12096
rect 50712 12044 50764 12096
rect 54668 12044 54720 12096
rect 56508 12044 56560 12096
rect 57704 12087 57756 12096
rect 57704 12053 57713 12087
rect 57713 12053 57747 12087
rect 57747 12053 57756 12087
rect 57704 12044 57756 12053
rect 61568 12044 61620 12096
rect 65340 12087 65392 12096
rect 65340 12053 65349 12087
rect 65349 12053 65383 12087
rect 65383 12053 65392 12087
rect 65340 12044 65392 12053
rect 67364 12087 67416 12096
rect 67364 12053 67373 12087
rect 67373 12053 67407 12087
rect 67407 12053 67416 12087
rect 67364 12044 67416 12053
rect 97540 12044 97592 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 65686 11942 65738 11994
rect 65750 11942 65802 11994
rect 65814 11942 65866 11994
rect 65878 11942 65930 11994
rect 96406 11942 96458 11994
rect 96470 11942 96522 11994
rect 96534 11942 96586 11994
rect 96598 11942 96650 11994
rect 2228 11840 2280 11892
rect 38660 11840 38712 11892
rect 10324 11815 10376 11824
rect 10324 11781 10333 11815
rect 10333 11781 10367 11815
rect 10367 11781 10376 11815
rect 10324 11772 10376 11781
rect 17132 11772 17184 11824
rect 17960 11772 18012 11824
rect 6920 11636 6972 11688
rect 9312 11568 9364 11620
rect 18420 11704 18472 11756
rect 26332 11772 26384 11824
rect 27160 11772 27212 11824
rect 28080 11704 28132 11756
rect 28632 11747 28684 11756
rect 28632 11713 28641 11747
rect 28641 11713 28675 11747
rect 28675 11713 28684 11747
rect 28632 11704 28684 11713
rect 36360 11704 36412 11756
rect 42064 11840 42116 11892
rect 42248 11840 42300 11892
rect 46848 11840 46900 11892
rect 47768 11840 47820 11892
rect 57980 11840 58032 11892
rect 58072 11840 58124 11892
rect 59268 11840 59320 11892
rect 62672 11840 62724 11892
rect 70124 11840 70176 11892
rect 70308 11840 70360 11892
rect 79692 11840 79744 11892
rect 38844 11772 38896 11824
rect 12532 11568 12584 11620
rect 12900 11568 12952 11620
rect 7564 11500 7616 11552
rect 17316 11568 17368 11620
rect 27528 11636 27580 11688
rect 25228 11568 25280 11620
rect 37924 11636 37976 11688
rect 15016 11543 15068 11552
rect 15016 11509 15025 11543
rect 15025 11509 15059 11543
rect 15059 11509 15068 11543
rect 15016 11500 15068 11509
rect 25504 11500 25556 11552
rect 28356 11500 28408 11552
rect 30380 11500 30432 11552
rect 32036 11500 32088 11552
rect 37556 11500 37608 11552
rect 37648 11500 37700 11552
rect 38016 11500 38068 11552
rect 38381 11679 38433 11688
rect 38381 11645 38393 11679
rect 38393 11645 38427 11679
rect 38427 11645 38433 11679
rect 38568 11679 38620 11688
rect 38381 11636 38433 11645
rect 38568 11645 38576 11679
rect 38576 11645 38610 11679
rect 38610 11645 38620 11679
rect 38568 11636 38620 11645
rect 38660 11679 38712 11688
rect 38660 11645 38669 11679
rect 38669 11645 38703 11679
rect 38703 11645 38712 11679
rect 39028 11704 39080 11756
rect 39396 11772 39448 11824
rect 45652 11772 45704 11824
rect 46204 11772 46256 11824
rect 56600 11772 56652 11824
rect 58992 11772 59044 11824
rect 65524 11772 65576 11824
rect 39764 11704 39816 11756
rect 41972 11704 42024 11756
rect 42064 11704 42116 11756
rect 69480 11704 69532 11756
rect 75552 11747 75604 11756
rect 38660 11636 38712 11645
rect 38752 11500 38804 11552
rect 62672 11636 62724 11688
rect 75552 11713 75561 11747
rect 75561 11713 75595 11747
rect 75595 11713 75604 11747
rect 75552 11704 75604 11713
rect 39580 11568 39632 11620
rect 67272 11568 67324 11620
rect 69480 11568 69532 11620
rect 85488 11815 85540 11824
rect 85488 11781 85497 11815
rect 85497 11781 85531 11815
rect 85531 11781 85540 11815
rect 85488 11772 85540 11781
rect 91008 11815 91060 11824
rect 91008 11781 91017 11815
rect 91017 11781 91051 11815
rect 91051 11781 91060 11815
rect 91008 11772 91060 11781
rect 67640 11500 67692 11552
rect 75460 11500 75512 11552
rect 92572 11500 92624 11552
rect 96712 11500 96764 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 50326 11398 50378 11450
rect 50390 11398 50442 11450
rect 50454 11398 50506 11450
rect 50518 11398 50570 11450
rect 81046 11398 81098 11450
rect 81110 11398 81162 11450
rect 81174 11398 81226 11450
rect 81238 11398 81290 11450
rect 12532 11296 12584 11348
rect 36544 11296 36596 11348
rect 38200 11296 38252 11348
rect 12348 11203 12400 11212
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 12348 11169 12357 11203
rect 12357 11169 12391 11203
rect 12391 11169 12400 11203
rect 12348 11160 12400 11169
rect 12532 11160 12584 11212
rect 12900 11203 12952 11212
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 13084 11160 13136 11212
rect 26792 11228 26844 11280
rect 28356 11271 28408 11280
rect 28356 11237 28365 11271
rect 28365 11237 28399 11271
rect 28399 11237 28408 11271
rect 28356 11228 28408 11237
rect 21732 11203 21784 11212
rect 21732 11169 21741 11203
rect 21741 11169 21775 11203
rect 21775 11169 21784 11203
rect 21732 11160 21784 11169
rect 26332 11160 26384 11212
rect 6920 11092 6972 11144
rect 7656 11092 7708 11144
rect 12808 11135 12860 11144
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 12808 11092 12860 11101
rect 26424 11092 26476 11144
rect 26884 11092 26936 11144
rect 27252 11160 27304 11212
rect 36452 11160 36504 11212
rect 37280 11160 37332 11212
rect 38384 11296 38436 11348
rect 38568 11296 38620 11348
rect 41972 11296 42024 11348
rect 55864 11296 55916 11348
rect 60372 11296 60424 11348
rect 38568 11203 38620 11212
rect 38568 11169 38577 11203
rect 38577 11169 38611 11203
rect 38611 11169 38620 11203
rect 38844 11228 38896 11280
rect 38568 11160 38620 11169
rect 4896 10956 4948 11008
rect 41604 11160 41656 11212
rect 42984 11228 43036 11280
rect 67456 11296 67508 11348
rect 69296 11296 69348 11348
rect 55496 11092 55548 11144
rect 55864 11160 55916 11212
rect 62948 11160 63000 11212
rect 67824 11228 67876 11280
rect 69848 11296 69900 11348
rect 97540 11339 97592 11348
rect 97540 11305 97549 11339
rect 97549 11305 97583 11339
rect 97583 11305 97592 11339
rect 97540 11296 97592 11305
rect 58072 11092 58124 11144
rect 59728 11092 59780 11144
rect 72332 11160 72384 11212
rect 73896 11160 73948 11212
rect 79784 11160 79836 11212
rect 82636 11160 82688 11212
rect 96712 11203 96764 11212
rect 96712 11169 96721 11203
rect 96721 11169 96755 11203
rect 96755 11169 96764 11203
rect 96712 11160 96764 11169
rect 86500 11024 86552 11076
rect 92664 11024 92716 11076
rect 12440 10956 12492 11008
rect 12532 10999 12584 11008
rect 12532 10965 12541 10999
rect 12541 10965 12575 10999
rect 12575 10965 12584 10999
rect 25228 10999 25280 11008
rect 12532 10956 12584 10965
rect 25228 10965 25237 10999
rect 25237 10965 25271 10999
rect 25271 10965 25280 10999
rect 25228 10956 25280 10965
rect 26240 10956 26292 11008
rect 28632 10956 28684 11008
rect 35808 10956 35860 11008
rect 61476 10956 61528 11008
rect 61568 10956 61620 11008
rect 62856 10956 62908 11008
rect 64328 10956 64380 11008
rect 83096 10956 83148 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 65686 10854 65738 10906
rect 65750 10854 65802 10906
rect 65814 10854 65866 10906
rect 65878 10854 65930 10906
rect 96406 10854 96458 10906
rect 96470 10854 96522 10906
rect 96534 10854 96586 10906
rect 96598 10854 96650 10906
rect 12440 10752 12492 10804
rect 28448 10752 28500 10804
rect 28632 10752 28684 10804
rect 42892 10752 42944 10804
rect 44640 10752 44692 10804
rect 45100 10752 45152 10804
rect 46388 10752 46440 10804
rect 57980 10752 58032 10804
rect 91560 10752 91612 10804
rect 12256 10684 12308 10736
rect 32772 10684 32824 10736
rect 25964 10616 26016 10668
rect 36544 10684 36596 10736
rect 44364 10684 44416 10736
rect 45376 10684 45428 10736
rect 49424 10684 49476 10736
rect 51724 10684 51776 10736
rect 61660 10684 61712 10736
rect 67272 10727 67324 10736
rect 67272 10693 67281 10727
rect 67281 10693 67315 10727
rect 67315 10693 67324 10727
rect 67272 10684 67324 10693
rect 41144 10616 41196 10668
rect 20076 10548 20128 10600
rect 27252 10548 27304 10600
rect 33232 10548 33284 10600
rect 33416 10548 33468 10600
rect 36452 10548 36504 10600
rect 5448 10480 5500 10532
rect 41788 10548 41840 10600
rect 44180 10591 44232 10600
rect 44180 10557 44189 10591
rect 44189 10557 44223 10591
rect 44223 10557 44232 10591
rect 44180 10548 44232 10557
rect 44272 10548 44324 10600
rect 46296 10616 46348 10668
rect 46572 10616 46624 10668
rect 61476 10616 61528 10668
rect 45192 10548 45244 10600
rect 47768 10548 47820 10600
rect 51724 10548 51776 10600
rect 51908 10548 51960 10600
rect 58164 10548 58216 10600
rect 37924 10480 37976 10532
rect 39672 10480 39724 10532
rect 12532 10412 12584 10464
rect 41696 10412 41748 10464
rect 50620 10412 50672 10464
rect 57336 10480 57388 10532
rect 61660 10548 61712 10600
rect 61844 10591 61896 10600
rect 61844 10557 61853 10591
rect 61853 10557 61887 10591
rect 61887 10557 61896 10591
rect 61844 10548 61896 10557
rect 64972 10548 65024 10600
rect 69112 10684 69164 10736
rect 87788 10684 87840 10736
rect 65248 10523 65300 10532
rect 62120 10412 62172 10464
rect 62948 10412 63000 10464
rect 63224 10455 63276 10464
rect 63224 10421 63233 10455
rect 63233 10421 63267 10455
rect 63267 10421 63276 10455
rect 63224 10412 63276 10421
rect 65248 10489 65257 10523
rect 65257 10489 65291 10523
rect 65291 10489 65300 10523
rect 65248 10480 65300 10489
rect 68652 10548 68704 10600
rect 85948 10616 86000 10668
rect 75092 10548 75144 10600
rect 71504 10480 71556 10532
rect 77944 10548 77996 10600
rect 82636 10548 82688 10600
rect 75276 10480 75328 10532
rect 68284 10412 68336 10464
rect 75184 10412 75236 10464
rect 96068 10412 96120 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 50326 10310 50378 10362
rect 50390 10310 50442 10362
rect 50454 10310 50506 10362
rect 50518 10310 50570 10362
rect 81046 10310 81098 10362
rect 81110 10310 81162 10362
rect 81174 10310 81226 10362
rect 81238 10310 81290 10362
rect 4896 10183 4948 10192
rect 4896 10149 4905 10183
rect 4905 10149 4939 10183
rect 4939 10149 4948 10183
rect 4896 10140 4948 10149
rect 9772 10208 9824 10260
rect 10876 10208 10928 10260
rect 25780 10208 25832 10260
rect 26240 10208 26292 10260
rect 26332 10208 26384 10260
rect 27252 10251 27304 10260
rect 27252 10217 27261 10251
rect 27261 10217 27295 10251
rect 27295 10217 27304 10251
rect 27252 10208 27304 10217
rect 28080 10251 28132 10260
rect 28080 10217 28089 10251
rect 28089 10217 28123 10251
rect 28123 10217 28132 10251
rect 28080 10208 28132 10217
rect 32772 10208 32824 10260
rect 46204 10208 46256 10260
rect 46480 10208 46532 10260
rect 50712 10208 50764 10260
rect 65248 10208 65300 10260
rect 67364 10208 67416 10260
rect 75184 10208 75236 10260
rect 18512 10072 18564 10124
rect 18788 10072 18840 10124
rect 20076 10072 20128 10124
rect 20812 10072 20864 10124
rect 21180 10072 21232 10124
rect 23388 10072 23440 10124
rect 27068 10072 27120 10124
rect 27988 10115 28040 10124
rect 27988 10081 27997 10115
rect 27997 10081 28031 10115
rect 28031 10081 28040 10115
rect 27988 10072 28040 10081
rect 36544 10140 36596 10192
rect 39212 10140 39264 10192
rect 42432 10140 42484 10192
rect 42800 10140 42852 10192
rect 45376 10140 45428 10192
rect 46296 10140 46348 10192
rect 86776 10140 86828 10192
rect 9128 10004 9180 10056
rect 10508 10004 10560 10056
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 15016 10004 15068 10056
rect 18604 10004 18656 10056
rect 6184 9936 6236 9988
rect 7656 9936 7708 9988
rect 18696 9936 18748 9988
rect 20628 9936 20680 9988
rect 24860 10004 24912 10056
rect 25136 10004 25188 10056
rect 25872 10047 25924 10056
rect 25872 10013 25881 10047
rect 25881 10013 25915 10047
rect 25915 10013 25924 10047
rect 25872 10004 25924 10013
rect 26976 10004 27028 10056
rect 28448 10004 28500 10056
rect 33416 10004 33468 10056
rect 33968 10072 34020 10124
rect 62672 10072 62724 10124
rect 63408 10072 63460 10124
rect 63500 10072 63552 10124
rect 37924 10004 37976 10056
rect 9680 9868 9732 9920
rect 25780 9868 25832 9920
rect 30380 9936 30432 9988
rect 31208 9936 31260 9988
rect 27068 9868 27120 9920
rect 33968 9868 34020 9920
rect 37556 9936 37608 9988
rect 52736 10004 52788 10056
rect 57796 10004 57848 10056
rect 58164 10004 58216 10056
rect 71504 10004 71556 10056
rect 75092 10072 75144 10124
rect 81716 10115 81768 10124
rect 81716 10081 81725 10115
rect 81725 10081 81759 10115
rect 81759 10081 81768 10115
rect 81716 10072 81768 10081
rect 43996 9936 44048 9988
rect 44088 9936 44140 9988
rect 53564 9936 53616 9988
rect 66536 9936 66588 9988
rect 75276 9936 75328 9988
rect 39672 9911 39724 9920
rect 39672 9877 39681 9911
rect 39681 9877 39715 9911
rect 39715 9877 39724 9911
rect 39672 9868 39724 9877
rect 39856 9868 39908 9920
rect 42800 9868 42852 9920
rect 42892 9868 42944 9920
rect 50988 9868 51040 9920
rect 55128 9868 55180 9920
rect 96896 9936 96948 9988
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 65686 9766 65738 9818
rect 65750 9766 65802 9818
rect 65814 9766 65866 9818
rect 65878 9766 65930 9818
rect 96406 9766 96458 9818
rect 96470 9766 96522 9818
rect 96534 9766 96586 9818
rect 96598 9766 96650 9818
rect 12624 9596 12676 9648
rect 14740 9596 14792 9648
rect 18512 9596 18564 9648
rect 20352 9639 20404 9648
rect 20352 9605 20361 9639
rect 20361 9605 20395 9639
rect 20395 9605 20404 9639
rect 20352 9596 20404 9605
rect 20628 9664 20680 9716
rect 62672 9664 62724 9716
rect 63408 9664 63460 9716
rect 68284 9664 68336 9716
rect 68376 9664 68428 9716
rect 73068 9664 73120 9716
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 3608 9503 3660 9512
rect 3608 9469 3617 9503
rect 3617 9469 3651 9503
rect 3651 9469 3660 9503
rect 3608 9460 3660 9469
rect 3700 9435 3752 9444
rect 3700 9401 3709 9435
rect 3709 9401 3743 9435
rect 3743 9401 3752 9435
rect 3700 9392 3752 9401
rect 5264 9392 5316 9444
rect 13636 9528 13688 9580
rect 19248 9528 19300 9580
rect 31576 9528 31628 9580
rect 35808 9528 35860 9580
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 15108 9460 15160 9512
rect 18788 9460 18840 9512
rect 19524 9503 19576 9512
rect 19524 9469 19533 9503
rect 19533 9469 19567 9503
rect 19567 9469 19576 9503
rect 19524 9460 19576 9469
rect 26884 9460 26936 9512
rect 35992 9503 36044 9512
rect 35992 9469 36001 9503
rect 36001 9469 36035 9503
rect 36035 9469 36044 9503
rect 35992 9460 36044 9469
rect 36268 9503 36320 9512
rect 36268 9469 36277 9503
rect 36277 9469 36311 9503
rect 36311 9469 36320 9503
rect 36268 9460 36320 9469
rect 36544 9460 36596 9512
rect 36912 9596 36964 9648
rect 89720 9596 89772 9648
rect 37372 9528 37424 9580
rect 54300 9571 54352 9580
rect 54300 9537 54309 9571
rect 54309 9537 54343 9571
rect 54343 9537 54352 9571
rect 54300 9528 54352 9537
rect 54760 9528 54812 9580
rect 72976 9528 73028 9580
rect 78680 9528 78732 9580
rect 82360 9528 82412 9580
rect 95516 9528 95568 9580
rect 37280 9460 37332 9512
rect 23388 9324 23440 9376
rect 25872 9324 25924 9376
rect 26240 9324 26292 9376
rect 37832 9392 37884 9444
rect 44916 9460 44968 9512
rect 51080 9503 51132 9512
rect 51080 9469 51089 9503
rect 51089 9469 51123 9503
rect 51123 9469 51132 9503
rect 51080 9460 51132 9469
rect 51540 9460 51592 9512
rect 53932 9460 53984 9512
rect 57336 9460 57388 9512
rect 40500 9392 40552 9444
rect 62396 9460 62448 9512
rect 62488 9460 62540 9512
rect 63224 9460 63276 9512
rect 63316 9460 63368 9512
rect 67180 9460 67232 9512
rect 86960 9460 87012 9512
rect 90732 9503 90784 9512
rect 90732 9469 90741 9503
rect 90741 9469 90775 9503
rect 90775 9469 90784 9503
rect 90732 9460 90784 9469
rect 90824 9503 90876 9512
rect 90824 9469 90833 9503
rect 90833 9469 90867 9503
rect 90867 9469 90876 9503
rect 90824 9460 90876 9469
rect 62856 9392 62908 9444
rect 65340 9392 65392 9444
rect 65524 9392 65576 9444
rect 68284 9392 68336 9444
rect 68744 9392 68796 9444
rect 73896 9392 73948 9444
rect 41512 9324 41564 9376
rect 49332 9324 49384 9376
rect 71872 9324 71924 9376
rect 85948 9324 86000 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 50326 9222 50378 9274
rect 50390 9222 50442 9274
rect 50454 9222 50506 9274
rect 50518 9222 50570 9274
rect 81046 9222 81098 9274
rect 81110 9222 81162 9274
rect 81174 9222 81226 9274
rect 81238 9222 81290 9274
rect 10968 9120 11020 9172
rect 12256 9163 12308 9172
rect 5356 9052 5408 9104
rect 9036 9052 9088 9104
rect 4804 8984 4856 9036
rect 5080 9027 5132 9036
rect 5080 8993 5089 9027
rect 5089 8993 5123 9027
rect 5123 8993 5132 9027
rect 5080 8984 5132 8993
rect 7472 8984 7524 9036
rect 11612 9027 11664 9036
rect 11612 8993 11621 9027
rect 11621 8993 11655 9027
rect 11655 8993 11664 9027
rect 11612 8984 11664 8993
rect 11796 9027 11848 9036
rect 11796 8993 11804 9027
rect 11804 8993 11838 9027
rect 11838 8993 11848 9027
rect 11796 8984 11848 8993
rect 12256 9129 12265 9163
rect 12265 9129 12299 9163
rect 12299 9129 12308 9163
rect 12256 9120 12308 9129
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 19340 9120 19392 9172
rect 30380 9120 30432 9172
rect 36912 9120 36964 9172
rect 49884 9120 49936 9172
rect 50804 9120 50856 9172
rect 51080 9120 51132 9172
rect 54484 9120 54536 9172
rect 12164 9027 12216 9036
rect 12164 8993 12173 9027
rect 12173 8993 12207 9027
rect 12207 8993 12216 9027
rect 12164 8984 12216 8993
rect 16396 8984 16448 9036
rect 35716 8984 35768 9036
rect 37004 9052 37056 9104
rect 37280 9052 37332 9104
rect 37372 8984 37424 9036
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 11520 8848 11572 8900
rect 15016 8916 15068 8968
rect 17684 8848 17736 8900
rect 15660 8780 15712 8832
rect 21272 8916 21324 8968
rect 35900 8916 35952 8968
rect 37648 9052 37700 9104
rect 39764 9095 39816 9104
rect 39764 9061 39773 9095
rect 39773 9061 39807 9095
rect 39807 9061 39816 9095
rect 39764 9052 39816 9061
rect 42616 9052 42668 9104
rect 37740 8984 37792 9036
rect 40316 8984 40368 9036
rect 44732 8984 44784 9036
rect 37648 8916 37700 8968
rect 43076 8916 43128 8968
rect 56784 9052 56836 9104
rect 59268 9052 59320 9104
rect 59452 9052 59504 9104
rect 62856 9052 62908 9104
rect 63868 9052 63920 9104
rect 67364 9052 67416 9104
rect 74264 9120 74316 9172
rect 87052 9052 87104 9104
rect 88524 9052 88576 9104
rect 48412 8984 48464 9036
rect 63040 9027 63092 9036
rect 26884 8848 26936 8900
rect 21732 8780 21784 8832
rect 22100 8780 22152 8832
rect 33692 8780 33744 8832
rect 33968 8780 34020 8832
rect 37556 8823 37608 8832
rect 37556 8789 37565 8823
rect 37565 8789 37599 8823
rect 37599 8789 37608 8823
rect 37556 8780 37608 8789
rect 47584 8848 47636 8900
rect 62028 8916 62080 8968
rect 63040 8993 63049 9027
rect 63049 8993 63083 9027
rect 63083 8993 63092 9027
rect 63040 8984 63092 8993
rect 88984 9027 89036 9036
rect 88984 8993 88993 9027
rect 88993 8993 89027 9027
rect 89027 8993 89036 9027
rect 88984 8984 89036 8993
rect 89352 9027 89404 9036
rect 89352 8993 89361 9027
rect 89361 8993 89395 9027
rect 89395 8993 89404 9027
rect 89352 8984 89404 8993
rect 55312 8848 55364 8900
rect 55588 8848 55640 8900
rect 56784 8848 56836 8900
rect 58072 8848 58124 8900
rect 61660 8848 61712 8900
rect 61752 8848 61804 8900
rect 63224 8916 63276 8968
rect 65524 8916 65576 8968
rect 74172 8959 74224 8968
rect 74172 8925 74181 8959
rect 74181 8925 74215 8959
rect 74215 8925 74224 8959
rect 74172 8916 74224 8925
rect 88432 8959 88484 8968
rect 88432 8925 88441 8959
rect 88441 8925 88475 8959
rect 88475 8925 88484 8959
rect 88432 8916 88484 8925
rect 45008 8780 45060 8832
rect 51816 8780 51868 8832
rect 52368 8780 52420 8832
rect 94136 9052 94188 9104
rect 95516 9095 95568 9104
rect 95516 9061 95525 9095
rect 95525 9061 95559 9095
rect 95559 9061 95568 9095
rect 95516 9052 95568 9061
rect 95148 9027 95200 9036
rect 95148 8993 95157 9027
rect 95157 8993 95191 9027
rect 95191 8993 95200 9027
rect 95148 8984 95200 8993
rect 64512 8780 64564 8832
rect 89720 8780 89772 8832
rect 94872 8780 94924 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 65686 8678 65738 8730
rect 65750 8678 65802 8730
rect 65814 8678 65866 8730
rect 65878 8678 65930 8730
rect 96406 8678 96458 8730
rect 96470 8678 96522 8730
rect 96534 8678 96586 8730
rect 96598 8678 96650 8730
rect 20444 8619 20496 8628
rect 20444 8585 20453 8619
rect 20453 8585 20487 8619
rect 20487 8585 20496 8619
rect 20444 8576 20496 8585
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 33416 8576 33468 8628
rect 39396 8576 39448 8628
rect 39948 8576 40000 8628
rect 41328 8576 41380 8628
rect 46480 8576 46532 8628
rect 47676 8576 47728 8628
rect 19892 8440 19944 8492
rect 20260 8440 20312 8492
rect 19340 8372 19392 8424
rect 19984 8415 20036 8424
rect 19984 8381 19992 8415
rect 19992 8381 20026 8415
rect 20026 8381 20036 8415
rect 19984 8372 20036 8381
rect 6644 8304 6696 8356
rect 9220 8304 9272 8356
rect 16212 8304 16264 8356
rect 16488 8304 16540 8356
rect 23020 8415 23072 8424
rect 23020 8381 23029 8415
rect 23029 8381 23063 8415
rect 23063 8381 23072 8415
rect 23020 8372 23072 8381
rect 31852 8440 31904 8492
rect 34336 8483 34388 8492
rect 34336 8449 34345 8483
rect 34345 8449 34379 8483
rect 34379 8449 34388 8483
rect 34336 8440 34388 8449
rect 34612 8440 34664 8492
rect 40408 8508 40460 8560
rect 50804 8508 50856 8560
rect 56600 8576 56652 8628
rect 60740 8576 60792 8628
rect 60832 8576 60884 8628
rect 67364 8576 67416 8628
rect 78956 8576 79008 8628
rect 94136 8619 94188 8628
rect 94136 8585 94145 8619
rect 94145 8585 94179 8619
rect 94179 8585 94188 8619
rect 94136 8576 94188 8585
rect 33416 8372 33468 8424
rect 33692 8415 33744 8424
rect 33692 8381 33701 8415
rect 33701 8381 33735 8415
rect 33735 8381 33744 8415
rect 33692 8372 33744 8381
rect 23388 8347 23440 8356
rect 3700 8236 3752 8288
rect 23388 8313 23397 8347
rect 23397 8313 23431 8347
rect 23431 8313 23440 8347
rect 23388 8304 23440 8313
rect 30288 8304 30340 8356
rect 34428 8304 34480 8356
rect 35716 8415 35768 8424
rect 35716 8381 35725 8415
rect 35725 8381 35759 8415
rect 35759 8381 35768 8415
rect 35716 8372 35768 8381
rect 38752 8372 38804 8424
rect 47492 8440 47544 8492
rect 50528 8440 50580 8492
rect 39028 8372 39080 8424
rect 39396 8372 39448 8424
rect 41512 8372 41564 8424
rect 49240 8415 49292 8424
rect 49240 8381 49249 8415
rect 49249 8381 49283 8415
rect 49283 8381 49292 8415
rect 49240 8372 49292 8381
rect 50436 8372 50488 8424
rect 51080 8440 51132 8492
rect 51540 8508 51592 8560
rect 55588 8508 55640 8560
rect 56508 8508 56560 8560
rect 68100 8508 68152 8560
rect 68284 8508 68336 8560
rect 94872 8508 94924 8560
rect 38660 8304 38712 8356
rect 25964 8236 26016 8288
rect 30932 8236 30984 8288
rect 37556 8236 37608 8288
rect 37648 8236 37700 8288
rect 48504 8304 48556 8356
rect 49332 8304 49384 8356
rect 49976 8304 50028 8356
rect 50804 8304 50856 8356
rect 53840 8372 53892 8424
rect 60832 8372 60884 8424
rect 61660 8372 61712 8424
rect 51172 8304 51224 8356
rect 62212 8372 62264 8424
rect 65524 8372 65576 8424
rect 65984 8415 66036 8424
rect 65984 8381 65993 8415
rect 65993 8381 66027 8415
rect 66027 8381 66036 8415
rect 65984 8372 66036 8381
rect 66168 8372 66220 8424
rect 67456 8415 67508 8424
rect 67456 8381 67465 8415
rect 67465 8381 67499 8415
rect 67499 8381 67508 8415
rect 67456 8372 67508 8381
rect 61844 8347 61896 8356
rect 61844 8313 61853 8347
rect 61853 8313 61887 8347
rect 61887 8313 61896 8347
rect 61844 8304 61896 8313
rect 63868 8304 63920 8356
rect 65248 8304 65300 8356
rect 66076 8304 66128 8356
rect 68100 8304 68152 8356
rect 94136 8304 94188 8356
rect 46204 8236 46256 8288
rect 74080 8236 74132 8288
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 50326 8134 50378 8186
rect 50390 8134 50442 8186
rect 50454 8134 50506 8186
rect 50518 8134 50570 8186
rect 81046 8134 81098 8186
rect 81110 8134 81162 8186
rect 81174 8134 81226 8186
rect 81238 8134 81290 8186
rect 10876 8032 10928 8084
rect 33324 8075 33376 8084
rect 1492 7896 1544 7948
rect 9496 7964 9548 8016
rect 2044 7939 2096 7948
rect 2044 7905 2053 7939
rect 2053 7905 2087 7939
rect 2087 7905 2096 7939
rect 2044 7896 2096 7905
rect 2872 7896 2924 7948
rect 10416 7939 10468 7948
rect 10416 7905 10425 7939
rect 10425 7905 10459 7939
rect 10459 7905 10468 7939
rect 10416 7896 10468 7905
rect 27344 7964 27396 8016
rect 33324 8041 33333 8075
rect 33333 8041 33367 8075
rect 33367 8041 33376 8075
rect 33324 8032 33376 8041
rect 33692 8032 33744 8084
rect 37648 8032 37700 8084
rect 40224 8032 40276 8084
rect 46204 8032 46256 8084
rect 46296 8032 46348 8084
rect 38844 7964 38896 8016
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 10600 7828 10652 7880
rect 25780 7896 25832 7948
rect 31852 7896 31904 7948
rect 32036 7896 32088 7948
rect 32220 7939 32272 7948
rect 32220 7905 32229 7939
rect 32229 7905 32263 7939
rect 32263 7905 32272 7939
rect 32220 7896 32272 7905
rect 37280 7939 37332 7948
rect 37280 7905 37289 7939
rect 37289 7905 37323 7939
rect 37323 7905 37332 7939
rect 37280 7896 37332 7905
rect 38016 7939 38068 7948
rect 32680 7828 32732 7880
rect 33048 7828 33100 7880
rect 37556 7871 37608 7880
rect 37556 7837 37565 7871
rect 37565 7837 37599 7871
rect 37599 7837 37608 7871
rect 37556 7828 37608 7837
rect 38016 7905 38025 7939
rect 38025 7905 38059 7939
rect 38059 7905 38068 7939
rect 38016 7896 38068 7905
rect 40040 7964 40092 8016
rect 39212 7896 39264 7948
rect 38108 7871 38160 7880
rect 38108 7837 38117 7871
rect 38117 7837 38151 7871
rect 38151 7837 38160 7871
rect 38108 7828 38160 7837
rect 38568 7828 38620 7880
rect 38660 7828 38712 7880
rect 39488 7896 39540 7948
rect 46204 7896 46256 7948
rect 49148 8032 49200 8084
rect 87512 8032 87564 8084
rect 47860 7964 47912 8016
rect 90180 7964 90232 8016
rect 81716 7896 81768 7948
rect 81900 7896 81952 7948
rect 83280 7896 83332 7948
rect 46112 7828 46164 7880
rect 46480 7828 46532 7880
rect 67732 7828 67784 7880
rect 73068 7828 73120 7880
rect 91284 7760 91336 7812
rect 10048 7692 10100 7744
rect 45376 7692 45428 7744
rect 45560 7692 45612 7744
rect 46480 7692 46532 7744
rect 46572 7692 46624 7744
rect 49700 7692 49752 7744
rect 50160 7692 50212 7744
rect 50712 7692 50764 7744
rect 54668 7692 54720 7744
rect 56232 7692 56284 7744
rect 56876 7692 56928 7744
rect 63960 7692 64012 7744
rect 66996 7692 67048 7744
rect 67272 7692 67324 7744
rect 77392 7692 77444 7744
rect 77760 7692 77812 7744
rect 77852 7692 77904 7744
rect 83372 7692 83424 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 65686 7590 65738 7642
rect 65750 7590 65802 7642
rect 65814 7590 65866 7642
rect 65878 7590 65930 7642
rect 96406 7590 96458 7642
rect 96470 7590 96522 7642
rect 96534 7590 96586 7642
rect 96598 7590 96650 7642
rect 1860 7488 1912 7540
rect 20904 7488 20956 7540
rect 23388 7488 23440 7540
rect 26792 7488 26844 7540
rect 31024 7488 31076 7540
rect 11888 7463 11940 7472
rect 11888 7429 11897 7463
rect 11897 7429 11931 7463
rect 11931 7429 11940 7463
rect 11888 7420 11940 7429
rect 16948 7420 17000 7472
rect 17776 7420 17828 7472
rect 25780 7420 25832 7472
rect 32588 7420 32640 7472
rect 2872 7352 2924 7404
rect 1492 7284 1544 7336
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 19340 7352 19392 7404
rect 22928 7352 22980 7404
rect 34704 7420 34756 7472
rect 37280 7420 37332 7472
rect 45284 7420 45336 7472
rect 45468 7420 45520 7472
rect 49608 7420 49660 7472
rect 49700 7420 49752 7472
rect 54024 7488 54076 7540
rect 54392 7488 54444 7540
rect 60188 7488 60240 7540
rect 65340 7488 65392 7540
rect 69572 7531 69624 7540
rect 69572 7497 69581 7531
rect 69581 7497 69615 7531
rect 69615 7497 69624 7531
rect 69572 7488 69624 7497
rect 9496 7327 9548 7336
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 9496 7284 9548 7293
rect 10048 7327 10100 7336
rect 10048 7293 10057 7327
rect 10057 7293 10091 7327
rect 10091 7293 10100 7327
rect 10048 7284 10100 7293
rect 20628 7284 20680 7336
rect 24860 7284 24912 7336
rect 25320 7284 25372 7336
rect 24124 7216 24176 7268
rect 34244 7352 34296 7404
rect 39028 7352 39080 7404
rect 39304 7352 39356 7404
rect 39856 7352 39908 7404
rect 40040 7352 40092 7404
rect 40960 7352 41012 7404
rect 53656 7352 53708 7404
rect 25688 7284 25740 7336
rect 25780 7327 25832 7336
rect 25780 7293 25789 7327
rect 25789 7293 25823 7327
rect 25823 7293 25832 7327
rect 25964 7327 26016 7336
rect 25780 7284 25832 7293
rect 25964 7293 25973 7327
rect 25973 7293 26007 7327
rect 26007 7293 26016 7327
rect 25964 7284 26016 7293
rect 26608 7284 26660 7336
rect 31852 7284 31904 7336
rect 38292 7284 38344 7336
rect 38476 7284 38528 7336
rect 42708 7284 42760 7336
rect 38660 7216 38712 7268
rect 38752 7216 38804 7268
rect 46572 7284 46624 7336
rect 49056 7284 49108 7336
rect 49424 7327 49476 7336
rect 49424 7293 49433 7327
rect 49433 7293 49467 7327
rect 49467 7293 49476 7327
rect 49424 7284 49476 7293
rect 49608 7327 49660 7336
rect 49608 7293 49617 7327
rect 49617 7293 49651 7327
rect 49651 7293 49660 7327
rect 49608 7284 49660 7293
rect 18052 7148 18104 7200
rect 20168 7148 20220 7200
rect 25964 7148 26016 7200
rect 48872 7216 48924 7268
rect 46296 7148 46348 7200
rect 48964 7148 49016 7200
rect 49700 7148 49752 7200
rect 50068 7284 50120 7336
rect 57704 7420 57756 7472
rect 58900 7420 58952 7472
rect 62948 7420 63000 7472
rect 64788 7420 64840 7472
rect 64972 7420 65024 7472
rect 61568 7352 61620 7404
rect 69480 7352 69532 7404
rect 61844 7284 61896 7336
rect 78680 7488 78732 7540
rect 71228 7420 71280 7472
rect 77852 7420 77904 7472
rect 82452 7420 82504 7472
rect 87236 7420 87288 7472
rect 87052 7395 87104 7404
rect 87052 7361 87061 7395
rect 87061 7361 87095 7395
rect 87095 7361 87104 7395
rect 87052 7352 87104 7361
rect 84200 7284 84252 7336
rect 97724 7284 97776 7336
rect 86684 7216 86736 7268
rect 50160 7148 50212 7200
rect 59912 7148 59964 7200
rect 77944 7148 77996 7200
rect 83924 7148 83976 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 50326 7046 50378 7098
rect 50390 7046 50442 7098
rect 50454 7046 50506 7098
rect 50518 7046 50570 7098
rect 81046 7046 81098 7098
rect 81110 7046 81162 7098
rect 81174 7046 81226 7098
rect 81238 7046 81290 7098
rect 3148 6944 3200 6996
rect 19340 6944 19392 6996
rect 20444 6944 20496 6996
rect 34244 6944 34296 6996
rect 39212 6944 39264 6996
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 34428 6876 34480 6928
rect 46020 6944 46072 6996
rect 46112 6944 46164 6996
rect 68192 6944 68244 6996
rect 42156 6876 42208 6928
rect 45100 6876 45152 6928
rect 45376 6876 45428 6928
rect 49332 6876 49384 6928
rect 49700 6876 49752 6928
rect 54760 6876 54812 6928
rect 72148 6876 72200 6928
rect 10968 6808 11020 6860
rect 19432 6808 19484 6860
rect 43352 6851 43404 6860
rect 5356 6740 5408 6792
rect 6460 6740 6512 6792
rect 33876 6740 33928 6792
rect 35440 6740 35492 6792
rect 36912 6740 36964 6792
rect 43352 6817 43361 6851
rect 43361 6817 43395 6851
rect 43395 6817 43404 6851
rect 43352 6808 43404 6817
rect 48596 6808 48648 6860
rect 49976 6740 50028 6792
rect 50712 6808 50764 6860
rect 63592 6851 63644 6860
rect 63592 6817 63601 6851
rect 63601 6817 63635 6851
rect 63635 6817 63644 6851
rect 63592 6808 63644 6817
rect 71964 6808 72016 6860
rect 72608 6851 72660 6860
rect 72608 6817 72617 6851
rect 72617 6817 72651 6851
rect 72651 6817 72660 6851
rect 72608 6808 72660 6817
rect 55680 6740 55732 6792
rect 61752 6740 61804 6792
rect 68468 6740 68520 6792
rect 78404 6808 78456 6860
rect 91468 6808 91520 6860
rect 98276 6808 98328 6860
rect 80520 6740 80572 6792
rect 95884 6740 95936 6792
rect 7472 6672 7524 6724
rect 56600 6672 56652 6724
rect 6460 6604 6512 6656
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 7748 6604 7800 6656
rect 21916 6604 21968 6656
rect 22008 6604 22060 6656
rect 28356 6604 28408 6656
rect 44824 6604 44876 6656
rect 45468 6604 45520 6656
rect 50804 6604 50856 6656
rect 83188 6672 83240 6724
rect 65984 6604 66036 6656
rect 72608 6604 72660 6656
rect 81348 6604 81400 6656
rect 87604 6604 87656 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 65686 6502 65738 6554
rect 65750 6502 65802 6554
rect 65814 6502 65866 6554
rect 65878 6502 65930 6554
rect 96406 6502 96458 6554
rect 96470 6502 96522 6554
rect 96534 6502 96586 6554
rect 96598 6502 96650 6554
rect 8392 6400 8444 6452
rect 72884 6400 72936 6452
rect 78312 6400 78364 6452
rect 93492 6400 93544 6452
rect 7196 6332 7248 6384
rect 8208 6332 8260 6384
rect 9128 6332 9180 6384
rect 15200 6332 15252 6384
rect 5356 6264 5408 6316
rect 11520 6264 11572 6316
rect 15476 6307 15528 6316
rect 3516 6196 3568 6248
rect 3976 6196 4028 6248
rect 6552 6196 6604 6248
rect 10232 6196 10284 6248
rect 15476 6273 15485 6307
rect 15485 6273 15519 6307
rect 15519 6273 15528 6307
rect 15476 6264 15528 6273
rect 15752 6332 15804 6384
rect 21088 6375 21140 6384
rect 21088 6341 21097 6375
rect 21097 6341 21131 6375
rect 21131 6341 21140 6375
rect 21088 6332 21140 6341
rect 21824 6332 21876 6384
rect 21916 6332 21968 6384
rect 48412 6332 48464 6384
rect 51448 6375 51500 6384
rect 51448 6341 51457 6375
rect 51457 6341 51491 6375
rect 51491 6341 51500 6375
rect 51448 6332 51500 6341
rect 62028 6332 62080 6384
rect 94412 6332 94464 6384
rect 81348 6264 81400 6316
rect 14188 6196 14240 6248
rect 15292 6239 15344 6248
rect 15292 6205 15301 6239
rect 15301 6205 15335 6239
rect 15335 6205 15344 6239
rect 15292 6196 15344 6205
rect 15384 6239 15436 6248
rect 15384 6205 15393 6239
rect 15393 6205 15427 6239
rect 15427 6205 15436 6239
rect 15384 6196 15436 6205
rect 20352 6196 20404 6248
rect 7932 6128 7984 6180
rect 11888 6128 11940 6180
rect 13544 6128 13596 6180
rect 15476 6128 15528 6180
rect 18420 6128 18472 6180
rect 21824 6196 21876 6248
rect 29000 6196 29052 6248
rect 29276 6196 29328 6248
rect 21364 6171 21416 6180
rect 7656 6060 7708 6112
rect 11612 6060 11664 6112
rect 15108 6060 15160 6112
rect 17316 6060 17368 6112
rect 20260 6060 20312 6112
rect 21364 6137 21373 6171
rect 21373 6137 21407 6171
rect 21407 6137 21416 6171
rect 21364 6128 21416 6137
rect 21640 6128 21692 6180
rect 33876 6128 33928 6180
rect 34428 6239 34480 6248
rect 34428 6205 34437 6239
rect 34437 6205 34471 6239
rect 34471 6205 34480 6239
rect 34428 6196 34480 6205
rect 42800 6196 42852 6248
rect 43812 6196 43864 6248
rect 52736 6239 52788 6248
rect 52736 6205 52745 6239
rect 52745 6205 52779 6239
rect 52779 6205 52788 6239
rect 52736 6196 52788 6205
rect 52000 6128 52052 6180
rect 20720 6103 20772 6112
rect 20720 6069 20729 6103
rect 20729 6069 20763 6103
rect 20763 6069 20772 6103
rect 20720 6060 20772 6069
rect 20812 6060 20864 6112
rect 42800 6060 42852 6112
rect 43352 6060 43404 6112
rect 51908 6060 51960 6112
rect 53196 6196 53248 6248
rect 69480 6196 69532 6248
rect 84200 6264 84252 6316
rect 86592 6307 86644 6316
rect 86592 6273 86601 6307
rect 86601 6273 86635 6307
rect 86635 6273 86644 6307
rect 86592 6264 86644 6273
rect 53656 6128 53708 6180
rect 81900 6239 81952 6248
rect 81900 6205 81909 6239
rect 81909 6205 81943 6239
rect 81943 6205 81952 6239
rect 81900 6196 81952 6205
rect 81440 6128 81492 6180
rect 84844 6196 84896 6248
rect 85948 6239 86000 6248
rect 85948 6205 85957 6239
rect 85957 6205 85991 6239
rect 85991 6205 86000 6239
rect 85948 6196 86000 6205
rect 61752 6060 61804 6112
rect 69480 6060 69532 6112
rect 97816 6264 97868 6316
rect 96988 6239 97040 6248
rect 96988 6205 96997 6239
rect 96997 6205 97031 6239
rect 97031 6205 97040 6239
rect 96988 6196 97040 6205
rect 97632 6239 97684 6248
rect 97632 6205 97641 6239
rect 97641 6205 97675 6239
rect 97675 6205 97684 6239
rect 97632 6196 97684 6205
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 50326 5958 50378 6010
rect 50390 5958 50442 6010
rect 50454 5958 50506 6010
rect 50518 5958 50570 6010
rect 81046 5958 81098 6010
rect 81110 5958 81162 6010
rect 81174 5958 81226 6010
rect 81238 5958 81290 6010
rect 1860 5720 1912 5772
rect 2780 5720 2832 5772
rect 20812 5856 20864 5908
rect 23388 5856 23440 5908
rect 71596 5856 71648 5908
rect 73896 5899 73948 5908
rect 73896 5865 73905 5899
rect 73905 5865 73939 5899
rect 73939 5865 73948 5899
rect 73896 5856 73948 5865
rect 91836 5856 91888 5908
rect 95884 5899 95936 5908
rect 6920 5720 6972 5772
rect 7656 5763 7708 5772
rect 5632 5652 5684 5704
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 11704 5788 11756 5840
rect 11888 5788 11940 5840
rect 17224 5788 17276 5840
rect 17316 5788 17368 5840
rect 22008 5788 22060 5840
rect 29736 5788 29788 5840
rect 15108 5720 15160 5772
rect 15200 5720 15252 5772
rect 21640 5720 21692 5772
rect 26516 5763 26568 5772
rect 7656 5584 7708 5636
rect 8760 5652 8812 5704
rect 22836 5652 22888 5704
rect 26240 5695 26292 5704
rect 8208 5584 8260 5636
rect 11704 5584 11756 5636
rect 23940 5584 23992 5636
rect 5080 5559 5132 5568
rect 5080 5525 5089 5559
rect 5089 5525 5123 5559
rect 5123 5525 5132 5559
rect 5080 5516 5132 5525
rect 8392 5516 8444 5568
rect 8484 5516 8536 5568
rect 15476 5516 15528 5568
rect 17224 5516 17276 5568
rect 24768 5516 24820 5568
rect 26240 5661 26249 5695
rect 26249 5661 26283 5695
rect 26283 5661 26292 5695
rect 26240 5652 26292 5661
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 32404 5720 32456 5772
rect 35992 5720 36044 5772
rect 36636 5788 36688 5840
rect 53472 5788 53524 5840
rect 58532 5788 58584 5840
rect 34796 5652 34848 5704
rect 37648 5584 37700 5636
rect 40684 5584 40736 5636
rect 44916 5720 44968 5772
rect 58992 5720 59044 5772
rect 74080 5763 74132 5772
rect 74080 5729 74089 5763
rect 74089 5729 74123 5763
rect 74123 5729 74132 5763
rect 74080 5720 74132 5729
rect 95332 5720 95384 5772
rect 95884 5865 95893 5899
rect 95893 5865 95927 5899
rect 95927 5865 95936 5899
rect 95884 5856 95936 5865
rect 46756 5652 46808 5704
rect 59452 5652 59504 5704
rect 83740 5652 83792 5704
rect 91468 5652 91520 5704
rect 31116 5516 31168 5568
rect 34060 5516 34112 5568
rect 36544 5516 36596 5568
rect 46204 5516 46256 5568
rect 52828 5516 52880 5568
rect 67640 5584 67692 5636
rect 69940 5584 69992 5636
rect 61476 5516 61528 5568
rect 62764 5516 62816 5568
rect 73988 5516 74040 5568
rect 76564 5516 76616 5568
rect 89352 5584 89404 5636
rect 96252 5720 96304 5772
rect 99012 5720 99064 5772
rect 95332 5516 95384 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 65686 5414 65738 5466
rect 65750 5414 65802 5466
rect 65814 5414 65866 5466
rect 65878 5414 65930 5466
rect 96406 5414 96458 5466
rect 96470 5414 96522 5466
rect 96534 5414 96586 5466
rect 96598 5414 96650 5466
rect 7564 5312 7616 5364
rect 16028 5312 16080 5364
rect 24308 5355 24360 5364
rect 5264 5108 5316 5160
rect 6736 5108 6788 5160
rect 8300 5108 8352 5160
rect 2044 5040 2096 5092
rect 480 4972 532 5024
rect 3424 5015 3476 5024
rect 3424 4981 3433 5015
rect 3433 4981 3467 5015
rect 3467 4981 3476 5015
rect 3424 4972 3476 4981
rect 4896 4972 4948 5024
rect 5632 4972 5684 5024
rect 8208 4972 8260 5024
rect 22928 5244 22980 5296
rect 24308 5321 24317 5355
rect 24317 5321 24351 5355
rect 24351 5321 24360 5355
rect 24308 5312 24360 5321
rect 29276 5244 29328 5296
rect 23204 5219 23256 5228
rect 9128 5151 9180 5160
rect 9128 5117 9137 5151
rect 9137 5117 9171 5151
rect 9171 5117 9180 5151
rect 9128 5108 9180 5117
rect 21732 5108 21784 5160
rect 23204 5185 23213 5219
rect 23213 5185 23247 5219
rect 23247 5185 23256 5219
rect 23204 5176 23256 5185
rect 31392 5176 31444 5228
rect 25044 5151 25096 5160
rect 25044 5117 25053 5151
rect 25053 5117 25087 5151
rect 25087 5117 25096 5151
rect 25044 5108 25096 5117
rect 25688 5151 25740 5160
rect 25688 5117 25697 5151
rect 25697 5117 25731 5151
rect 25731 5117 25740 5151
rect 25688 5108 25740 5117
rect 26332 5151 26384 5160
rect 26332 5117 26341 5151
rect 26341 5117 26375 5151
rect 26375 5117 26384 5151
rect 26332 5108 26384 5117
rect 27804 5151 27856 5160
rect 27804 5117 27813 5151
rect 27813 5117 27847 5151
rect 27847 5117 27856 5151
rect 27804 5108 27856 5117
rect 33508 5108 33560 5160
rect 18604 5040 18656 5092
rect 31668 5040 31720 5092
rect 34612 5244 34664 5296
rect 38016 5244 38068 5296
rect 43444 5176 43496 5228
rect 34152 5151 34204 5160
rect 34152 5117 34161 5151
rect 34161 5117 34195 5151
rect 34195 5117 34204 5151
rect 34152 5108 34204 5117
rect 36636 5151 36688 5160
rect 36636 5117 36645 5151
rect 36645 5117 36679 5151
rect 36679 5117 36688 5151
rect 36636 5108 36688 5117
rect 36820 5151 36872 5160
rect 36820 5117 36829 5151
rect 36829 5117 36863 5151
rect 36863 5117 36872 5151
rect 36820 5108 36872 5117
rect 37188 5108 37240 5160
rect 38752 5151 38804 5160
rect 38752 5117 38761 5151
rect 38761 5117 38795 5151
rect 38795 5117 38804 5151
rect 38752 5108 38804 5117
rect 39212 5151 39264 5160
rect 39212 5117 39221 5151
rect 39221 5117 39255 5151
rect 39255 5117 39264 5151
rect 39212 5108 39264 5117
rect 45008 5176 45060 5228
rect 45284 5219 45336 5228
rect 45284 5185 45293 5219
rect 45293 5185 45327 5219
rect 45327 5185 45336 5219
rect 45284 5176 45336 5185
rect 46296 5244 46348 5296
rect 55772 5244 55824 5296
rect 55956 5312 56008 5364
rect 66168 5312 66220 5364
rect 73988 5312 74040 5364
rect 74080 5312 74132 5364
rect 82176 5312 82228 5364
rect 90824 5312 90876 5364
rect 52000 5176 52052 5228
rect 52184 5176 52236 5228
rect 55864 5176 55916 5228
rect 36452 5015 36504 5024
rect 36452 4981 36461 5015
rect 36461 4981 36495 5015
rect 36495 4981 36504 5015
rect 36452 4972 36504 4981
rect 36820 4972 36872 5024
rect 44088 5040 44140 5092
rect 54576 5108 54628 5160
rect 57888 5244 57940 5296
rect 64972 5244 65024 5296
rect 65156 5244 65208 5296
rect 65524 5244 65576 5296
rect 67088 5244 67140 5296
rect 68100 5244 68152 5296
rect 68560 5244 68612 5296
rect 56232 5176 56284 5228
rect 59084 5176 59136 5228
rect 65340 5176 65392 5228
rect 71044 5176 71096 5228
rect 58900 5108 58952 5160
rect 64604 5108 64656 5160
rect 64880 5151 64932 5160
rect 64880 5117 64889 5151
rect 64889 5117 64923 5151
rect 64923 5117 64932 5151
rect 64880 5108 64932 5117
rect 65064 5151 65116 5160
rect 65064 5117 65073 5151
rect 65073 5117 65107 5151
rect 65107 5117 65116 5151
rect 65064 5108 65116 5117
rect 65156 5108 65208 5160
rect 82176 5176 82228 5228
rect 82636 5176 82688 5228
rect 76932 5151 76984 5160
rect 76932 5117 76941 5151
rect 76941 5117 76975 5151
rect 76975 5117 76984 5151
rect 76932 5108 76984 5117
rect 77484 5108 77536 5160
rect 87328 5151 87380 5160
rect 87328 5117 87337 5151
rect 87337 5117 87371 5151
rect 87371 5117 87380 5151
rect 87328 5108 87380 5117
rect 87604 5151 87656 5160
rect 87604 5117 87613 5151
rect 87613 5117 87647 5151
rect 87647 5117 87656 5151
rect 87604 5108 87656 5117
rect 59268 5040 59320 5092
rect 64788 5040 64840 5092
rect 52000 4972 52052 5024
rect 65524 4972 65576 5024
rect 68836 4972 68888 5024
rect 82176 5040 82228 5092
rect 87236 4972 87288 5024
rect 88524 5108 88576 5160
rect 90732 5151 90784 5160
rect 90732 5117 90741 5151
rect 90741 5117 90775 5151
rect 90775 5117 90784 5151
rect 90732 5108 90784 5117
rect 90824 5108 90876 5160
rect 91468 5151 91520 5160
rect 91468 5117 91477 5151
rect 91477 5117 91511 5151
rect 91511 5117 91520 5151
rect 91468 5108 91520 5117
rect 92940 5151 92992 5160
rect 92940 5117 92949 5151
rect 92949 5117 92983 5151
rect 92983 5117 92992 5151
rect 92940 5108 92992 5117
rect 91836 5040 91888 5092
rect 89812 4972 89864 5024
rect 95700 5108 95752 5160
rect 97816 5151 97868 5160
rect 95240 5040 95292 5092
rect 97816 5117 97825 5151
rect 97825 5117 97859 5151
rect 97859 5117 97868 5151
rect 97816 5108 97868 5117
rect 98460 5040 98512 5092
rect 96160 4972 96212 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 50326 4870 50378 4922
rect 50390 4870 50442 4922
rect 50454 4870 50506 4922
rect 50518 4870 50570 4922
rect 81046 4870 81098 4922
rect 81110 4870 81162 4922
rect 81174 4870 81226 4922
rect 81238 4870 81290 4922
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 2504 4811 2556 4820
rect 2504 4777 2513 4811
rect 2513 4777 2547 4811
rect 2547 4777 2556 4811
rect 2504 4768 2556 4777
rect 6644 4743 6696 4752
rect 6644 4709 6653 4743
rect 6653 4709 6687 4743
rect 6687 4709 6696 4743
rect 6644 4700 6696 4709
rect 848 4632 900 4684
rect 8944 4768 8996 4820
rect 25136 4768 25188 4820
rect 7288 4743 7340 4752
rect 7288 4709 7297 4743
rect 7297 4709 7331 4743
rect 7331 4709 7340 4743
rect 7288 4700 7340 4709
rect 8116 4700 8168 4752
rect 20076 4700 20128 4752
rect 24952 4700 25004 4752
rect 25320 4700 25372 4752
rect 25964 4700 26016 4752
rect 8852 4632 8904 4684
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 11888 4675 11940 4684
rect 11888 4641 11897 4675
rect 11897 4641 11931 4675
rect 11931 4641 11940 4675
rect 11888 4632 11940 4641
rect 12440 4632 12492 4684
rect 14280 4632 14332 4684
rect 15200 4632 15252 4684
rect 16120 4675 16172 4684
rect 16120 4641 16129 4675
rect 16129 4641 16163 4675
rect 16163 4641 16172 4675
rect 16120 4632 16172 4641
rect 17316 4675 17368 4684
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 17960 4675 18012 4684
rect 17960 4641 17969 4675
rect 17969 4641 18003 4675
rect 18003 4641 18012 4675
rect 17960 4632 18012 4641
rect 18604 4675 18656 4684
rect 18604 4641 18613 4675
rect 18613 4641 18647 4675
rect 18647 4641 18656 4675
rect 18604 4632 18656 4641
rect 19892 4632 19944 4684
rect 20996 4675 21048 4684
rect 20996 4641 21005 4675
rect 21005 4641 21039 4675
rect 21039 4641 21048 4675
rect 20996 4632 21048 4641
rect 21732 4632 21784 4684
rect 22652 4675 22704 4684
rect 22652 4641 22661 4675
rect 22661 4641 22695 4675
rect 22695 4641 22704 4675
rect 22652 4632 22704 4641
rect 23204 4632 23256 4684
rect 25872 4632 25924 4684
rect 26056 4675 26108 4684
rect 26056 4641 26065 4675
rect 26065 4641 26099 4675
rect 26099 4641 26108 4675
rect 26056 4632 26108 4641
rect 27436 4700 27488 4752
rect 32956 4768 33008 4820
rect 33324 4768 33376 4820
rect 37372 4768 37424 4820
rect 52920 4768 52972 4820
rect 36544 4700 36596 4752
rect 39948 4700 40000 4752
rect 50988 4700 51040 4752
rect 26884 4632 26936 4684
rect 27068 4632 27120 4684
rect 29092 4675 29144 4684
rect 29092 4641 29101 4675
rect 29101 4641 29135 4675
rect 29135 4641 29144 4675
rect 29092 4632 29144 4641
rect 32956 4632 33008 4684
rect 34244 4675 34296 4684
rect 34244 4641 34253 4675
rect 34253 4641 34287 4675
rect 34287 4641 34296 4675
rect 34244 4632 34296 4641
rect 36084 4675 36136 4684
rect 36084 4641 36093 4675
rect 36093 4641 36127 4675
rect 36127 4641 36136 4675
rect 36084 4632 36136 4641
rect 36636 4632 36688 4684
rect 37648 4675 37700 4684
rect 37648 4641 37657 4675
rect 37657 4641 37691 4675
rect 37691 4641 37700 4675
rect 37648 4632 37700 4641
rect 39488 4675 39540 4684
rect 39488 4641 39497 4675
rect 39497 4641 39531 4675
rect 39531 4641 39540 4675
rect 39488 4632 39540 4641
rect 40316 4632 40368 4684
rect 41512 4632 41564 4684
rect 43996 4675 44048 4684
rect 43996 4641 44005 4675
rect 44005 4641 44039 4675
rect 44039 4641 44048 4675
rect 43996 4632 44048 4641
rect 44548 4632 44600 4684
rect 45836 4632 45888 4684
rect 47032 4675 47084 4684
rect 47032 4641 47041 4675
rect 47041 4641 47075 4675
rect 47075 4641 47084 4675
rect 47032 4632 47084 4641
rect 47584 4632 47636 4684
rect 49240 4632 49292 4684
rect 52368 4632 52420 4684
rect 52552 4675 52604 4684
rect 52552 4641 52561 4675
rect 52561 4641 52595 4675
rect 52595 4641 52604 4675
rect 52552 4632 52604 4641
rect 53472 4675 53524 4684
rect 53472 4641 53481 4675
rect 53481 4641 53515 4675
rect 53515 4641 53524 4675
rect 53472 4632 53524 4641
rect 53656 4675 53708 4684
rect 53656 4641 53665 4675
rect 53665 4641 53699 4675
rect 53699 4641 53708 4675
rect 53656 4632 53708 4641
rect 54300 4675 54352 4684
rect 54300 4641 54309 4675
rect 54309 4641 54343 4675
rect 54343 4641 54352 4675
rect 54300 4632 54352 4641
rect 6184 4564 6236 4616
rect 8300 4564 8352 4616
rect 21180 4564 21232 4616
rect 1676 4496 1728 4548
rect 7104 4539 7156 4548
rect 7104 4505 7113 4539
rect 7113 4505 7147 4539
rect 7147 4505 7156 4539
rect 7104 4496 7156 4505
rect 7380 4496 7432 4548
rect 19984 4496 20036 4548
rect 22836 4496 22888 4548
rect 36452 4564 36504 4616
rect 37740 4564 37792 4616
rect 49516 4564 49568 4616
rect 55128 4700 55180 4752
rect 62028 4700 62080 4752
rect 55312 4632 55364 4684
rect 57336 4632 57388 4684
rect 61844 4632 61896 4684
rect 62396 4700 62448 4752
rect 66168 4700 66220 4752
rect 71044 4700 71096 4752
rect 78220 4743 78272 4752
rect 62304 4675 62356 4684
rect 62304 4641 62313 4675
rect 62313 4641 62347 4675
rect 62347 4641 62356 4675
rect 62304 4632 62356 4641
rect 62580 4632 62632 4684
rect 64236 4675 64288 4684
rect 64236 4641 64245 4675
rect 64245 4641 64279 4675
rect 64279 4641 64288 4675
rect 64236 4632 64288 4641
rect 64328 4632 64380 4684
rect 65432 4632 65484 4684
rect 65984 4632 66036 4684
rect 68376 4675 68428 4684
rect 68376 4641 68385 4675
rect 68385 4641 68419 4675
rect 68419 4641 68428 4675
rect 68376 4632 68428 4641
rect 70768 4675 70820 4684
rect 70768 4641 70777 4675
rect 70777 4641 70811 4675
rect 70811 4641 70820 4675
rect 70768 4632 70820 4641
rect 73804 4675 73856 4684
rect 73804 4641 73813 4675
rect 73813 4641 73847 4675
rect 73847 4641 73856 4675
rect 73804 4632 73856 4641
rect 76288 4675 76340 4684
rect 76288 4641 76297 4675
rect 76297 4641 76331 4675
rect 76331 4641 76340 4675
rect 76288 4632 76340 4641
rect 77944 4675 77996 4684
rect 77944 4641 77953 4675
rect 77953 4641 77987 4675
rect 77987 4641 77996 4675
rect 77944 4632 77996 4641
rect 78220 4709 78229 4743
rect 78229 4709 78263 4743
rect 78263 4709 78272 4743
rect 78220 4700 78272 4709
rect 78404 4768 78456 4820
rect 97540 4768 97592 4820
rect 78680 4675 78732 4684
rect 78680 4641 78689 4675
rect 78689 4641 78723 4675
rect 78723 4641 78732 4675
rect 78680 4632 78732 4641
rect 78772 4632 78824 4684
rect 79416 4632 79468 4684
rect 80060 4632 80112 4684
rect 82912 4675 82964 4684
rect 8208 4428 8260 4480
rect 28632 4471 28684 4480
rect 28632 4437 28641 4471
rect 28641 4437 28675 4471
rect 28675 4437 28684 4471
rect 28632 4428 28684 4437
rect 33048 4428 33100 4480
rect 36820 4428 36872 4480
rect 52092 4496 52144 4548
rect 42156 4428 42208 4480
rect 46388 4428 46440 4480
rect 61016 4564 61068 4616
rect 63868 4564 63920 4616
rect 58256 4496 58308 4548
rect 62120 4496 62172 4548
rect 62856 4496 62908 4548
rect 64420 4564 64472 4616
rect 64972 4496 65024 4548
rect 78956 4564 79008 4616
rect 78404 4496 78456 4548
rect 80520 4564 80572 4616
rect 82912 4641 82921 4675
rect 82921 4641 82955 4675
rect 82955 4641 82964 4675
rect 82912 4632 82964 4641
rect 83556 4675 83608 4684
rect 83556 4641 83565 4675
rect 83565 4641 83599 4675
rect 83599 4641 83608 4675
rect 83556 4632 83608 4641
rect 84292 4700 84344 4752
rect 85488 4700 85540 4752
rect 87604 4700 87656 4752
rect 85396 4675 85448 4684
rect 85396 4641 85405 4675
rect 85405 4641 85439 4675
rect 85439 4641 85448 4675
rect 85396 4632 85448 4641
rect 86040 4675 86092 4684
rect 86040 4641 86049 4675
rect 86049 4641 86083 4675
rect 86083 4641 86092 4675
rect 86040 4632 86092 4641
rect 86960 4632 87012 4684
rect 88800 4675 88852 4684
rect 88800 4641 88809 4675
rect 88809 4641 88843 4675
rect 88843 4641 88852 4675
rect 88800 4632 88852 4641
rect 89076 4632 89128 4684
rect 89720 4632 89772 4684
rect 90272 4632 90324 4684
rect 91100 4632 91152 4684
rect 91652 4632 91704 4684
rect 92756 4632 92808 4684
rect 93860 4632 93912 4684
rect 94228 4632 94280 4684
rect 95332 4675 95384 4684
rect 95332 4641 95341 4675
rect 95341 4641 95375 4675
rect 95375 4641 95384 4675
rect 95332 4632 95384 4641
rect 95976 4675 96028 4684
rect 95976 4641 95985 4675
rect 95985 4641 96019 4675
rect 96019 4641 96028 4675
rect 95976 4632 96028 4641
rect 96712 4632 96764 4684
rect 97264 4675 97316 4684
rect 97264 4641 97273 4675
rect 97273 4641 97307 4675
rect 97307 4641 97316 4675
rect 97264 4632 97316 4641
rect 88340 4564 88392 4616
rect 90732 4496 90784 4548
rect 53472 4428 53524 4480
rect 62028 4428 62080 4480
rect 62304 4428 62356 4480
rect 67640 4428 67692 4480
rect 74172 4428 74224 4480
rect 89352 4428 89404 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 65686 4326 65738 4378
rect 65750 4326 65802 4378
rect 65814 4326 65866 4378
rect 65878 4326 65930 4378
rect 96406 4326 96458 4378
rect 96470 4326 96522 4378
rect 96534 4326 96586 4378
rect 96598 4326 96650 4378
rect 2964 4131 3016 4140
rect 2964 4097 2973 4131
rect 2973 4097 3007 4131
rect 3007 4097 3016 4131
rect 2964 4088 3016 4097
rect 5264 4088 5316 4140
rect 6184 4088 6236 4140
rect 7104 4088 7156 4140
rect 1216 4020 1268 4072
rect 3148 4020 3200 4072
rect 4712 4063 4764 4072
rect 4712 4029 4721 4063
rect 4721 4029 4755 4063
rect 4755 4029 4764 4063
rect 4712 4020 4764 4029
rect 664 3952 716 4004
rect 2228 3995 2280 4004
rect 2228 3961 2237 3995
rect 2237 3961 2271 3995
rect 2271 3961 2280 3995
rect 2228 3952 2280 3961
rect 3332 3952 3384 4004
rect 5448 4020 5500 4072
rect 6552 4020 6604 4072
rect 7748 4063 7800 4072
rect 7748 4029 7757 4063
rect 7757 4029 7791 4063
rect 7791 4029 7800 4063
rect 7748 4020 7800 4029
rect 5264 3952 5316 4004
rect 9404 4063 9456 4072
rect 9404 4029 9413 4063
rect 9413 4029 9447 4063
rect 9447 4029 9456 4063
rect 9404 4020 9456 4029
rect 9496 4020 9548 4072
rect 10140 4020 10192 4072
rect 11428 4020 11480 4072
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 13176 4020 13228 4029
rect 5080 3884 5132 3936
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 7840 3884 7892 3936
rect 8576 3884 8628 3936
rect 8944 3884 8996 3936
rect 12256 3884 12308 3936
rect 13084 3952 13136 4004
rect 13728 4020 13780 4072
rect 15476 4020 15528 4072
rect 33508 4224 33560 4276
rect 46296 4224 46348 4276
rect 47952 4224 48004 4276
rect 21916 4156 21968 4208
rect 33140 4156 33192 4208
rect 16764 4020 16816 4072
rect 18328 4020 18380 4072
rect 19248 4020 19300 4072
rect 23020 4063 23072 4072
rect 18788 3952 18840 4004
rect 19156 3995 19208 4004
rect 19156 3961 19165 3995
rect 19165 3961 19199 3995
rect 19199 3961 19208 3995
rect 19156 3952 19208 3961
rect 20352 3952 20404 4004
rect 23020 4029 23029 4063
rect 23029 4029 23063 4063
rect 23063 4029 23072 4063
rect 23020 4020 23072 4029
rect 23480 4063 23532 4072
rect 23480 4029 23489 4063
rect 23489 4029 23523 4063
rect 23523 4029 23532 4063
rect 23480 4020 23532 4029
rect 23848 4020 23900 4072
rect 24492 4020 24544 4072
rect 25964 4020 26016 4072
rect 15292 3884 15344 3936
rect 16028 3884 16080 3936
rect 18328 3884 18380 3936
rect 18972 3884 19024 3936
rect 19340 3884 19392 3936
rect 25320 3952 25372 4004
rect 25780 3952 25832 4004
rect 26516 4020 26568 4072
rect 28080 4020 28132 4072
rect 28724 4020 28776 4072
rect 29368 4020 29420 4072
rect 31208 4063 31260 4072
rect 31208 4029 31217 4063
rect 31217 4029 31251 4063
rect 31251 4029 31260 4063
rect 31208 4020 31260 4029
rect 26424 3952 26476 4004
rect 29920 3952 29972 4004
rect 23388 3884 23440 3936
rect 26884 3884 26936 3936
rect 27804 3884 27856 3936
rect 35624 4088 35676 4140
rect 37280 4088 37332 4140
rect 32956 4020 33008 4072
rect 33600 4020 33652 4072
rect 34336 4020 34388 4072
rect 34796 4020 34848 4072
rect 35716 4020 35768 4072
rect 36820 4063 36872 4072
rect 36820 4029 36829 4063
rect 36829 4029 36863 4063
rect 36863 4029 36872 4063
rect 36820 4020 36872 4029
rect 38660 4063 38712 4072
rect 38660 4029 38669 4063
rect 38669 4029 38703 4063
rect 38703 4029 38712 4063
rect 38660 4020 38712 4029
rect 39396 4088 39448 4140
rect 39948 4063 40000 4072
rect 39948 4029 39957 4063
rect 39957 4029 39991 4063
rect 39991 4029 40000 4063
rect 39948 4020 40000 4029
rect 38568 3952 38620 4004
rect 39212 3952 39264 4004
rect 39672 3952 39724 4004
rect 40960 3952 41012 4004
rect 36360 3884 36412 3936
rect 36544 3884 36596 3936
rect 42340 3884 42392 3936
rect 42708 4156 42760 4208
rect 48504 4156 48556 4208
rect 55772 4088 55824 4140
rect 42708 4020 42760 4072
rect 45376 4063 45428 4072
rect 43352 3952 43404 4004
rect 45376 4029 45385 4063
rect 45385 4029 45419 4063
rect 45419 4029 45428 4063
rect 45376 4020 45428 4029
rect 46020 4063 46072 4072
rect 46020 4029 46029 4063
rect 46029 4029 46063 4063
rect 46063 4029 46072 4063
rect 46020 4020 46072 4029
rect 45192 3952 45244 4004
rect 46388 3952 46440 4004
rect 48228 4020 48280 4072
rect 48872 4020 48924 4072
rect 49516 4020 49568 4072
rect 50160 4020 50212 4072
rect 50804 4020 50856 4072
rect 51264 3952 51316 4004
rect 52644 4063 52696 4072
rect 52644 4029 52653 4063
rect 52653 4029 52687 4063
rect 52687 4029 52696 4063
rect 52644 4020 52696 4029
rect 53104 4020 53156 4072
rect 53656 3952 53708 4004
rect 54944 4020 54996 4072
rect 55588 4020 55640 4072
rect 56232 4020 56284 4072
rect 56784 4020 56836 4072
rect 57428 4020 57480 4072
rect 60924 4088 60976 4140
rect 61016 4088 61068 4140
rect 58624 4020 58676 4072
rect 52828 3884 52880 3936
rect 53932 3884 53984 3936
rect 59084 3952 59136 4004
rect 59820 3952 59872 4004
rect 60740 4020 60792 4072
rect 62304 4088 62356 4140
rect 62028 4020 62080 4072
rect 63500 4088 63552 4140
rect 63224 4020 63276 4072
rect 64788 4088 64840 4140
rect 65340 4088 65392 4140
rect 69572 4088 69624 4140
rect 66536 4020 66588 4072
rect 67180 4020 67232 4072
rect 67824 4020 67876 4072
rect 68928 4020 68980 4072
rect 70216 4088 70268 4140
rect 87144 4088 87196 4140
rect 90640 4088 90692 4140
rect 71412 4020 71464 4072
rect 72056 4020 72108 4072
rect 72608 4020 72660 4072
rect 73252 4020 73304 4072
rect 74448 4020 74500 4072
rect 75092 4020 75144 4072
rect 75736 4020 75788 4072
rect 77116 4063 77168 4072
rect 77116 4029 77125 4063
rect 77125 4029 77159 4063
rect 77159 4029 77168 4063
rect 77116 4020 77168 4029
rect 78312 4063 78364 4072
rect 78312 4029 78321 4063
rect 78321 4029 78355 4063
rect 78355 4029 78364 4063
rect 78312 4020 78364 4029
rect 78956 4063 79008 4072
rect 78956 4029 78965 4063
rect 78965 4029 78999 4063
rect 78999 4029 79008 4063
rect 78956 4020 79008 4029
rect 80796 4063 80848 4072
rect 80796 4029 80805 4063
rect 80805 4029 80839 4063
rect 80839 4029 80848 4063
rect 80796 4020 80848 4029
rect 81348 4020 81400 4072
rect 81992 4020 82044 4072
rect 82728 4063 82780 4072
rect 82728 4029 82737 4063
rect 82737 4029 82771 4063
rect 82771 4029 82780 4063
rect 82728 4020 82780 4029
rect 83648 4063 83700 4072
rect 83648 4029 83657 4063
rect 83657 4029 83691 4063
rect 83691 4029 83700 4063
rect 83648 4020 83700 4029
rect 84200 4020 84252 4072
rect 84844 4020 84896 4072
rect 87604 4020 87656 4072
rect 91192 4063 91244 4072
rect 60924 3952 60976 4004
rect 80888 3952 80940 4004
rect 85672 3952 85724 4004
rect 55680 3884 55732 3936
rect 91192 4029 91201 4063
rect 91201 4029 91235 4063
rect 91235 4029 91244 4063
rect 91192 4020 91244 4029
rect 91376 4063 91428 4072
rect 91376 4029 91385 4063
rect 91385 4029 91419 4063
rect 91419 4029 91428 4063
rect 91376 4020 91428 4029
rect 92020 4088 92072 4140
rect 97080 4088 97132 4140
rect 91744 3952 91796 4004
rect 92388 4020 92440 4072
rect 93584 4020 93636 4072
rect 94136 4020 94188 4072
rect 95424 4020 95476 4072
rect 97908 4063 97960 4072
rect 97908 4029 97917 4063
rect 97917 4029 97951 4063
rect 97951 4029 97960 4063
rect 97908 4020 97960 4029
rect 99288 3952 99340 4004
rect 98000 3927 98052 3936
rect 98000 3893 98009 3927
rect 98009 3893 98043 3927
rect 98043 3893 98052 3927
rect 98000 3884 98052 3893
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 50326 3782 50378 3834
rect 50390 3782 50442 3834
rect 50454 3782 50506 3834
rect 50518 3782 50570 3834
rect 81046 3782 81098 3834
rect 81110 3782 81162 3834
rect 81174 3782 81226 3834
rect 81238 3782 81290 3834
rect 5080 3680 5132 3732
rect 5356 3680 5408 3732
rect 11152 3680 11204 3732
rect 3056 3655 3108 3664
rect 3056 3621 3065 3655
rect 3065 3621 3099 3655
rect 3099 3621 3108 3655
rect 3056 3612 3108 3621
rect 4804 3612 4856 3664
rect 5540 3655 5592 3664
rect 5540 3621 5549 3655
rect 5549 3621 5583 3655
rect 5583 3621 5592 3655
rect 5540 3612 5592 3621
rect 6276 3655 6328 3664
rect 6276 3621 6285 3655
rect 6285 3621 6319 3655
rect 6319 3621 6328 3655
rect 6276 3612 6328 3621
rect 8024 3612 8076 3664
rect 1952 3544 2004 3596
rect 112 3476 164 3528
rect 1124 3476 1176 3528
rect 2412 3476 2464 3528
rect 1308 3408 1360 3460
rect 3884 3544 3936 3596
rect 5356 3544 5408 3596
rect 7196 3544 7248 3596
rect 9956 3612 10008 3664
rect 13268 3655 13320 3664
rect 13268 3621 13277 3655
rect 13277 3621 13311 3655
rect 13311 3621 13320 3655
rect 13268 3612 13320 3621
rect 10324 3587 10376 3596
rect 8024 3476 8076 3528
rect 8944 3476 8996 3528
rect 10324 3553 10333 3587
rect 10333 3553 10367 3587
rect 10367 3553 10376 3587
rect 10324 3544 10376 3553
rect 13636 3544 13688 3596
rect 19340 3680 19392 3732
rect 20628 3680 20680 3732
rect 17592 3612 17644 3664
rect 17868 3655 17920 3664
rect 17868 3621 17894 3655
rect 17894 3621 17920 3655
rect 17868 3612 17920 3621
rect 18144 3612 18196 3664
rect 20168 3612 20220 3664
rect 27528 3680 27580 3732
rect 29092 3680 29144 3732
rect 34704 3680 34756 3732
rect 21548 3655 21600 3664
rect 21548 3621 21557 3655
rect 21557 3621 21591 3655
rect 21591 3621 21600 3655
rect 21548 3612 21600 3621
rect 21824 3612 21876 3664
rect 36544 3612 36596 3664
rect 16212 3544 16264 3596
rect 17040 3544 17092 3596
rect 16672 3476 16724 3528
rect 17224 3544 17276 3596
rect 18512 3587 18564 3596
rect 18512 3553 18521 3587
rect 18521 3553 18555 3587
rect 18555 3553 18564 3587
rect 18512 3544 18564 3553
rect 20076 3587 20128 3596
rect 20076 3553 20085 3587
rect 20085 3553 20119 3587
rect 20119 3553 20128 3587
rect 20076 3544 20128 3553
rect 21180 3544 21232 3596
rect 21916 3544 21968 3596
rect 22836 3587 22888 3596
rect 22836 3553 22845 3587
rect 22845 3553 22879 3587
rect 22879 3553 22888 3587
rect 22836 3544 22888 3553
rect 24032 3587 24084 3596
rect 24032 3553 24041 3587
rect 24041 3553 24075 3587
rect 24075 3553 24084 3587
rect 24032 3544 24084 3553
rect 24676 3544 24728 3596
rect 25320 3544 25372 3596
rect 26792 3587 26844 3596
rect 26792 3553 26801 3587
rect 26801 3553 26835 3587
rect 26835 3553 26844 3587
rect 26792 3544 26844 3553
rect 27712 3587 27764 3596
rect 27712 3553 27721 3587
rect 27721 3553 27755 3587
rect 27755 3553 27764 3587
rect 27712 3544 27764 3553
rect 28908 3587 28960 3596
rect 28908 3553 28917 3587
rect 28917 3553 28951 3587
rect 28951 3553 28960 3587
rect 28908 3544 28960 3553
rect 29920 3544 29972 3596
rect 30564 3544 30616 3596
rect 31944 3587 31996 3596
rect 31944 3553 31953 3587
rect 31953 3553 31987 3587
rect 31987 3553 31996 3587
rect 31944 3544 31996 3553
rect 17868 3476 17920 3528
rect 13268 3408 13320 3460
rect 13452 3408 13504 3460
rect 14464 3408 14516 3460
rect 14740 3408 14792 3460
rect 16488 3408 16540 3460
rect 17132 3408 17184 3460
rect 9220 3340 9272 3392
rect 9864 3340 9916 3392
rect 10508 3340 10560 3392
rect 11612 3340 11664 3392
rect 12900 3340 12952 3392
rect 14096 3340 14148 3392
rect 16028 3340 16080 3392
rect 20628 3476 20680 3528
rect 22284 3476 22336 3528
rect 18236 3408 18288 3460
rect 18144 3340 18196 3392
rect 19432 3340 19484 3392
rect 20812 3408 20864 3460
rect 22008 3408 22060 3460
rect 25596 3408 25648 3460
rect 31852 3476 31904 3528
rect 32864 3544 32916 3596
rect 34428 3587 34480 3596
rect 34428 3553 34437 3587
rect 34437 3553 34471 3587
rect 34471 3553 34480 3587
rect 34428 3544 34480 3553
rect 35440 3544 35492 3596
rect 37464 3680 37516 3732
rect 37832 3680 37884 3732
rect 39488 3680 39540 3732
rect 49700 3680 49752 3732
rect 44640 3612 44692 3664
rect 45100 3612 45152 3664
rect 48688 3612 48740 3664
rect 49608 3612 49660 3664
rect 76380 3680 76432 3732
rect 78128 3680 78180 3732
rect 78680 3680 78732 3732
rect 79324 3680 79376 3732
rect 62488 3612 62540 3664
rect 37740 3587 37792 3596
rect 35624 3476 35676 3528
rect 37740 3553 37749 3587
rect 37749 3553 37783 3587
rect 37783 3553 37792 3587
rect 37740 3544 37792 3553
rect 38108 3544 38160 3596
rect 39304 3544 39356 3596
rect 40500 3544 40552 3596
rect 41696 3587 41748 3596
rect 41696 3553 41705 3587
rect 41705 3553 41739 3587
rect 41739 3553 41748 3587
rect 41696 3544 41748 3553
rect 42340 3587 42392 3596
rect 42340 3553 42349 3587
rect 42349 3553 42383 3587
rect 42383 3553 42392 3587
rect 42340 3544 42392 3553
rect 42984 3587 43036 3596
rect 42984 3553 42993 3587
rect 42993 3553 43027 3587
rect 43027 3553 43036 3587
rect 42984 3544 43036 3553
rect 44824 3587 44876 3596
rect 42248 3476 42300 3528
rect 44824 3553 44833 3587
rect 44833 3553 44867 3587
rect 44867 3553 44876 3587
rect 44824 3544 44876 3553
rect 46572 3544 46624 3596
rect 47308 3544 47360 3596
rect 47952 3544 48004 3596
rect 48412 3476 48464 3528
rect 49784 3587 49836 3596
rect 49784 3553 49793 3587
rect 49793 3553 49827 3587
rect 49827 3553 49836 3587
rect 49784 3544 49836 3553
rect 50896 3544 50948 3596
rect 52092 3587 52144 3596
rect 52092 3553 52101 3587
rect 52101 3553 52135 3587
rect 52135 3553 52144 3587
rect 52092 3544 52144 3553
rect 52736 3587 52788 3596
rect 52736 3553 52745 3587
rect 52745 3553 52779 3587
rect 52779 3553 52788 3587
rect 52736 3544 52788 3553
rect 53288 3544 53340 3596
rect 53932 3544 53984 3596
rect 54576 3544 54628 3596
rect 55128 3544 55180 3596
rect 56324 3544 56376 3596
rect 57152 3544 57204 3596
rect 58164 3587 58216 3596
rect 58164 3553 58173 3587
rect 58173 3553 58207 3587
rect 58207 3553 58216 3587
rect 58164 3544 58216 3553
rect 58808 3587 58860 3596
rect 58808 3553 58817 3587
rect 58817 3553 58851 3587
rect 58851 3553 58860 3587
rect 58808 3544 58860 3553
rect 60648 3587 60700 3596
rect 57980 3476 58032 3528
rect 60648 3553 60657 3587
rect 60657 3553 60691 3587
rect 60691 3553 60700 3587
rect 60648 3544 60700 3553
rect 61292 3544 61344 3596
rect 64052 3612 64104 3664
rect 61844 3476 61896 3528
rect 63040 3476 63092 3528
rect 63684 3476 63736 3528
rect 64880 3544 64932 3596
rect 71320 3612 71372 3664
rect 78588 3612 78640 3664
rect 66720 3544 66772 3596
rect 67916 3587 67968 3596
rect 67916 3553 67925 3587
rect 67925 3553 67959 3587
rect 67959 3553 67968 3587
rect 67916 3544 67968 3553
rect 68560 3587 68612 3596
rect 68560 3553 68569 3587
rect 68569 3553 68603 3587
rect 68603 3553 68612 3587
rect 68560 3544 68612 3553
rect 69204 3587 69256 3596
rect 69204 3553 69213 3587
rect 69213 3553 69247 3587
rect 69247 3553 69256 3587
rect 69204 3544 69256 3553
rect 69756 3544 69808 3596
rect 70400 3544 70452 3596
rect 71044 3544 71096 3596
rect 71596 3544 71648 3596
rect 72792 3544 72844 3596
rect 74080 3587 74132 3596
rect 74080 3553 74089 3587
rect 74089 3553 74123 3587
rect 74123 3553 74132 3587
rect 74080 3544 74132 3553
rect 74632 3544 74684 3596
rect 75920 3587 75972 3596
rect 75920 3553 75929 3587
rect 75929 3553 75963 3587
rect 75963 3553 75972 3587
rect 75920 3544 75972 3553
rect 76472 3544 76524 3596
rect 77668 3544 77720 3596
rect 65524 3476 65576 3528
rect 74908 3476 74960 3528
rect 80244 3612 80296 3664
rect 82360 3680 82412 3732
rect 83556 3680 83608 3732
rect 87880 3680 87932 3732
rect 88800 3680 88852 3732
rect 89352 3680 89404 3732
rect 88708 3612 88760 3664
rect 43076 3408 43128 3460
rect 21824 3340 21876 3392
rect 23940 3340 23992 3392
rect 26240 3340 26292 3392
rect 26700 3340 26752 3392
rect 32404 3340 32456 3392
rect 32864 3340 32916 3392
rect 35808 3340 35860 3392
rect 38936 3340 38988 3392
rect 54024 3340 54076 3392
rect 55772 3408 55824 3460
rect 79600 3544 79652 3596
rect 80152 3544 80204 3596
rect 83004 3587 83056 3596
rect 83004 3553 83013 3587
rect 83013 3553 83047 3587
rect 83047 3553 83056 3587
rect 83004 3544 83056 3553
rect 83832 3544 83884 3596
rect 84384 3544 84436 3596
rect 85028 3544 85080 3596
rect 86224 3587 86276 3596
rect 86224 3553 86233 3587
rect 86233 3553 86267 3587
rect 86267 3553 86276 3587
rect 86224 3544 86276 3553
rect 86868 3587 86920 3596
rect 86868 3553 86877 3587
rect 86877 3553 86911 3587
rect 86911 3553 86920 3587
rect 86868 3544 86920 3553
rect 87512 3544 87564 3596
rect 89904 3612 89956 3664
rect 91744 3612 91796 3664
rect 88064 3476 88116 3528
rect 56876 3340 56928 3392
rect 61660 3340 61712 3392
rect 62028 3340 62080 3392
rect 62856 3340 62908 3392
rect 63224 3340 63276 3392
rect 74540 3340 74592 3392
rect 79140 3451 79192 3460
rect 79140 3417 79149 3451
rect 79149 3417 79183 3451
rect 79183 3417 79192 3451
rect 79140 3408 79192 3417
rect 81532 3451 81584 3460
rect 81532 3417 81541 3451
rect 81541 3417 81575 3451
rect 81575 3417 81584 3451
rect 81532 3408 81584 3417
rect 83740 3408 83792 3460
rect 89260 3408 89312 3460
rect 90548 3476 90600 3528
rect 91100 3476 91152 3528
rect 93032 3476 93084 3528
rect 95056 3544 95108 3596
rect 96804 3655 96856 3664
rect 96804 3621 96813 3655
rect 96813 3621 96847 3655
rect 96847 3621 96856 3655
rect 96804 3612 96856 3621
rect 94780 3476 94832 3528
rect 96160 3476 96212 3528
rect 99472 3476 99524 3528
rect 94964 3451 95016 3460
rect 94964 3417 94973 3451
rect 94973 3417 95007 3451
rect 95007 3417 95016 3451
rect 94964 3408 95016 3417
rect 98644 3408 98696 3460
rect 78036 3340 78088 3392
rect 97448 3340 97500 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 65686 3238 65738 3290
rect 65750 3238 65802 3290
rect 65814 3238 65866 3290
rect 65878 3238 65930 3290
rect 96406 3238 96458 3290
rect 96470 3238 96522 3290
rect 96534 3238 96586 3290
rect 96598 3238 96650 3290
rect 5172 3136 5224 3188
rect 5448 3136 5500 3188
rect 9680 3136 9732 3188
rect 13268 3136 13320 3188
rect 14372 3179 14424 3188
rect 5080 3111 5132 3120
rect 5080 3077 5089 3111
rect 5089 3077 5123 3111
rect 5123 3077 5132 3111
rect 5080 3068 5132 3077
rect 2136 3043 2188 3052
rect 2136 3009 2145 3043
rect 2145 3009 2179 3043
rect 2179 3009 2188 3043
rect 2136 3000 2188 3009
rect 3792 3000 3844 3052
rect 4160 3000 4212 3052
rect 4896 3000 4948 3052
rect 8208 3068 8260 3120
rect 10324 3068 10376 3120
rect 1492 2932 1544 2984
rect 2320 2932 2372 2984
rect 2872 2932 2924 2984
rect 7472 3000 7524 3052
rect 7564 3000 7616 3052
rect 9128 3000 9180 3052
rect 11796 3000 11848 3052
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 6000 2932 6052 2984
rect 7932 2932 7984 2984
rect 10232 2932 10284 2984
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 13268 2975 13320 2984
rect 13268 2941 13277 2975
rect 13277 2941 13311 2975
rect 13311 2941 13320 2975
rect 13268 2932 13320 2941
rect 4620 2864 4672 2916
rect 6368 2864 6420 2916
rect 9036 2864 9088 2916
rect 12348 2907 12400 2916
rect 12348 2873 12357 2907
rect 12357 2873 12391 2907
rect 12391 2873 12400 2907
rect 12348 2864 12400 2873
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 14464 3136 14516 3188
rect 15936 3179 15988 3188
rect 14188 3068 14240 3120
rect 15016 3068 15068 3120
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 16672 3136 16724 3188
rect 20168 3136 20220 3188
rect 20444 3136 20496 3188
rect 20904 3136 20956 3188
rect 21640 3136 21692 3188
rect 21824 3136 21876 3188
rect 19064 3068 19116 3120
rect 19156 3068 19208 3120
rect 35808 3136 35860 3188
rect 38016 3136 38068 3188
rect 38200 3136 38252 3188
rect 39488 3136 39540 3188
rect 39580 3136 39632 3188
rect 74540 3136 74592 3188
rect 74816 3179 74868 3188
rect 74816 3145 74825 3179
rect 74825 3145 74859 3179
rect 74859 3145 74868 3179
rect 74816 3136 74868 3145
rect 76380 3179 76432 3188
rect 76380 3145 76389 3179
rect 76389 3145 76423 3179
rect 76423 3145 76432 3179
rect 76380 3136 76432 3145
rect 78496 3179 78548 3188
rect 78496 3145 78505 3179
rect 78505 3145 78539 3179
rect 78539 3145 78548 3179
rect 78496 3136 78548 3145
rect 78588 3136 78640 3188
rect 80888 3136 80940 3188
rect 65524 3068 65576 3120
rect 66812 3111 66864 3120
rect 66812 3077 66821 3111
rect 66821 3077 66855 3111
rect 66855 3077 66864 3111
rect 66812 3068 66864 3077
rect 69296 3068 69348 3120
rect 70032 3068 70084 3120
rect 13912 2932 13964 2984
rect 15016 2975 15068 2984
rect 15016 2941 15025 2975
rect 15025 2941 15059 2975
rect 15059 2941 15068 2975
rect 15016 2932 15068 2941
rect 17408 3000 17460 3052
rect 18512 3000 18564 3052
rect 34704 3000 34756 3052
rect 35532 3043 35584 3052
rect 35532 3009 35541 3043
rect 35541 3009 35575 3043
rect 35575 3009 35584 3043
rect 35532 3000 35584 3009
rect 15752 2975 15804 2984
rect 15752 2941 15761 2975
rect 15761 2941 15795 2975
rect 15795 2941 15804 2975
rect 15752 2932 15804 2941
rect 16948 2932 17000 2984
rect 18144 2932 18196 2984
rect 18788 2932 18840 2984
rect 19340 2932 19392 2984
rect 20168 2932 20220 2984
rect 22100 2932 22152 2984
rect 22192 2932 22244 2984
rect 23480 2932 23532 2984
rect 25136 2932 25188 2984
rect 25596 2975 25648 2984
rect 25596 2941 25605 2975
rect 25605 2941 25639 2975
rect 25639 2941 25648 2975
rect 25596 2932 25648 2941
rect 2504 2796 2556 2848
rect 3424 2796 3476 2848
rect 9312 2796 9364 2848
rect 13452 2796 13504 2848
rect 18052 2864 18104 2916
rect 18696 2864 18748 2916
rect 20444 2864 20496 2916
rect 20628 2864 20680 2916
rect 19984 2796 20036 2848
rect 20076 2796 20128 2848
rect 21364 2796 21416 2848
rect 24860 2864 24912 2916
rect 26976 2932 27028 2984
rect 27620 2975 27672 2984
rect 27620 2941 27629 2975
rect 27629 2941 27663 2975
rect 27663 2941 27672 2975
rect 27620 2932 27672 2941
rect 28816 2932 28868 2984
rect 26240 2864 26292 2916
rect 27344 2864 27396 2916
rect 28448 2864 28500 2916
rect 29552 2932 29604 2984
rect 30104 2932 30156 2984
rect 30748 2932 30800 2984
rect 31392 2932 31444 2984
rect 32588 2932 32640 2984
rect 33232 2932 33284 2984
rect 33784 2932 33836 2984
rect 35348 2975 35400 2984
rect 35348 2941 35357 2975
rect 35357 2941 35391 2975
rect 35391 2941 35400 2975
rect 35348 2932 35400 2941
rect 42156 3000 42208 3052
rect 42432 3000 42484 3052
rect 34612 2864 34664 2916
rect 36176 2864 36228 2916
rect 36268 2864 36320 2916
rect 37464 2932 37516 2984
rect 39488 2932 39540 2984
rect 41144 2932 41196 2984
rect 43536 2932 43588 2984
rect 45744 2975 45796 2984
rect 37648 2864 37700 2916
rect 25228 2796 25280 2848
rect 25504 2796 25556 2848
rect 26148 2796 26200 2848
rect 35532 2796 35584 2848
rect 35716 2796 35768 2848
rect 35808 2796 35860 2848
rect 38016 2796 38068 2848
rect 41604 2864 41656 2916
rect 43628 2907 43680 2916
rect 43628 2873 43637 2907
rect 43637 2873 43671 2907
rect 43671 2873 43680 2907
rect 43628 2864 43680 2873
rect 44180 2864 44232 2916
rect 45744 2941 45753 2975
rect 45753 2941 45787 2975
rect 45787 2941 45796 2975
rect 45744 2932 45796 2941
rect 45560 2907 45612 2916
rect 45560 2873 45569 2907
rect 45569 2873 45603 2907
rect 45603 2873 45612 2907
rect 45560 2864 45612 2873
rect 46204 2932 46256 2984
rect 46848 2932 46900 2984
rect 49056 3000 49108 3052
rect 48136 2932 48188 2984
rect 49148 2932 49200 2984
rect 49792 2932 49844 2984
rect 50804 3000 50856 3052
rect 50988 3000 51040 3052
rect 55220 3043 55272 3052
rect 55220 3009 55229 3043
rect 55229 3009 55263 3043
rect 55263 3009 55272 3043
rect 55220 3000 55272 3009
rect 40132 2796 40184 2848
rect 41236 2796 41288 2848
rect 43168 2796 43220 2848
rect 44364 2796 44416 2848
rect 46112 2796 46164 2848
rect 46204 2796 46256 2848
rect 48044 2796 48096 2848
rect 49240 2864 49292 2916
rect 50160 2864 50212 2916
rect 51356 2864 51408 2916
rect 51448 2864 51500 2916
rect 54024 2932 54076 2984
rect 55312 2907 55364 2916
rect 55312 2873 55321 2907
rect 55321 2873 55355 2907
rect 55355 2873 55364 2907
rect 55312 2864 55364 2873
rect 49608 2796 49660 2848
rect 49792 2796 49844 2848
rect 49976 2796 50028 2848
rect 51080 2796 51132 2848
rect 53564 2796 53616 2848
rect 54760 2796 54812 2848
rect 58348 3000 58400 3052
rect 60832 3000 60884 3052
rect 64420 3000 64472 3052
rect 56692 2975 56744 2984
rect 56692 2941 56701 2975
rect 56701 2941 56735 2975
rect 56735 2941 56744 2975
rect 56692 2932 56744 2941
rect 55772 2864 55824 2916
rect 57612 2932 57664 2984
rect 59360 2975 59412 2984
rect 59360 2941 59369 2975
rect 59369 2941 59403 2975
rect 59403 2941 59412 2975
rect 59360 2932 59412 2941
rect 59452 2932 59504 2984
rect 60096 2932 60148 2984
rect 60924 2932 60976 2984
rect 62120 2932 62172 2984
rect 62764 2975 62816 2984
rect 62764 2941 62773 2975
rect 62773 2941 62807 2975
rect 62807 2941 62816 2975
rect 62764 2932 62816 2941
rect 63592 2975 63644 2984
rect 63592 2941 63601 2975
rect 63601 2941 63635 2975
rect 63635 2941 63644 2975
rect 63592 2932 63644 2941
rect 64328 2932 64380 2984
rect 65524 2932 65576 2984
rect 67272 3000 67324 3052
rect 57796 2864 57848 2916
rect 60280 2864 60332 2916
rect 61568 2907 61620 2916
rect 61568 2873 61577 2907
rect 61577 2873 61611 2907
rect 61611 2873 61620 2907
rect 61568 2864 61620 2873
rect 64512 2907 64564 2916
rect 64512 2873 64521 2907
rect 64521 2873 64555 2907
rect 64555 2873 64564 2907
rect 64512 2864 64564 2873
rect 64696 2907 64748 2916
rect 64696 2873 64705 2907
rect 64705 2873 64739 2907
rect 64739 2873 64748 2907
rect 64696 2864 64748 2873
rect 66904 2907 66956 2916
rect 66904 2873 66913 2907
rect 66913 2873 66947 2907
rect 66947 2873 66956 2907
rect 66904 2864 66956 2873
rect 56600 2796 56652 2848
rect 58992 2796 59044 2848
rect 61476 2796 61528 2848
rect 62672 2796 62724 2848
rect 66168 2796 66220 2848
rect 70124 3000 70176 3052
rect 71320 2975 71372 2984
rect 67364 2864 67416 2916
rect 71320 2941 71329 2975
rect 71329 2941 71363 2975
rect 71363 2941 71372 2975
rect 71320 2932 71372 2941
rect 71504 2975 71556 2984
rect 71504 2941 71512 2975
rect 71512 2941 71546 2975
rect 71546 2941 71556 2975
rect 71504 2932 71556 2941
rect 69388 2864 69440 2916
rect 70584 2907 70636 2916
rect 70584 2873 70593 2907
rect 70593 2873 70627 2907
rect 70627 2873 70636 2907
rect 70584 2864 70636 2873
rect 70860 2864 70912 2916
rect 74908 3000 74960 3052
rect 81808 3136 81860 3188
rect 82912 3136 82964 3188
rect 83464 3136 83516 3188
rect 85948 3136 86000 3188
rect 88340 3136 88392 3188
rect 89996 3136 90048 3188
rect 94412 3179 94464 3188
rect 94412 3145 94421 3179
rect 94421 3145 94455 3179
rect 94455 3145 94464 3179
rect 94412 3136 94464 3145
rect 95792 3179 95844 3188
rect 95792 3145 95801 3179
rect 95801 3145 95835 3179
rect 95835 3145 95844 3179
rect 95792 3136 95844 3145
rect 96068 3136 96120 3188
rect 92204 3068 92256 3120
rect 92940 3068 92992 3120
rect 71872 2975 71924 2984
rect 71872 2941 71881 2975
rect 71881 2941 71915 2975
rect 71915 2941 71924 2975
rect 71872 2932 71924 2941
rect 72240 2932 72292 2984
rect 73436 2932 73488 2984
rect 74816 2932 74868 2984
rect 75276 2932 75328 2984
rect 74908 2864 74960 2916
rect 76656 2907 76708 2916
rect 76656 2873 76665 2907
rect 76665 2873 76699 2907
rect 76699 2873 76708 2907
rect 76656 2864 76708 2873
rect 77576 2932 77628 2984
rect 78496 2932 78548 2984
rect 80888 2932 80940 2984
rect 82636 2932 82688 2984
rect 83280 2932 83332 2984
rect 85672 2932 85724 2984
rect 87604 2932 87656 2984
rect 87972 2975 88024 2984
rect 87972 2941 87981 2975
rect 87981 2941 88015 2975
rect 88015 2941 88024 2975
rect 87972 2932 88024 2941
rect 91560 2975 91612 2984
rect 91560 2941 91569 2975
rect 91569 2941 91603 2975
rect 91603 2941 91612 2975
rect 91560 2932 91612 2941
rect 92296 2975 92348 2984
rect 92296 2941 92305 2975
rect 92305 2941 92339 2975
rect 92339 2941 92348 2975
rect 92296 2932 92348 2941
rect 93952 2975 94004 2984
rect 93952 2941 93961 2975
rect 93961 2941 93995 2975
rect 93995 2941 94004 2975
rect 93952 2932 94004 2941
rect 79784 2864 79836 2916
rect 80336 2864 80388 2916
rect 85856 2907 85908 2916
rect 68192 2796 68244 2848
rect 69296 2796 69348 2848
rect 71964 2839 72016 2848
rect 71964 2805 71973 2839
rect 71973 2805 72007 2839
rect 72007 2805 72016 2839
rect 71964 2796 72016 2805
rect 72424 2796 72476 2848
rect 77944 2796 77996 2848
rect 85856 2873 85865 2907
rect 85865 2873 85899 2907
rect 85899 2873 85908 2907
rect 85856 2864 85908 2873
rect 85948 2864 86000 2916
rect 90088 2864 90140 2916
rect 93124 2907 93176 2916
rect 93124 2873 93133 2907
rect 93133 2873 93167 2907
rect 93167 2873 93176 2907
rect 93124 2864 93176 2873
rect 82176 2796 82228 2848
rect 87052 2796 87104 2848
rect 88800 2796 88852 2848
rect 90824 2796 90876 2848
rect 91928 2796 91980 2848
rect 92848 2796 92900 2848
rect 93400 2864 93452 2916
rect 93860 2864 93912 2916
rect 94412 2932 94464 2984
rect 96160 3000 96212 3052
rect 95792 2932 95844 2984
rect 93768 2796 93820 2848
rect 94596 2796 94648 2848
rect 95332 2796 95384 2848
rect 95608 2864 95660 2916
rect 96804 2932 96856 2984
rect 97724 3000 97776 3052
rect 98828 3000 98880 3052
rect 96896 2907 96948 2916
rect 96896 2873 96905 2907
rect 96905 2873 96939 2907
rect 96939 2873 96948 2907
rect 96896 2864 96948 2873
rect 98368 2864 98420 2916
rect 97724 2796 97776 2848
rect 99840 2796 99892 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 50326 2694 50378 2746
rect 50390 2694 50442 2746
rect 50454 2694 50506 2746
rect 50518 2694 50570 2746
rect 81046 2694 81098 2746
rect 81110 2694 81162 2746
rect 81174 2694 81226 2746
rect 81238 2694 81290 2746
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 13176 2592 13228 2644
rect 7656 2524 7708 2576
rect 10140 2567 10192 2576
rect 10140 2533 10149 2567
rect 10149 2533 10183 2567
rect 10183 2533 10192 2567
rect 10140 2524 10192 2533
rect 13360 2524 13412 2576
rect 15844 2592 15896 2644
rect 17776 2524 17828 2576
rect 18880 2524 18932 2576
rect 20536 2567 20588 2576
rect 20536 2533 20545 2567
rect 20545 2533 20579 2567
rect 20579 2533 20588 2567
rect 20536 2524 20588 2533
rect 21732 2524 21784 2576
rect 23112 2567 23164 2576
rect 23112 2533 23121 2567
rect 23121 2533 23155 2567
rect 23155 2533 23164 2567
rect 23112 2524 23164 2533
rect 23756 2567 23808 2576
rect 23756 2533 23765 2567
rect 23765 2533 23799 2567
rect 23799 2533 23808 2567
rect 23756 2524 23808 2533
rect 296 2456 348 2508
rect 3700 2456 3752 2508
rect 5172 2456 5224 2508
rect 5724 2456 5776 2508
rect 8392 2456 8444 2508
rect 9588 2456 9640 2508
rect 10876 2499 10928 2508
rect 10876 2465 10885 2499
rect 10885 2465 10919 2499
rect 10919 2465 10928 2499
rect 10876 2456 10928 2465
rect 11428 2456 11480 2508
rect 12624 2456 12676 2508
rect 14464 2456 14516 2508
rect 15108 2456 15160 2508
rect 16304 2456 16356 2508
rect 17684 2456 17736 2508
rect 19984 2456 20036 2508
rect 21180 2456 21232 2508
rect 26976 2524 27028 2576
rect 28448 2567 28500 2576
rect 28448 2533 28457 2567
rect 28457 2533 28491 2567
rect 28491 2533 28500 2567
rect 28448 2524 28500 2533
rect 28632 2592 28684 2644
rect 33140 2592 33192 2644
rect 33416 2592 33468 2644
rect 31024 2567 31076 2576
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 11520 2388 11572 2440
rect 16212 2388 16264 2440
rect 6092 2320 6144 2372
rect 21272 2320 21324 2372
rect 12164 2252 12216 2304
rect 13636 2252 13688 2304
rect 15568 2252 15620 2304
rect 25320 2456 25372 2508
rect 26240 2499 26292 2508
rect 26240 2465 26249 2499
rect 26249 2465 26283 2499
rect 26283 2465 26292 2499
rect 26240 2456 26292 2465
rect 27252 2499 27304 2508
rect 27252 2465 27261 2499
rect 27261 2465 27295 2499
rect 27295 2465 27304 2499
rect 27252 2456 27304 2465
rect 29736 2456 29788 2508
rect 31024 2533 31033 2567
rect 31033 2533 31067 2567
rect 31067 2533 31076 2567
rect 31024 2524 31076 2533
rect 32496 2567 32548 2576
rect 31760 2499 31812 2508
rect 23664 2388 23716 2440
rect 28172 2388 28224 2440
rect 31760 2465 31769 2499
rect 31769 2465 31803 2499
rect 31803 2465 31812 2499
rect 31760 2456 31812 2465
rect 32496 2533 32505 2567
rect 32505 2533 32539 2567
rect 32539 2533 32548 2567
rect 32496 2524 32548 2533
rect 33692 2567 33744 2576
rect 33692 2533 33701 2567
rect 33701 2533 33735 2567
rect 33735 2533 33744 2567
rect 33692 2524 33744 2533
rect 34060 2524 34112 2576
rect 35256 2524 35308 2576
rect 35992 2524 36044 2576
rect 36176 2524 36228 2576
rect 38292 2592 38344 2644
rect 36452 2499 36504 2508
rect 30932 2388 30984 2440
rect 36452 2465 36461 2499
rect 36461 2465 36495 2499
rect 36495 2465 36504 2499
rect 36452 2456 36504 2465
rect 36912 2499 36964 2508
rect 36912 2465 36921 2499
rect 36921 2465 36955 2499
rect 36955 2465 36964 2499
rect 36912 2456 36964 2465
rect 38752 2524 38804 2576
rect 39120 2567 39172 2576
rect 39120 2533 39129 2567
rect 39129 2533 39163 2567
rect 39163 2533 39172 2567
rect 39120 2524 39172 2533
rect 39856 2567 39908 2576
rect 39856 2533 39865 2567
rect 39865 2533 39899 2567
rect 39899 2533 39908 2567
rect 39856 2524 39908 2533
rect 40592 2567 40644 2576
rect 40592 2533 40601 2567
rect 40601 2533 40635 2567
rect 40635 2533 40644 2567
rect 40592 2524 40644 2533
rect 44732 2592 44784 2644
rect 42432 2567 42484 2576
rect 39396 2456 39448 2508
rect 39488 2456 39540 2508
rect 42432 2533 42441 2567
rect 42441 2533 42475 2567
rect 42475 2533 42484 2567
rect 42432 2524 42484 2533
rect 44088 2524 44140 2576
rect 44456 2567 44508 2576
rect 44456 2533 44465 2567
rect 44465 2533 44499 2567
rect 44499 2533 44508 2567
rect 44456 2524 44508 2533
rect 46112 2592 46164 2644
rect 48320 2635 48372 2644
rect 48320 2601 48329 2635
rect 48329 2601 48363 2635
rect 48363 2601 48372 2635
rect 48320 2592 48372 2601
rect 46756 2524 46808 2576
rect 47768 2567 47820 2576
rect 47768 2533 47777 2567
rect 47777 2533 47811 2567
rect 47811 2533 47820 2567
rect 47768 2524 47820 2533
rect 49792 2592 49844 2644
rect 49976 2592 50028 2644
rect 54024 2592 54076 2644
rect 57336 2592 57388 2644
rect 42248 2456 42300 2508
rect 42524 2456 42576 2508
rect 47676 2456 47728 2508
rect 49884 2456 49936 2508
rect 51540 2524 51592 2576
rect 52368 2567 52420 2576
rect 52368 2533 52377 2567
rect 52377 2533 52411 2567
rect 52411 2533 52420 2567
rect 52368 2524 52420 2533
rect 53748 2524 53800 2576
rect 54116 2524 54168 2576
rect 55036 2567 55088 2576
rect 55036 2533 55045 2567
rect 55045 2533 55079 2567
rect 55079 2533 55088 2567
rect 55036 2524 55088 2533
rect 55404 2524 55456 2576
rect 37924 2388 37976 2440
rect 40684 2388 40736 2440
rect 45008 2388 45060 2440
rect 21824 2320 21876 2372
rect 23020 2320 23072 2372
rect 22468 2252 22520 2304
rect 24216 2252 24268 2304
rect 27896 2320 27948 2372
rect 29092 2320 29144 2372
rect 30380 2320 30432 2372
rect 32220 2320 32272 2372
rect 34704 2320 34756 2372
rect 37188 2320 37240 2372
rect 39028 2320 39080 2372
rect 28540 2252 28592 2304
rect 29736 2252 29788 2304
rect 31576 2252 31628 2304
rect 33968 2252 34020 2304
rect 36452 2252 36504 2304
rect 37096 2252 37148 2304
rect 43812 2320 43864 2372
rect 51632 2456 51684 2508
rect 52460 2456 52512 2508
rect 56140 2524 56192 2576
rect 60280 2592 60332 2644
rect 61384 2592 61436 2644
rect 62120 2592 62172 2644
rect 58348 2567 58400 2576
rect 58348 2533 58357 2567
rect 58357 2533 58391 2567
rect 58391 2533 58400 2567
rect 58348 2524 58400 2533
rect 59176 2567 59228 2576
rect 59176 2533 59185 2567
rect 59185 2533 59219 2567
rect 59219 2533 59228 2567
rect 59176 2524 59228 2533
rect 60464 2567 60516 2576
rect 60464 2533 60473 2567
rect 60473 2533 60507 2567
rect 60507 2533 60516 2567
rect 60464 2524 60516 2533
rect 60740 2524 60792 2576
rect 58072 2456 58124 2508
rect 61200 2499 61252 2508
rect 61200 2465 61209 2499
rect 61209 2465 61243 2499
rect 61243 2465 61252 2499
rect 61200 2456 61252 2465
rect 61384 2456 61436 2508
rect 63132 2567 63184 2576
rect 63132 2533 63141 2567
rect 63141 2533 63175 2567
rect 63175 2533 63184 2567
rect 63132 2524 63184 2533
rect 63776 2567 63828 2576
rect 63776 2533 63785 2567
rect 63785 2533 63819 2567
rect 63819 2533 63828 2567
rect 63776 2524 63828 2533
rect 63868 2524 63920 2576
rect 64420 2456 64472 2508
rect 65432 2524 65484 2576
rect 66628 2592 66680 2644
rect 66996 2635 67048 2644
rect 66996 2601 67005 2635
rect 67005 2601 67039 2635
rect 67039 2601 67048 2635
rect 68100 2635 68152 2644
rect 66996 2592 67048 2601
rect 68100 2601 68109 2635
rect 68109 2601 68143 2635
rect 68143 2601 68152 2635
rect 68836 2635 68888 2644
rect 68100 2592 68152 2601
rect 68836 2601 68845 2635
rect 68845 2601 68879 2635
rect 68879 2601 68888 2635
rect 68836 2592 68888 2601
rect 71688 2592 71740 2644
rect 74172 2635 74224 2644
rect 70308 2524 70360 2576
rect 71228 2524 71280 2576
rect 74172 2601 74181 2635
rect 74181 2601 74215 2635
rect 74215 2601 74224 2635
rect 74172 2592 74224 2601
rect 74724 2592 74776 2644
rect 79508 2635 79560 2644
rect 79508 2601 79517 2635
rect 79517 2601 79551 2635
rect 79551 2601 79560 2635
rect 80244 2635 80296 2644
rect 79508 2592 79560 2601
rect 69296 2456 69348 2508
rect 71780 2499 71832 2508
rect 71780 2465 71789 2499
rect 71789 2465 71823 2499
rect 71823 2465 71832 2499
rect 71780 2456 71832 2465
rect 71872 2456 71924 2508
rect 72148 2456 72200 2508
rect 75368 2524 75420 2576
rect 76104 2524 76156 2576
rect 77852 2567 77904 2576
rect 76380 2499 76432 2508
rect 76380 2465 76389 2499
rect 76389 2465 76423 2499
rect 76423 2465 76432 2499
rect 76380 2456 76432 2465
rect 76564 2456 76616 2508
rect 77852 2533 77861 2567
rect 77861 2533 77895 2567
rect 77895 2533 77904 2567
rect 77852 2524 77904 2533
rect 80244 2601 80253 2635
rect 80253 2601 80287 2635
rect 80287 2601 80296 2635
rect 85764 2635 85816 2644
rect 80244 2592 80296 2601
rect 85764 2601 85773 2635
rect 85773 2601 85807 2635
rect 85807 2601 85816 2635
rect 85764 2592 85816 2601
rect 86408 2592 86460 2644
rect 82452 2524 82504 2576
rect 83096 2524 83148 2576
rect 86960 2524 87012 2576
rect 87788 2567 87840 2576
rect 87788 2533 87797 2567
rect 87797 2533 87831 2567
rect 87831 2533 87840 2567
rect 87788 2524 87840 2533
rect 88892 2592 88944 2644
rect 90180 2635 90232 2644
rect 90180 2601 90189 2635
rect 90189 2601 90223 2635
rect 90223 2601 90232 2635
rect 90916 2635 90968 2644
rect 90180 2592 90232 2601
rect 90916 2601 90925 2635
rect 90925 2601 90959 2635
rect 90959 2601 90968 2635
rect 92112 2635 92164 2644
rect 90916 2592 90968 2601
rect 92112 2601 92121 2635
rect 92121 2601 92155 2635
rect 92155 2601 92164 2635
rect 92112 2592 92164 2601
rect 94504 2592 94556 2644
rect 94044 2524 94096 2576
rect 97724 2524 97776 2576
rect 50528 2388 50580 2440
rect 55956 2388 56008 2440
rect 63408 2388 63460 2440
rect 41972 2252 42024 2304
rect 45468 2252 45520 2304
rect 50436 2320 50488 2372
rect 54116 2320 54168 2372
rect 47400 2252 47452 2304
rect 51724 2252 51776 2304
rect 57152 2320 57204 2372
rect 60372 2320 60424 2372
rect 63316 2320 63368 2372
rect 66812 2320 66864 2372
rect 68468 2320 68520 2372
rect 58072 2252 58124 2304
rect 59636 2252 59688 2304
rect 60740 2252 60792 2304
rect 62028 2252 62080 2304
rect 63960 2252 64012 2304
rect 66260 2252 66312 2304
rect 69296 2252 69348 2304
rect 71688 2388 71740 2440
rect 75000 2388 75052 2440
rect 79232 2456 79284 2508
rect 84292 2456 84344 2508
rect 84660 2499 84712 2508
rect 84660 2465 84669 2499
rect 84669 2465 84703 2499
rect 84703 2465 84712 2499
rect 84660 2456 84712 2465
rect 85304 2456 85356 2508
rect 88616 2499 88668 2508
rect 88616 2465 88625 2499
rect 88625 2465 88659 2499
rect 88659 2465 88668 2499
rect 88616 2456 88668 2465
rect 88800 2456 88852 2508
rect 84752 2388 84804 2440
rect 88248 2388 88300 2440
rect 92664 2456 92716 2508
rect 91284 2388 91336 2440
rect 95792 2499 95844 2508
rect 95792 2465 95801 2499
rect 95801 2465 95835 2499
rect 95835 2465 95844 2499
rect 95792 2456 95844 2465
rect 93952 2388 94004 2440
rect 94228 2388 94280 2440
rect 94320 2388 94372 2440
rect 97540 2456 97592 2508
rect 72700 2320 72752 2372
rect 72884 2320 72936 2372
rect 72148 2252 72200 2304
rect 72516 2295 72568 2304
rect 72516 2261 72525 2295
rect 72525 2261 72559 2295
rect 72559 2261 72568 2295
rect 72516 2252 72568 2261
rect 73068 2252 73120 2304
rect 75460 2320 75512 2372
rect 82820 2363 82872 2372
rect 82820 2329 82829 2363
rect 82829 2329 82863 2363
rect 82863 2329 82872 2363
rect 82820 2320 82872 2329
rect 87696 2320 87748 2372
rect 78680 2295 78732 2304
rect 78680 2261 78689 2295
rect 78689 2261 78723 2295
rect 78723 2261 78732 2295
rect 78680 2252 78732 2261
rect 83372 2252 83424 2304
rect 84016 2252 84068 2304
rect 88340 2295 88392 2304
rect 88340 2261 88349 2295
rect 88349 2261 88383 2295
rect 88383 2261 88392 2295
rect 88340 2252 88392 2261
rect 88616 2252 88668 2304
rect 88892 2252 88944 2304
rect 92572 2320 92624 2372
rect 99656 2320 99708 2372
rect 93308 2252 93360 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 65686 2150 65738 2202
rect 65750 2150 65802 2202
rect 65814 2150 65866 2202
rect 65878 2150 65930 2202
rect 96406 2150 96458 2202
rect 96470 2150 96522 2202
rect 96534 2150 96586 2202
rect 96598 2150 96650 2202
rect 18420 2048 18472 2100
rect 31760 2048 31812 2100
rect 48688 2048 48740 2100
rect 51632 2048 51684 2100
rect 56416 2048 56468 2100
rect 61200 2048 61252 2100
rect 61752 2048 61804 2100
rect 62120 2048 62172 2100
rect 63960 2048 64012 2100
rect 67548 2048 67600 2100
rect 69296 2048 69348 2100
rect 70032 2048 70084 2100
rect 71688 2048 71740 2100
rect 76380 2048 76432 2100
rect 80428 2048 80480 2100
rect 81164 2048 81216 2100
rect 82728 2048 82780 2100
rect 89536 2048 89588 2100
rect 93308 2048 93360 2100
rect 2044 1980 2096 2032
rect 3976 1912 4028 1964
rect 4344 1912 4396 1964
rect 21272 1912 21324 1964
rect 26240 1912 26292 1964
rect 25320 1844 25372 1896
rect 27252 1980 27304 2032
rect 31300 1980 31352 2032
rect 31668 1980 31720 2032
rect 33048 1980 33100 2032
rect 26792 1912 26844 1964
rect 38568 1980 38620 2032
rect 54392 1980 54444 2032
rect 63408 1980 63460 2032
rect 68744 1980 68796 2032
rect 72516 1980 72568 2032
rect 72700 1980 72752 2032
rect 78680 1980 78732 2032
rect 47676 1912 47728 1964
rect 53840 1912 53892 1964
rect 71780 1912 71832 1964
rect 82268 1912 82320 1964
rect 33508 1844 33560 1896
rect 51908 1844 51960 1896
rect 52644 1844 52696 1896
rect 66352 1844 66404 1896
rect 76564 1844 76616 1896
rect 31484 1776 31536 1828
rect 18052 1708 18104 1760
rect 33324 1708 33376 1760
rect 35256 1436 35308 1488
rect 37188 1436 37240 1488
rect 58440 1436 58492 1488
rect 60372 1436 60424 1488
rect 65708 1436 65760 1488
rect 66260 1436 66312 1488
rect 66352 1436 66404 1488
rect 68468 1436 68520 1488
rect 74264 1436 74316 1488
rect 74724 1436 74776 1488
rect 32772 1368 32824 1420
rect 33968 1368 34020 1420
rect 34060 1368 34112 1420
rect 34704 1368 34756 1420
rect 36452 1368 36504 1420
rect 37924 1368 37976 1420
rect 48688 1368 48740 1420
rect 50528 1368 50580 1420
rect 52920 1368 52972 1420
rect 54024 1368 54076 1420
rect 60188 1368 60240 1420
rect 62028 1368 62080 1420
rect 65064 1368 65116 1420
rect 66812 1368 66864 1420
rect 71228 1368 71280 1420
rect 72884 1368 72936 1420
rect 73620 1368 73672 1420
rect 75000 1368 75052 1420
rect 77300 1368 77352 1420
rect 79232 1368 79284 1420
rect 16396 1300 16448 1352
rect 30288 1300 30340 1352
rect 31760 1300 31812 1352
rect 43628 1300 43680 1352
rect 48964 1300 49016 1352
rect 58072 1300 58124 1352
rect 59728 1300 59780 1352
rect 62396 1300 62448 1352
rect 91376 1300 91428 1352
rect 38568 1232 38620 1284
rect 43076 1232 43128 1284
rect 43260 1232 43312 1284
rect 25872 1164 25924 1216
rect 36728 1164 36780 1216
rect 65248 1232 65300 1284
rect 72148 1164 72200 1216
rect 58348 1096 58400 1148
rect 63592 1096 63644 1148
rect 95792 1096 95844 1148
rect 12348 1028 12400 1080
rect 58256 1028 58308 1080
rect 92664 1028 92716 1080
rect 26056 960 26108 1012
rect 70676 960 70728 1012
rect 9312 892 9364 944
rect 33876 892 33928 944
rect 44272 892 44324 944
rect 46664 892 46716 944
rect 89812 892 89864 944
rect 13636 824 13688 876
rect 53012 824 53064 876
rect 59268 824 59320 876
rect 88340 824 88392 876
rect 34520 756 34572 808
rect 73528 756 73580 808
rect 25596 688 25648 740
rect 62212 688 62264 740
rect 20444 620 20496 672
rect 2596 552 2648 604
rect 37740 552 37792 604
rect 38568 552 38620 604
rect 42248 620 42300 672
rect 78036 620 78088 672
rect 44916 552 44968 604
rect 50804 552 50856 604
rect 15660 484 15712 536
rect 38384 416 38436 468
rect 71504 552 71556 604
rect 54852 484 54904 536
rect 71320 484 71372 536
rect 49332 416 49384 468
rect 72332 416 72384 468
rect 6460 348 6512 400
rect 92480 348 92532 400
rect 25964 280 26016 332
rect 92848 280 92900 332
rect 5264 212 5316 264
rect 62396 212 62448 264
rect 20260 144 20312 196
rect 73712 144 73764 196
rect 16212 76 16264 128
rect 48780 76 48832 128
rect 87144 76 87196 128
rect 37556 8 37608 60
rect 38384 8 38436 60
rect 39764 8 39816 60
rect 70860 8 70912 60
<< metal2 >>
rect 386 39200 442 40000
rect 1214 39200 1270 40000
rect 2134 39200 2190 40000
rect 2962 39200 3018 40000
rect 3882 39200 3938 40000
rect 4710 39200 4766 40000
rect 5630 39200 5686 40000
rect 6458 39200 6514 40000
rect 7378 39200 7434 40000
rect 8206 39200 8262 40000
rect 9126 39200 9182 40000
rect 9954 39200 10010 40000
rect 10874 39200 10930 40000
rect 11702 39200 11758 40000
rect 12622 39200 12678 40000
rect 13542 39200 13598 40000
rect 13728 39228 13780 39234
rect 400 37398 428 39200
rect 1228 37482 1256 39200
rect 1228 37466 1440 37482
rect 1228 37460 1452 37466
rect 1228 37454 1400 37460
rect 1400 37402 1452 37408
rect 388 37392 440 37398
rect 388 37334 440 37340
rect 2148 36854 2176 39200
rect 2976 37330 3004 39200
rect 3332 37868 3384 37874
rect 3332 37810 3384 37816
rect 2964 37324 3016 37330
rect 2964 37266 3016 37272
rect 2320 37256 2372 37262
rect 2320 37198 2372 37204
rect 2136 36848 2188 36854
rect 2136 36790 2188 36796
rect 2332 36718 2360 37198
rect 3148 37120 3200 37126
rect 3148 37062 3200 37068
rect 2596 36916 2648 36922
rect 2596 36858 2648 36864
rect 2320 36712 2372 36718
rect 2320 36654 2372 36660
rect 2502 29608 2558 29617
rect 2502 29543 2504 29552
rect 2556 29543 2558 29552
rect 2504 29514 2556 29520
rect 2504 28144 2556 28150
rect 2504 28086 2556 28092
rect 1492 24744 1544 24750
rect 1492 24686 1544 24692
rect 1768 24744 1820 24750
rect 1768 24686 1820 24692
rect 2136 24744 2188 24750
rect 2136 24686 2188 24692
rect 1398 20088 1454 20097
rect 1398 20023 1454 20032
rect 1412 19922 1440 20023
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1124 17604 1176 17610
rect 1124 17546 1176 17552
rect 480 5024 532 5030
rect 480 4966 532 4972
rect 112 3528 164 3534
rect 112 3470 164 3476
rect 124 800 152 3470
rect 296 2508 348 2514
rect 296 2450 348 2456
rect 308 800 336 2450
rect 492 800 520 4966
rect 848 4684 900 4690
rect 848 4626 900 4632
rect 664 4004 716 4010
rect 664 3946 716 3952
rect 676 800 704 3946
rect 860 800 888 4626
rect 1136 3534 1164 17546
rect 1504 7954 1532 24686
rect 1780 23866 1808 24686
rect 1768 23860 1820 23866
rect 1768 23802 1820 23808
rect 1860 23316 1912 23322
rect 1860 23258 1912 23264
rect 1872 21146 1900 23258
rect 2044 22704 2096 22710
rect 2044 22646 2096 22652
rect 1860 21140 1912 21146
rect 1860 21082 1912 21088
rect 1952 18692 2004 18698
rect 1952 18634 2004 18640
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1504 7342 1532 7890
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1872 7546 1900 7822
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1216 4072 1268 4078
rect 1216 4014 1268 4020
rect 1124 3528 1176 3534
rect 1124 3470 1176 3476
rect 1228 2122 1256 4014
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 1136 2094 1256 2122
rect 1136 800 1164 2094
rect 1320 800 1348 3402
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1504 800 1532 2926
rect 1688 800 1716 4490
rect 1872 800 1900 5714
rect 1964 4826 1992 18634
rect 2056 17490 2084 22646
rect 2148 20618 2176 24686
rect 2320 23248 2372 23254
rect 2320 23190 2372 23196
rect 2148 20590 2268 20618
rect 2134 17776 2190 17785
rect 2134 17711 2190 17720
rect 2148 17678 2176 17711
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2056 17462 2176 17490
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 2056 7954 2084 17274
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1964 1850 1992 3538
rect 2056 2038 2084 5034
rect 2148 3058 2176 17462
rect 2240 11898 2268 20590
rect 2332 17338 2360 23190
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 2424 21010 2452 21490
rect 2412 21004 2464 21010
rect 2412 20946 2464 20952
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2424 17202 2452 17614
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2516 4826 2544 28086
rect 2608 17746 2636 36858
rect 3056 25424 3108 25430
rect 3056 25366 3108 25372
rect 3068 24750 3096 25366
rect 2872 24744 2924 24750
rect 2872 24686 2924 24692
rect 3056 24744 3108 24750
rect 3056 24686 3108 24692
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2700 23798 2728 24550
rect 2688 23792 2740 23798
rect 2688 23734 2740 23740
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2884 7954 2912 24686
rect 2964 24608 3016 24614
rect 2964 24550 3016 24556
rect 2976 20602 3004 24550
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2976 16658 3004 17682
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2964 15632 3016 15638
rect 2964 15574 3016 15580
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2688 7880 2740 7886
rect 2686 7848 2688 7857
rect 2740 7848 2742 7857
rect 2686 7783 2742 7792
rect 2884 7410 2912 7890
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2044 2032 2096 2038
rect 2044 1974 2096 1980
rect 1964 1822 2176 1850
rect 2148 800 2176 1822
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2240 785 2268 3946
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2332 800 2360 2926
rect 2226 776 2282 785
rect 2226 711 2282 720
rect 2318 0 2374 800
rect 2424 241 2452 3470
rect 2792 2938 2820 5714
rect 2976 4146 3004 15574
rect 3160 7002 3188 37062
rect 3238 36816 3294 36825
rect 3238 36751 3240 36760
rect 3292 36751 3294 36760
rect 3240 36722 3292 36728
rect 3240 24812 3292 24818
rect 3240 24754 3292 24760
rect 3252 20058 3280 24754
rect 3344 24750 3372 37810
rect 3896 37398 3924 39200
rect 4344 38140 4396 38146
rect 4344 38082 4396 38088
rect 3884 37392 3936 37398
rect 3884 37334 3936 37340
rect 4356 37330 4384 38082
rect 4724 37670 4752 39200
rect 5644 37890 5672 39200
rect 5460 37862 5672 37890
rect 4712 37664 4764 37670
rect 4712 37606 4764 37612
rect 5460 37330 5488 37862
rect 5724 37732 5776 37738
rect 5724 37674 5776 37680
rect 5736 37330 5764 37674
rect 6472 37466 6500 39200
rect 7012 37800 7064 37806
rect 7012 37742 7064 37748
rect 6460 37460 6512 37466
rect 6460 37402 6512 37408
rect 7024 37398 7052 37742
rect 7012 37392 7064 37398
rect 7012 37334 7064 37340
rect 4344 37324 4396 37330
rect 4344 37266 4396 37272
rect 5448 37324 5500 37330
rect 5448 37266 5500 37272
rect 5724 37324 5776 37330
rect 5724 37266 5776 37272
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 7392 36854 7420 39200
rect 7380 36848 7432 36854
rect 7380 36790 7432 36796
rect 8220 36718 8248 39200
rect 8392 37664 8444 37670
rect 8392 37606 8444 37612
rect 8484 37664 8536 37670
rect 8484 37606 8536 37612
rect 8404 37466 8432 37606
rect 8392 37460 8444 37466
rect 8392 37402 8444 37408
rect 8496 37398 8524 37606
rect 9140 37398 9168 39200
rect 8484 37392 8536 37398
rect 8484 37334 8536 37340
rect 9128 37392 9180 37398
rect 9128 37334 9180 37340
rect 9968 36854 9996 39200
rect 10784 38888 10836 38894
rect 10784 38830 10836 38836
rect 10416 38072 10468 38078
rect 10416 38014 10468 38020
rect 9956 36848 10008 36854
rect 9956 36790 10008 36796
rect 3516 36712 3568 36718
rect 3516 36654 3568 36660
rect 8208 36712 8260 36718
rect 8208 36654 8260 36660
rect 3424 31476 3476 31482
rect 3424 31418 3476 31424
rect 3332 24744 3384 24750
rect 3332 24686 3384 24692
rect 3436 20874 3464 31418
rect 3528 29102 3556 36654
rect 7472 36644 7524 36650
rect 7472 36586 7524 36592
rect 10324 36644 10376 36650
rect 10324 36586 10376 36592
rect 4896 36236 4948 36242
rect 4896 36178 4948 36184
rect 6184 36236 6236 36242
rect 6184 36178 6236 36184
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 3608 31680 3660 31686
rect 3608 31622 3660 31628
rect 3516 29096 3568 29102
rect 3516 29038 3568 29044
rect 3528 28626 3556 29038
rect 3516 28620 3568 28626
rect 3516 28562 3568 28568
rect 3620 28218 3648 31622
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4908 31210 4936 36178
rect 6196 31754 6224 36178
rect 6460 36032 6512 36038
rect 6460 35974 6512 35980
rect 6104 31726 6224 31754
rect 4896 31204 4948 31210
rect 4896 31146 4948 31152
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 3608 28212 3660 28218
rect 3608 28154 3660 28160
rect 3792 28212 3844 28218
rect 3792 28154 3844 28160
rect 3804 28014 3832 28154
rect 4080 28014 4108 28698
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 3792 28008 3844 28014
rect 3792 27950 3844 27956
rect 4068 28008 4120 28014
rect 4068 27950 4120 27956
rect 3976 27872 4028 27878
rect 3976 27814 4028 27820
rect 3988 27674 4016 27814
rect 3976 27668 4028 27674
rect 3976 27610 4028 27616
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4712 26444 4764 26450
rect 4712 26386 4764 26392
rect 4620 26308 4672 26314
rect 4620 26250 4672 26256
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 3700 24744 3752 24750
rect 3700 24686 3752 24692
rect 3712 24410 3740 24686
rect 3700 24404 3752 24410
rect 3700 24346 3752 24352
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 3424 20868 3476 20874
rect 3424 20810 3476 20816
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 3240 20052 3292 20058
rect 3240 19994 3292 20000
rect 3792 19984 3844 19990
rect 3792 19926 3844 19932
rect 3608 13456 3660 13462
rect 3608 13398 3660 13404
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 3436 9518 3464 12106
rect 3620 9518 3648 13398
rect 3240 9512 3292 9518
rect 3238 9480 3240 9489
rect 3424 9512 3476 9518
rect 3292 9480 3294 9489
rect 3424 9454 3476 9460
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3238 9415 3294 9424
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3712 8294 3740 9386
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3516 6248 3568 6254
rect 3054 6216 3110 6225
rect 3516 6190 3568 6196
rect 3054 6151 3110 6160
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3068 3670 3096 6151
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2700 2910 2820 2938
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2516 800 2544 2790
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2410 232 2466 241
rect 2410 167 2466 176
rect 2502 0 2558 800
rect 2608 610 2636 2382
rect 2700 800 2728 2910
rect 2884 800 2912 2926
rect 3160 800 3188 4014
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3344 800 3372 3946
rect 3436 2854 3464 4966
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3528 800 3556 6190
rect 3804 3058 3832 19926
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4632 6338 4660 26250
rect 4724 24886 4752 26386
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 4724 24426 4752 24822
rect 4724 24398 4844 24426
rect 4712 24268 4764 24274
rect 4712 24210 4764 24216
rect 4724 22982 4752 24210
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4724 6914 4752 22918
rect 4816 9042 4844 24398
rect 4908 21010 4936 31146
rect 6104 30258 6132 31726
rect 6092 30252 6144 30258
rect 6092 30194 6144 30200
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 6000 28416 6052 28422
rect 6000 28358 6052 28364
rect 5368 28150 5396 28358
rect 5356 28144 5408 28150
rect 5356 28086 5408 28092
rect 5356 26852 5408 26858
rect 5356 26794 5408 26800
rect 5368 26586 5396 26794
rect 5356 26580 5408 26586
rect 5356 26522 5408 26528
rect 5172 26444 5224 26450
rect 5172 26386 5224 26392
rect 5080 26376 5132 26382
rect 5080 26318 5132 26324
rect 5092 24682 5120 26318
rect 5080 24676 5132 24682
rect 5080 24618 5132 24624
rect 5184 22094 5212 26386
rect 5356 24676 5408 24682
rect 5356 24618 5408 24624
rect 5092 22066 5212 22094
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 5000 18222 5028 19246
rect 4988 18216 5040 18222
rect 4988 18158 5040 18164
rect 5092 13802 5120 22066
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10198 4936 10950
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 5092 9042 5120 13738
rect 5276 9450 5304 18566
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 4724 6886 5028 6914
rect 4632 6310 4844 6338
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3712 800 3740 2450
rect 3896 800 3924 3538
rect 3988 1970 4016 6190
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4172 2394 4200 2994
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4080 2366 4200 2394
rect 4080 1986 4108 2366
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 3976 1964 4028 1970
rect 4080 1958 4200 1986
rect 3976 1906 4028 1912
rect 4172 800 4200 1958
rect 4344 1964 4396 1970
rect 4344 1906 4396 1912
rect 4356 800 4384 1906
rect 4632 1442 4660 2858
rect 4540 1414 4660 1442
rect 4540 800 4568 1414
rect 4724 800 4752 4014
rect 4816 3670 4844 6310
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4908 3058 4936 4966
rect 5000 4162 5028 6886
rect 5080 5568 5132 5574
rect 5078 5536 5080 5545
rect 5132 5536 5134 5545
rect 5078 5471 5134 5480
rect 5184 4298 5212 8910
rect 5276 5166 5304 9386
rect 5368 9110 5396 24618
rect 5448 21616 5500 21622
rect 5448 21558 5500 21564
rect 5460 21010 5488 21558
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5540 20868 5592 20874
rect 5540 20810 5592 20816
rect 5552 20466 5580 20810
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5552 18426 5580 19178
rect 5644 18970 5672 20878
rect 5920 20874 5948 20946
rect 5908 20868 5960 20874
rect 5908 20810 5960 20816
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5460 10538 5488 14350
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 6322 5396 6734
rect 5446 6352 5502 6361
rect 5356 6316 5408 6322
rect 5446 6287 5502 6296
rect 5356 6258 5408 6264
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5184 4270 5304 4298
rect 5000 4134 5212 4162
rect 5276 4146 5304 4270
rect 5460 4162 5488 6287
rect 5080 3936 5132 3942
rect 5000 3896 5080 3924
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 5000 800 5028 3896
rect 5080 3878 5132 3884
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5092 3126 5120 3674
rect 5184 3194 5212 4134
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5368 4134 5488 4162
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5184 800 5212 2450
rect 2596 604 2648 610
rect 2596 546 2648 552
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5276 270 5304 3946
rect 5368 3738 5396 4134
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5368 800 5396 3538
rect 5460 3194 5488 4014
rect 5552 3670 5580 16050
rect 6012 12434 6040 28358
rect 6104 18358 6132 30194
rect 6472 29578 6500 35974
rect 6736 35012 6788 35018
rect 6736 34954 6788 34960
rect 6748 31754 6776 34954
rect 6748 31726 6868 31754
rect 6460 29572 6512 29578
rect 6460 29514 6512 29520
rect 6736 28620 6788 28626
rect 6736 28562 6788 28568
rect 6748 26450 6776 28562
rect 6736 26444 6788 26450
rect 6736 26386 6788 26392
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6196 21078 6224 21830
rect 6184 21072 6236 21078
rect 6184 21014 6236 21020
rect 6196 20942 6224 21014
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6276 20460 6328 20466
rect 6276 20402 6328 20408
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 6012 12406 6132 12434
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 5710 5672 6802
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5644 2774 5672 4966
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5552 2746 5672 2774
rect 5552 800 5580 2746
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5736 800 5764 2450
rect 6012 800 6040 2926
rect 6104 2378 6132 12406
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 6196 4622 6224 9930
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6092 2372 6144 2378
rect 6092 2314 6144 2320
rect 6196 800 6224 4082
rect 6288 3670 6316 20402
rect 6656 17542 6684 20742
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6748 16250 6776 19314
rect 6840 18902 6868 31726
rect 7288 27056 7340 27062
rect 7288 26998 7340 27004
rect 6920 23316 6972 23322
rect 6920 23258 6972 23264
rect 6932 23186 6960 23258
rect 6920 23180 6972 23186
rect 6920 23122 6972 23128
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6656 14006 6684 14214
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6748 11150 6776 14962
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6932 11150 6960 11630
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6460 6792 6512 6798
rect 6512 6752 6592 6780
rect 6460 6734 6512 6740
rect 6564 6662 6592 6752
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6368 2916 6420 2922
rect 6368 2858 6420 2864
rect 6380 800 6408 2858
rect 5264 264 5316 270
rect 5264 206 5316 212
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6472 406 6500 6598
rect 6564 6254 6592 6598
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6656 4758 6684 8298
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6564 800 6592 4014
rect 6748 800 6776 5102
rect 6932 2938 6960 5714
rect 7024 3942 7052 12378
rect 7208 6390 7236 15438
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7300 4758 7328 26998
rect 7484 15094 7512 36586
rect 8392 36576 8444 36582
rect 8392 36518 8444 36524
rect 8404 36378 8432 36518
rect 8300 36372 8352 36378
rect 8300 36314 8352 36320
rect 8392 36372 8444 36378
rect 8392 36314 8444 36320
rect 7564 34672 7616 34678
rect 7564 34614 7616 34620
rect 7576 23186 7604 34614
rect 8312 30394 8340 36314
rect 9956 34400 10008 34406
rect 9956 34342 10008 34348
rect 9968 34066 9996 34342
rect 9956 34060 10008 34066
rect 9956 34002 10008 34008
rect 9956 33924 10008 33930
rect 9956 33866 10008 33872
rect 8944 31340 8996 31346
rect 8944 31282 8996 31288
rect 8300 30388 8352 30394
rect 8300 30330 8352 30336
rect 7564 23180 7616 23186
rect 7564 23122 7616 23128
rect 8116 20868 8168 20874
rect 8116 20810 8168 20816
rect 7932 18352 7984 18358
rect 7932 18294 7984 18300
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7484 9042 7512 15030
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7380 4548 7432 4554
rect 7380 4490 7432 4496
rect 7116 4146 7144 4490
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 6932 2910 7052 2938
rect 7024 800 7052 2910
rect 7208 800 7236 3538
rect 7392 800 7420 4490
rect 7484 3058 7512 6666
rect 7576 5370 7604 11494
rect 7668 11150 7696 12718
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7668 9994 7696 11086
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7668 5778 7696 6054
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7654 5672 7710 5681
rect 7654 5607 7656 5616
rect 7708 5607 7710 5616
rect 7656 5578 7708 5584
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7760 4162 7788 6598
rect 7668 4134 7788 4162
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7576 800 7604 2994
rect 7668 2582 7696 4134
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7760 800 7788 4014
rect 7852 3942 7880 17002
rect 7944 12850 7972 18294
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7944 2990 7972 6122
rect 8036 3670 8064 17274
rect 8128 17066 8156 20810
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8128 4758 8156 15370
rect 8220 14414 8248 18770
rect 8576 18692 8628 18698
rect 8576 18634 8628 18640
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8312 18086 8340 18226
rect 8588 18154 8616 18634
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8220 12782 8248 14350
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8220 5642 8248 6326
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8404 5574 8432 6394
rect 8760 5704 8812 5710
rect 8758 5672 8760 5681
rect 8812 5672 8814 5681
rect 8758 5607 8814 5616
rect 8392 5568 8444 5574
rect 8484 5568 8536 5574
rect 8392 5510 8444 5516
rect 8482 5536 8484 5545
rect 8536 5536 8538 5545
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8220 4486 8248 4966
rect 8312 4622 8340 5102
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 8036 800 8064 3470
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8220 800 8248 3062
rect 8404 2650 8432 5510
rect 8482 5471 8538 5480
rect 8956 4826 8984 31282
rect 9312 31272 9364 31278
rect 9312 31214 9364 31220
rect 9324 30394 9352 31214
rect 9312 30388 9364 30394
rect 9312 30330 9364 30336
rect 9036 28960 9088 28966
rect 9036 28902 9088 28908
rect 9048 9110 9076 28902
rect 9128 24948 9180 24954
rect 9128 24890 9180 24896
rect 9140 10062 9168 24890
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 9232 8362 9260 23122
rect 9324 18290 9352 30330
rect 9404 29096 9456 29102
rect 9404 29038 9456 29044
rect 9416 23118 9444 29038
rect 9496 23860 9548 23866
rect 9496 23802 9548 23808
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9324 11626 9352 18226
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 6390 9168 7278
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8404 800 8432 2450
rect 8588 800 8616 3878
rect 8864 800 8892 4626
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 3534 8984 3878
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9140 3058 9168 5102
rect 9416 4078 9444 19858
rect 9508 8022 9536 23802
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9784 14822 9812 23054
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9876 16250 9904 22034
rect 9968 22001 9996 33866
rect 10140 30932 10192 30938
rect 10140 30874 10192 30880
rect 10152 30258 10180 30874
rect 10336 30394 10364 36586
rect 10324 30388 10376 30394
rect 10324 30330 10376 30336
rect 10140 30252 10192 30258
rect 10140 30194 10192 30200
rect 10336 26518 10364 30330
rect 10324 26512 10376 26518
rect 10324 26454 10376 26460
rect 9954 21992 10010 22001
rect 9954 21927 10010 21936
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9876 13870 9904 14894
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9784 10266 9812 13806
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 9508 7342 9536 7958
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 9048 800 9076 2858
rect 9232 800 9260 3334
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9324 950 9352 2790
rect 9508 2774 9536 4014
rect 9692 3194 9720 9862
rect 10046 7984 10102 7993
rect 10046 7919 10102 7928
rect 10060 7886 10088 7919
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 7342 10088 7686
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10152 6914 10180 19110
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10336 13938 10364 16662
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 12434 10272 13670
rect 10244 12406 10364 12434
rect 10336 11830 10364 12406
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10428 7954 10456 38014
rect 10796 37466 10824 38830
rect 10784 37460 10836 37466
rect 10784 37402 10836 37408
rect 10888 37346 10916 39200
rect 11060 37936 11112 37942
rect 11060 37878 11112 37884
rect 11072 37466 11100 37878
rect 11716 37466 11744 39200
rect 12348 37732 12400 37738
rect 12348 37674 12400 37680
rect 11060 37460 11112 37466
rect 11060 37402 11112 37408
rect 11704 37460 11756 37466
rect 11704 37402 11756 37408
rect 12360 37398 12388 37674
rect 11152 37392 11204 37398
rect 10888 37330 11008 37346
rect 11152 37334 11204 37340
rect 12348 37392 12400 37398
rect 12348 37334 12400 37340
rect 10888 37324 11020 37330
rect 10888 37318 10968 37324
rect 10968 37266 11020 37272
rect 10968 36168 11020 36174
rect 10968 36110 11020 36116
rect 10784 30252 10836 30258
rect 10784 30194 10836 30200
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10520 10062 10548 18294
rect 10612 16114 10640 24142
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10612 7886 10640 13874
rect 10796 12374 10824 30194
rect 10876 30184 10928 30190
rect 10876 30126 10928 30132
rect 10888 24206 10916 30126
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10874 18184 10930 18193
rect 10874 18119 10930 18128
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10888 12306 10916 18119
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10888 8090 10916 10202
rect 10980 9178 11008 36110
rect 11164 30802 11192 37334
rect 12636 36854 12664 39200
rect 13556 37330 13584 39200
rect 14370 39200 14426 40000
rect 15290 39200 15346 40000
rect 16118 39200 16174 40000
rect 17038 39200 17094 40000
rect 17866 39200 17922 40000
rect 18786 39200 18842 40000
rect 19614 39200 19670 40000
rect 20534 39200 20590 40000
rect 21362 39200 21418 40000
rect 21916 39296 21968 39302
rect 21916 39238 21968 39244
rect 13728 39170 13780 39176
rect 13544 37324 13596 37330
rect 13544 37266 13596 37272
rect 12624 36848 12676 36854
rect 12624 36790 12676 36796
rect 12992 36236 13044 36242
rect 12992 36178 13044 36184
rect 11888 35692 11940 35698
rect 11888 35634 11940 35640
rect 11612 32292 11664 32298
rect 11612 32234 11664 32240
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 11428 30796 11480 30802
rect 11428 30738 11480 30744
rect 11244 27532 11296 27538
rect 11244 27474 11296 27480
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 11164 24070 11192 27406
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 9968 6886 10180 6914
rect 9968 3670 9996 6886
rect 10980 6866 11008 9114
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10140 4072 10192 4078
rect 10060 4032 10140 4060
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9416 2746 9536 2774
rect 9312 944 9364 950
rect 9312 886 9364 892
rect 9416 800 9444 2746
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9600 800 9628 2450
rect 9876 800 9904 3334
rect 10060 800 10088 4032
rect 10140 4014 10192 4020
rect 10244 3890 10272 6190
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10152 3862 10272 3890
rect 10152 2582 10180 3862
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10336 3126 10364 3538
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 10244 800 10272 2926
rect 10520 2774 10548 3334
rect 10428 2746 10548 2774
rect 10428 800 10456 2746
rect 10612 800 10640 4626
rect 11072 2650 11100 20742
rect 11164 16998 11192 24006
rect 11256 22642 11284 27474
rect 11440 23254 11468 30738
rect 11520 27532 11572 27538
rect 11520 27474 11572 27480
rect 11532 26246 11560 27474
rect 11520 26240 11572 26246
rect 11520 26182 11572 26188
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 11428 22160 11480 22166
rect 11428 22102 11480 22108
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11164 10062 11192 14214
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10888 800 10916 2450
rect 11164 1442 11192 3674
rect 11072 1414 11192 1442
rect 11072 800 11100 1414
rect 11256 800 11284 4626
rect 11440 4078 11468 22102
rect 11624 22094 11652 32234
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11808 27606 11836 27950
rect 11796 27600 11848 27606
rect 11796 27542 11848 27548
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 11716 26042 11744 27474
rect 11704 26036 11756 26042
rect 11704 25978 11756 25984
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11532 22066 11652 22094
rect 11532 8906 11560 22066
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11624 9042 11652 16730
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11532 6322 11560 8842
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11624 6118 11652 8978
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11716 5930 11744 22578
rect 11794 9072 11850 9081
rect 11794 9007 11796 9016
rect 11848 9007 11850 9016
rect 11796 8978 11848 8984
rect 11532 5902 11744 5930
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11440 800 11468 2450
rect 11532 2446 11560 5902
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11716 5642 11744 5782
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11624 800 11652 3334
rect 11808 3058 11836 8978
rect 11900 7478 11928 35634
rect 13004 35562 13032 36178
rect 12992 35556 13044 35562
rect 12992 35498 13044 35504
rect 12164 35216 12216 35222
rect 12164 35158 12216 35164
rect 12072 30184 12124 30190
rect 12072 30126 12124 30132
rect 12084 30054 12112 30126
rect 12072 30048 12124 30054
rect 12072 29990 12124 29996
rect 12084 29102 12112 29990
rect 12072 29096 12124 29102
rect 12072 29038 12124 29044
rect 12176 21486 12204 35158
rect 13266 34640 13322 34649
rect 13266 34575 13322 34584
rect 12256 32428 12308 32434
rect 12256 32370 12308 32376
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 12084 19786 12112 21422
rect 12176 20806 12204 21422
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12072 19780 12124 19786
rect 12072 19722 12124 19728
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12176 9042 12204 18362
rect 12268 15162 12296 32370
rect 13280 31890 13308 34575
rect 13636 32768 13688 32774
rect 13636 32710 13688 32716
rect 13648 32570 13676 32710
rect 13636 32564 13688 32570
rect 13636 32506 13688 32512
rect 13740 32450 13768 39170
rect 13912 38752 13964 38758
rect 13912 38694 13964 38700
rect 13820 37800 13872 37806
rect 13820 37742 13872 37748
rect 13648 32422 13768 32450
rect 13084 31884 13136 31890
rect 13084 31826 13136 31832
rect 13268 31884 13320 31890
rect 13268 31826 13320 31832
rect 12440 31816 12492 31822
rect 12440 31758 12492 31764
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12452 12434 12480 31758
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12728 27130 12756 27270
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 12820 24818 12848 27474
rect 12992 27328 13044 27334
rect 12992 27270 13044 27276
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 12624 24404 12676 24410
rect 12624 24346 12676 24352
rect 12636 21486 12664 24346
rect 12728 22506 12756 24754
rect 13004 22574 13032 27270
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12716 22500 12768 22506
rect 12716 22442 12768 22448
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12820 20262 12848 21422
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 13096 14890 13124 31826
rect 13452 29776 13504 29782
rect 13452 29718 13504 29724
rect 13464 26314 13492 29718
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 13452 26308 13504 26314
rect 13452 26250 13504 26256
rect 13452 24744 13504 24750
rect 13452 24686 13504 24692
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 13372 23730 13400 24346
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13084 14884 13136 14890
rect 13084 14826 13136 14832
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 13096 14074 13124 14214
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12452 12406 12664 12434
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12544 11354 12572 11562
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12346 11248 12402 11257
rect 12346 11183 12348 11192
rect 12400 11183 12402 11192
rect 12532 11212 12584 11218
rect 12348 11154 12400 11160
rect 12532 11154 12584 11160
rect 12544 11121 12572 11154
rect 12530 11112 12586 11121
rect 12530 11047 12586 11056
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12452 10810 12480 10950
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 12268 9178 12296 10678
rect 12544 10470 12572 10950
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12636 9654 12664 12406
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12728 9518 12756 12718
rect 12912 11626 12940 13126
rect 13004 12782 13032 13262
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 13096 12714 13124 13194
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12806 11248 12862 11257
rect 12912 11218 12940 11562
rect 13082 11248 13138 11257
rect 12806 11183 12862 11192
rect 12900 11212 12952 11218
rect 12820 11150 12848 11183
rect 13082 11183 13084 11192
rect 12900 11154 12952 11160
rect 13136 11183 13138 11192
rect 13084 11154 13136 11160
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 12162 7440 12218 7449
rect 12162 7375 12218 7384
rect 11888 6180 11940 6186
rect 11888 6122 11940 6128
rect 11900 5846 11928 6122
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11900 800 11928 4626
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12084 800 12112 2926
rect 12176 2310 12204 7375
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12268 800 12296 3878
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 12360 1086 12388 2858
rect 12348 1080 12400 1086
rect 12348 1022 12400 1028
rect 12452 800 12480 4626
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13084 4004 13136 4010
rect 13084 3946 13136 3952
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12636 800 12664 2450
rect 12912 800 12940 3334
rect 13096 800 13124 3946
rect 13188 2650 13216 4014
rect 13280 3670 13308 13466
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 13280 3194 13308 3402
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13280 800 13308 2926
rect 13372 2582 13400 18022
rect 13464 3466 13492 24686
rect 13556 22166 13584 26522
rect 13544 22160 13596 22166
rect 13544 22102 13596 22108
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13556 18086 13584 18906
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13556 13530 13584 13942
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13648 9586 13676 32422
rect 13832 32366 13860 37742
rect 13924 37398 13952 38694
rect 14384 37398 14412 39200
rect 15108 38004 15160 38010
rect 15108 37946 15160 37952
rect 14924 37800 14976 37806
rect 14924 37742 14976 37748
rect 13912 37392 13964 37398
rect 13912 37334 13964 37340
rect 14372 37392 14424 37398
rect 14372 37334 14424 37340
rect 14096 36168 14148 36174
rect 14096 36110 14148 36116
rect 13912 36032 13964 36038
rect 13912 35974 13964 35980
rect 13820 32360 13872 32366
rect 13820 32302 13872 32308
rect 13728 31952 13780 31958
rect 13728 31894 13780 31900
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13740 7970 13768 31894
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13832 25265 13860 28086
rect 13924 27470 13952 35974
rect 14004 32836 14056 32842
rect 14004 32778 14056 32784
rect 14016 32502 14044 32778
rect 14004 32496 14056 32502
rect 14004 32438 14056 32444
rect 14004 32360 14056 32366
rect 14004 32302 14056 32308
rect 14016 30598 14044 32302
rect 14004 30592 14056 30598
rect 14004 30534 14056 30540
rect 14108 30410 14136 36110
rect 14464 35080 14516 35086
rect 14464 35022 14516 35028
rect 14188 30592 14240 30598
rect 14188 30534 14240 30540
rect 14016 30382 14136 30410
rect 14016 30258 14044 30382
rect 14200 30274 14228 30534
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 14108 30246 14228 30274
rect 14016 29102 14044 30194
rect 14004 29096 14056 29102
rect 14004 29038 14056 29044
rect 14004 27940 14056 27946
rect 14004 27882 14056 27888
rect 13912 27464 13964 27470
rect 13912 27406 13964 27412
rect 14016 26450 14044 27882
rect 14108 27878 14136 30246
rect 14280 28484 14332 28490
rect 14280 28426 14332 28432
rect 14292 28218 14320 28426
rect 14476 28218 14504 35022
rect 14936 31754 14964 37742
rect 15120 37398 15148 37946
rect 15108 37392 15160 37398
rect 15108 37334 15160 37340
rect 15304 36854 15332 39200
rect 15384 38208 15436 38214
rect 15384 38150 15436 38156
rect 15292 36848 15344 36854
rect 15292 36790 15344 36796
rect 15014 33960 15070 33969
rect 15014 33895 15070 33904
rect 14660 31726 14964 31754
rect 14556 29028 14608 29034
rect 14556 28970 14608 28976
rect 14660 28994 14688 31726
rect 14280 28212 14332 28218
rect 14280 28154 14332 28160
rect 14464 28212 14516 28218
rect 14464 28154 14516 28160
rect 14096 27872 14148 27878
rect 14096 27814 14148 27820
rect 14108 26994 14136 27814
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14188 27124 14240 27130
rect 14188 27066 14240 27072
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 14004 26444 14056 26450
rect 14004 26386 14056 26392
rect 13818 25256 13874 25265
rect 13818 25191 13874 25200
rect 14016 24954 14044 26386
rect 14004 24948 14056 24954
rect 14004 24890 14056 24896
rect 14200 23254 14228 27066
rect 14278 25256 14334 25265
rect 14278 25191 14334 25200
rect 14188 23248 14240 23254
rect 14188 23190 14240 23196
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13832 12646 13860 18702
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13648 7942 13768 7970
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 13556 3058 13584 6122
rect 13648 3602 13676 7942
rect 14200 6254 14228 23190
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14292 4842 14320 25191
rect 14200 4814 14320 4842
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 13464 800 13492 2790
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13648 882 13676 2246
rect 13636 876 13688 882
rect 13636 818 13688 824
rect 13740 800 13768 4014
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13924 800 13952 2926
rect 14108 800 14136 3334
rect 14200 3126 14228 4814
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14188 3120 14240 3126
rect 14188 3062 14240 3068
rect 14292 800 14320 4626
rect 14384 3194 14412 27406
rect 14568 21010 14596 28970
rect 14660 28966 14964 28994
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 14752 23186 14780 24550
rect 14936 23186 14964 28966
rect 14740 23180 14792 23186
rect 14740 23122 14792 23128
rect 14924 23180 14976 23186
rect 14924 23122 14976 23128
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14568 16182 14596 20946
rect 14752 20806 14780 23122
rect 15028 22778 15056 33895
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 15212 29510 15240 31826
rect 15396 31754 15424 38150
rect 15936 37664 15988 37670
rect 15936 37606 15988 37612
rect 15476 36712 15528 36718
rect 15476 36654 15528 36660
rect 15304 31726 15424 31754
rect 15488 31754 15516 36654
rect 15488 31726 15700 31754
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15108 28416 15160 28422
rect 15108 28358 15160 28364
rect 15120 28014 15148 28358
rect 15108 28008 15160 28014
rect 15108 27950 15160 27956
rect 15200 27600 15252 27606
rect 15200 27542 15252 27548
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 15120 25974 15148 26318
rect 15108 25968 15160 25974
rect 15108 25910 15160 25916
rect 15212 25498 15240 27542
rect 15200 25492 15252 25498
rect 15200 25434 15252 25440
rect 15212 25158 15240 25434
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15108 24336 15160 24342
rect 15108 24278 15160 24284
rect 15016 22772 15068 22778
rect 15016 22714 15068 22720
rect 15120 22710 15148 24278
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 15212 22710 15240 22986
rect 15108 22704 15160 22710
rect 15108 22646 15160 22652
rect 15200 22704 15252 22710
rect 15200 22646 15252 22652
rect 15108 22500 15160 22506
rect 15108 22442 15160 22448
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14752 9654 14780 20742
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15028 10062 15056 11494
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 15028 8974 15056 9998
rect 15120 9518 15148 22442
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15120 5778 15148 6054
rect 15212 5778 15240 6326
rect 15304 6254 15332 31726
rect 15476 30116 15528 30122
rect 15476 30058 15528 30064
rect 15488 29850 15516 30058
rect 15476 29844 15528 29850
rect 15476 29786 15528 29792
rect 15568 29096 15620 29102
rect 15568 29038 15620 29044
rect 15476 27396 15528 27402
rect 15476 27338 15528 27344
rect 15488 25702 15516 27338
rect 15476 25696 15528 25702
rect 15476 25638 15528 25644
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15396 6254 15424 25094
rect 15488 6322 15516 25638
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15488 5574 15516 6122
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14476 3194 14504 3402
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14476 800 14504 2450
rect 14752 800 14780 3402
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 15028 2990 15056 3062
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 15212 2774 15240 4626
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 14936 2746 15240 2774
rect 14936 800 14964 2746
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15120 800 15148 2450
rect 15304 800 15332 3878
rect 15488 800 15516 4014
rect 15580 2310 15608 29038
rect 15672 28801 15700 31726
rect 15844 30048 15896 30054
rect 15844 29990 15896 29996
rect 15856 29238 15884 29990
rect 15844 29232 15896 29238
rect 15844 29174 15896 29180
rect 15658 28792 15714 28801
rect 15658 28727 15714 28736
rect 15660 28620 15712 28626
rect 15856 28608 15884 29174
rect 15712 28580 15884 28608
rect 15660 28562 15712 28568
rect 15856 27470 15884 28580
rect 15844 27464 15896 27470
rect 15844 27406 15896 27412
rect 15856 26908 15884 27406
rect 15948 27130 15976 37606
rect 16132 37398 16160 39200
rect 16488 38412 16540 38418
rect 16488 38354 16540 38360
rect 16500 37466 16528 38354
rect 16856 38140 16908 38146
rect 16856 38082 16908 38088
rect 16868 38026 16896 38082
rect 16868 37998 16988 38026
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 16120 37392 16172 37398
rect 16120 37334 16172 37340
rect 16120 34604 16172 34610
rect 16120 34546 16172 34552
rect 16028 32292 16080 32298
rect 16028 32234 16080 32240
rect 16040 32026 16068 32234
rect 16028 32020 16080 32026
rect 16028 31962 16080 31968
rect 16026 28792 16082 28801
rect 16026 28727 16082 28736
rect 16040 27470 16068 28727
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 15856 26880 15976 26908
rect 15948 25974 15976 26880
rect 15936 25968 15988 25974
rect 15936 25910 15988 25916
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15672 22506 15700 23122
rect 15660 22500 15712 22506
rect 15660 22442 15712 22448
rect 15948 21010 15976 25910
rect 16132 22094 16160 34546
rect 16764 33108 16816 33114
rect 16764 33050 16816 33056
rect 16672 32972 16724 32978
rect 16672 32914 16724 32920
rect 16396 29844 16448 29850
rect 16396 29786 16448 29792
rect 16040 22066 16160 22094
rect 16408 22094 16436 29786
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16592 28150 16620 28494
rect 16580 28144 16632 28150
rect 16580 28086 16632 28092
rect 16488 24812 16540 24818
rect 16488 24754 16540 24760
rect 16500 22438 16528 24754
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16408 22066 16528 22094
rect 15936 21004 15988 21010
rect 15936 20946 15988 20952
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 6460 400 6512 406
rect 6460 342 6512 348
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 13910 0 13966 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15672 542 15700 8774
rect 15764 6390 15792 20878
rect 15844 20324 15896 20330
rect 15844 20266 15896 20272
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15752 2984 15804 2990
rect 15752 2926 15804 2932
rect 15764 800 15792 2926
rect 15856 2650 15884 20266
rect 16040 13190 16068 22066
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16316 18766 16344 21286
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16316 18034 16344 18702
rect 16132 18006 16344 18034
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16132 12434 16160 18006
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16316 15434 16344 17818
rect 16396 16516 16448 16522
rect 16396 16458 16448 16464
rect 16408 15502 16436 16458
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 15948 12406 16160 12434
rect 15948 3194 15976 12406
rect 16026 11112 16082 11121
rect 16026 11047 16082 11056
rect 16040 5370 16068 11047
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16040 3942 16068 5306
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 16040 1714 16068 3334
rect 15948 1686 16068 1714
rect 15948 800 15976 1686
rect 16132 800 16160 4626
rect 16224 3602 16252 8298
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 16304 2508 16356 2514
rect 16304 2450 16356 2456
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 15660 536 15712 542
rect 15660 478 15712 484
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16224 134 16252 2382
rect 16316 800 16344 2450
rect 16408 1358 16436 8978
rect 16500 8362 16528 22066
rect 16684 9178 16712 32914
rect 16776 31958 16804 33050
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 16764 31952 16816 31958
rect 16764 31894 16816 31900
rect 16868 31822 16896 32846
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 16856 31136 16908 31142
rect 16856 31078 16908 31084
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16776 28014 16804 28494
rect 16764 28008 16816 28014
rect 16764 27950 16816 27956
rect 16868 20534 16896 31078
rect 16960 30734 16988 37998
rect 17052 37466 17080 39200
rect 17500 38276 17552 38282
rect 17500 38218 17552 38224
rect 17040 37460 17092 37466
rect 17040 37402 17092 37408
rect 17408 36644 17460 36650
rect 17408 36586 17460 36592
rect 17316 32224 17368 32230
rect 17316 32166 17368 32172
rect 17040 31952 17092 31958
rect 17040 31894 17092 31900
rect 17052 31754 17080 31894
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 17040 31748 17092 31754
rect 17040 31690 17092 31696
rect 16948 30728 17000 30734
rect 16948 30670 17000 30676
rect 16960 24274 16988 30670
rect 17144 30598 17172 31758
rect 17224 31748 17276 31754
rect 17224 31690 17276 31696
rect 17132 30592 17184 30598
rect 17132 30534 17184 30540
rect 17132 30320 17184 30326
rect 17132 30262 17184 30268
rect 17144 29306 17172 30262
rect 17236 30190 17264 31690
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 17224 30048 17276 30054
rect 17224 29990 17276 29996
rect 17132 29300 17184 29306
rect 17132 29242 17184 29248
rect 17236 29170 17264 29990
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17040 28620 17092 28626
rect 17040 28562 17092 28568
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 17052 23186 17080 28562
rect 17224 28416 17276 28422
rect 17224 28358 17276 28364
rect 17132 28008 17184 28014
rect 17130 27976 17132 27985
rect 17184 27976 17186 27985
rect 17130 27911 17186 27920
rect 17236 25906 17264 28358
rect 17328 26926 17356 32166
rect 17420 28082 17448 36586
rect 17408 28076 17460 28082
rect 17408 28018 17460 28024
rect 17316 26920 17368 26926
rect 17316 26862 17368 26868
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 17144 24274 17172 24754
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 17236 22778 17264 23258
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17328 22642 17356 22986
rect 17316 22636 17368 22642
rect 17316 22578 17368 22584
rect 17316 22092 17368 22098
rect 17316 22034 17368 22040
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17144 21486 17172 21966
rect 17328 21622 17356 22034
rect 17420 21690 17448 28018
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17316 21616 17368 21622
rect 17512 21570 17540 38218
rect 17684 37732 17736 37738
rect 17684 37674 17736 37680
rect 17696 37398 17724 37674
rect 17684 37392 17736 37398
rect 17684 37334 17736 37340
rect 17880 36854 17908 39200
rect 18696 38480 18748 38486
rect 18696 38422 18748 38428
rect 17960 38140 18012 38146
rect 17960 38082 18012 38088
rect 17972 37466 18000 38082
rect 17960 37460 18012 37466
rect 17960 37402 18012 37408
rect 17868 36848 17920 36854
rect 17868 36790 17920 36796
rect 18708 36242 18736 38422
rect 18800 37398 18828 39200
rect 19248 38140 19300 38146
rect 19248 38082 19300 38088
rect 19260 37398 19288 38082
rect 19628 37754 19656 39200
rect 19984 38820 20036 38826
rect 19984 38762 20036 38768
rect 19628 37726 19932 37754
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19904 37398 19932 37726
rect 18788 37392 18840 37398
rect 18788 37334 18840 37340
rect 19248 37392 19300 37398
rect 19248 37334 19300 37340
rect 19892 37392 19944 37398
rect 19892 37334 19944 37340
rect 19340 36848 19392 36854
rect 19340 36790 19392 36796
rect 19524 36848 19576 36854
rect 19524 36790 19576 36796
rect 19064 36576 19116 36582
rect 19064 36518 19116 36524
rect 18696 36236 18748 36242
rect 18696 36178 18748 36184
rect 18696 34468 18748 34474
rect 18696 34410 18748 34416
rect 18708 34066 18736 34410
rect 18696 34060 18748 34066
rect 18696 34002 18748 34008
rect 18236 33992 18288 33998
rect 18236 33934 18288 33940
rect 18880 33992 18932 33998
rect 18880 33934 18932 33940
rect 17684 33652 17736 33658
rect 17684 33594 17736 33600
rect 17590 33552 17646 33561
rect 17590 33487 17592 33496
rect 17644 33487 17646 33496
rect 17592 33458 17644 33464
rect 17592 31748 17644 31754
rect 17592 31690 17644 31696
rect 17604 31414 17632 31690
rect 17592 31408 17644 31414
rect 17592 31350 17644 31356
rect 17592 27328 17644 27334
rect 17592 27270 17644 27276
rect 17604 27130 17632 27270
rect 17592 27124 17644 27130
rect 17592 27066 17644 27072
rect 17592 26308 17644 26314
rect 17592 26250 17644 26256
rect 17316 21558 17368 21564
rect 17420 21542 17540 21570
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17144 20874 17172 21422
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17132 20868 17184 20874
rect 17132 20810 17184 20816
rect 17236 20806 17264 21354
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16868 12646 16896 20470
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16960 13326 16988 18566
rect 17144 18290 17172 18566
rect 17236 18426 17264 18634
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17052 16658 17080 17138
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17144 16658 17172 16730
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17236 16250 17264 16390
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17328 15994 17356 18906
rect 17052 15966 17356 15994
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 17052 12434 17080 15966
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17236 15366 17264 15846
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 16960 12406 17080 12434
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16960 7478 16988 12406
rect 17144 11830 17172 15302
rect 17328 14618 17356 15506
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17236 12918 17264 13738
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 17236 7970 17264 12582
rect 17328 11626 17356 14554
rect 17420 12850 17448 21542
rect 17500 21412 17552 21418
rect 17500 21354 17552 21360
rect 17512 21146 17540 21354
rect 17500 21140 17552 21146
rect 17500 21082 17552 21088
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17512 15706 17540 20810
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17604 15570 17632 26250
rect 17696 15570 17724 33594
rect 17868 30184 17920 30190
rect 17868 30126 17920 30132
rect 17776 28416 17828 28422
rect 17776 28358 17828 28364
rect 17788 28150 17816 28358
rect 17776 28144 17828 28150
rect 17776 28086 17828 28092
rect 17788 25226 17816 28086
rect 17880 27010 17908 30126
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17972 27146 18000 27814
rect 17972 27118 18092 27146
rect 17880 26982 18000 27010
rect 17868 26920 17920 26926
rect 17868 26862 17920 26868
rect 17776 25220 17828 25226
rect 17776 25162 17828 25168
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17788 16454 17816 21626
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17684 14544 17736 14550
rect 17684 14486 17736 14492
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17316 11620 17368 11626
rect 17316 11562 17368 11568
rect 17052 7942 17264 7970
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16396 1352 16448 1358
rect 16396 1294 16448 1300
rect 16500 800 16528 3402
rect 16684 3194 16712 3470
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16776 800 16804 4014
rect 17052 3602 17080 7942
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17328 5846 17356 6054
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17236 5574 17264 5782
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17236 3505 17264 3538
rect 17222 3496 17278 3505
rect 17132 3460 17184 3466
rect 17222 3431 17278 3440
rect 17132 3402 17184 3408
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16960 800 16988 2926
rect 17144 800 17172 3402
rect 17328 800 17356 4626
rect 17420 3058 17448 12786
rect 17696 8906 17724 14486
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 17788 7562 17816 16050
rect 17880 16046 17908 26862
rect 17972 26790 18000 26982
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 18064 24614 18092 27118
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 18052 24608 18104 24614
rect 18052 24550 18104 24556
rect 18064 22094 18092 24550
rect 17972 22066 18092 22094
rect 17972 21010 18000 22066
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 18156 19922 18184 27066
rect 18248 23526 18276 33934
rect 18512 33924 18564 33930
rect 18512 33866 18564 33872
rect 18524 30666 18552 33866
rect 18892 33454 18920 33934
rect 18880 33448 18932 33454
rect 18880 33390 18932 33396
rect 18696 33312 18748 33318
rect 18696 33254 18748 33260
rect 18512 30660 18564 30666
rect 18512 30602 18564 30608
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18236 23520 18288 23526
rect 18236 23462 18288 23468
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17972 18290 18000 18702
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 18064 16046 18092 19382
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 18340 16182 18368 16458
rect 18328 16176 18380 16182
rect 18328 16118 18380 16124
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17880 15570 17908 15642
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 18156 15366 18184 15914
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17972 12306 18000 14894
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17972 11830 18000 12242
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17696 7534 17816 7562
rect 17592 3664 17644 3670
rect 17590 3632 17592 3641
rect 17644 3632 17646 3641
rect 17590 3567 17646 3576
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17696 2666 17724 7534
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17512 2638 17724 2666
rect 17512 1193 17540 2638
rect 17788 2582 17816 7414
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17880 3534 17908 3606
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17866 3360 17922 3369
rect 17866 3295 17922 3304
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17684 2508 17736 2514
rect 17604 2468 17684 2496
rect 17498 1184 17554 1193
rect 17498 1119 17554 1128
rect 17604 800 17632 2468
rect 17684 2450 17736 2456
rect 17880 1714 17908 3295
rect 17788 1686 17908 1714
rect 17788 800 17816 1686
rect 17972 800 18000 4626
rect 18064 2922 18092 7142
rect 18340 4078 18368 16118
rect 18432 15570 18460 24754
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18432 11762 18460 15506
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18524 10130 18552 30602
rect 18604 28008 18656 28014
rect 18602 27976 18604 27985
rect 18656 27976 18658 27985
rect 18602 27911 18658 27920
rect 18708 12434 18736 33254
rect 19076 31822 19104 36518
rect 19156 35624 19208 35630
rect 19156 35566 19208 35572
rect 19168 35290 19196 35566
rect 19156 35284 19208 35290
rect 19156 35226 19208 35232
rect 19352 34542 19380 36790
rect 19536 36718 19564 36790
rect 19524 36712 19576 36718
rect 19524 36654 19576 36660
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19996 35154 20024 38762
rect 20548 37210 20576 39200
rect 21376 37398 21404 39200
rect 21364 37392 21416 37398
rect 21364 37334 21416 37340
rect 20812 37324 20864 37330
rect 20812 37266 20864 37272
rect 20548 37182 20760 37210
rect 20732 36854 20760 37182
rect 20352 36848 20404 36854
rect 20352 36790 20404 36796
rect 20720 36848 20772 36854
rect 20720 36790 20772 36796
rect 20260 36644 20312 36650
rect 20260 36586 20312 36592
rect 20168 35760 20220 35766
rect 20168 35702 20220 35708
rect 19984 35148 20036 35154
rect 19984 35090 20036 35096
rect 19340 34536 19392 34542
rect 19340 34478 19392 34484
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19892 33516 19944 33522
rect 19892 33458 19944 33464
rect 19156 33448 19208 33454
rect 19156 33390 19208 33396
rect 19064 31816 19116 31822
rect 19064 31758 19116 31764
rect 19168 31498 19196 33390
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19340 31748 19392 31754
rect 19340 31690 19392 31696
rect 19076 31470 19196 31498
rect 18970 31376 19026 31385
rect 18970 31311 18972 31320
rect 19024 31311 19026 31320
rect 18972 31282 19024 31288
rect 19076 31226 19104 31470
rect 19352 31414 19380 31690
rect 19340 31408 19392 31414
rect 19168 31356 19340 31362
rect 19168 31350 19392 31356
rect 19524 31408 19576 31414
rect 19524 31350 19576 31356
rect 19614 31376 19670 31385
rect 19168 31346 19380 31350
rect 19156 31340 19380 31346
rect 19208 31334 19380 31340
rect 19156 31282 19208 31288
rect 19432 31272 19484 31278
rect 19352 31232 19432 31260
rect 19352 31226 19380 31232
rect 19076 31198 19380 31226
rect 19432 31214 19484 31220
rect 19536 31210 19564 31350
rect 19614 31311 19616 31320
rect 19668 31311 19670 31320
rect 19616 31282 19668 31288
rect 19524 31204 19576 31210
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 18800 28422 18828 30534
rect 18972 29504 19024 29510
rect 18972 29446 19024 29452
rect 18788 28416 18840 28422
rect 18788 28358 18840 28364
rect 18878 28112 18934 28121
rect 18878 28047 18934 28056
rect 18892 28014 18920 28047
rect 18880 28008 18932 28014
rect 18880 27950 18932 27956
rect 18892 25838 18920 27950
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18800 15570 18828 21014
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 18984 14890 19012 29446
rect 19076 29306 19104 31198
rect 19524 31146 19576 31152
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19432 30864 19484 30870
rect 19432 30806 19484 30812
rect 19064 29300 19116 29306
rect 19064 29242 19116 29248
rect 19076 28121 19104 29242
rect 19248 28416 19300 28422
rect 19248 28358 19300 28364
rect 19062 28112 19118 28121
rect 19062 28047 19118 28056
rect 19064 28008 19116 28014
rect 19064 27950 19116 27956
rect 19154 27976 19210 27985
rect 19076 26450 19104 27950
rect 19154 27911 19210 27920
rect 19168 27878 19196 27911
rect 19260 27878 19288 28358
rect 19340 27940 19392 27946
rect 19340 27882 19392 27888
rect 19156 27872 19208 27878
rect 19156 27814 19208 27820
rect 19248 27872 19300 27878
rect 19248 27814 19300 27820
rect 19064 26444 19116 26450
rect 19064 26386 19116 26392
rect 19064 25832 19116 25838
rect 19064 25774 19116 25780
rect 19076 24342 19104 25774
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 19248 22500 19300 22506
rect 19248 22442 19300 22448
rect 19260 19990 19288 22442
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19352 17882 19380 27882
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 18984 14770 19012 14826
rect 19156 14816 19208 14822
rect 18984 14764 19156 14770
rect 18984 14758 19208 14764
rect 18984 14742 19196 14758
rect 18984 14482 19012 14742
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18616 12406 18736 12434
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18524 9654 18552 10066
rect 18616 10062 18644 12406
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18144 3664 18196 3670
rect 18142 3632 18144 3641
rect 18196 3632 18198 3641
rect 18142 3567 18198 3576
rect 18234 3496 18290 3505
rect 18234 3431 18236 3440
rect 18288 3431 18290 3440
rect 18236 3402 18288 3408
rect 18144 3392 18196 3398
rect 18142 3360 18144 3369
rect 18196 3360 18198 3369
rect 18142 3295 18198 3304
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 18064 1766 18092 2858
rect 18052 1760 18104 1766
rect 18052 1702 18104 1708
rect 18156 800 18184 2926
rect 18340 800 18368 3878
rect 18432 2106 18460 6122
rect 18616 5098 18644 9998
rect 18696 9988 18748 9994
rect 18696 9930 18748 9936
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18524 3058 18552 3538
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18420 2100 18472 2106
rect 18420 2042 18472 2048
rect 18616 800 18644 4626
rect 18708 2922 18736 9930
rect 18800 9518 18828 10066
rect 19260 9586 19288 15982
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19352 15162 19380 15506
rect 19444 15502 19472 30806
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19904 28422 19932 33458
rect 20180 31754 20208 35702
rect 19996 31726 20208 31754
rect 19892 28416 19944 28422
rect 19892 28358 19944 28364
rect 19892 28144 19944 28150
rect 19892 28086 19944 28092
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19904 27130 19932 28086
rect 19892 27124 19944 27130
rect 19892 27066 19944 27072
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19892 25764 19944 25770
rect 19892 25706 19944 25712
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19904 25294 19932 25706
rect 19892 25288 19944 25294
rect 19892 25230 19944 25236
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19536 23866 19564 24006
rect 19628 23866 19656 24142
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19616 23860 19668 23866
rect 19616 23802 19668 23808
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19524 15088 19576 15094
rect 19338 15056 19394 15065
rect 19338 14991 19394 15000
rect 19522 15056 19524 15065
rect 19616 15088 19668 15094
rect 19576 15056 19578 15065
rect 19616 15030 19668 15036
rect 19706 15056 19762 15065
rect 19522 14991 19578 15000
rect 19352 14890 19380 14991
rect 19430 14920 19486 14929
rect 19340 14884 19392 14890
rect 19628 14890 19656 15030
rect 19706 14991 19762 15000
rect 19720 14958 19748 14991
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19430 14855 19432 14864
rect 19340 14826 19392 14832
rect 19484 14855 19486 14864
rect 19616 14884 19668 14890
rect 19432 14826 19484 14832
rect 19616 14826 19668 14832
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19338 14648 19394 14657
rect 19580 14640 19876 14660
rect 19338 14583 19394 14592
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18800 4010 18828 9454
rect 19352 9178 19380 14583
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19536 9364 19564 9454
rect 19444 9336 19564 9364
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19352 8430 19380 9114
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19352 7002 19380 7346
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19444 6866 19472 9336
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19904 8498 19932 23054
rect 19892 8492 19944 8498
rect 19892 8434 19944 8440
rect 19996 8430 20024 31726
rect 20076 31204 20128 31210
rect 20076 31146 20128 31152
rect 20088 31113 20116 31146
rect 20074 31104 20130 31113
rect 20074 31039 20130 31048
rect 20272 29594 20300 36586
rect 20364 31754 20392 36790
rect 20536 33380 20588 33386
rect 20536 33322 20588 33328
rect 20548 31754 20576 33322
rect 20364 31726 20484 31754
rect 20548 31726 20668 31754
rect 20272 29566 20392 29594
rect 20168 28416 20220 28422
rect 20168 28358 20220 28364
rect 20076 28144 20128 28150
rect 20076 28086 20128 28092
rect 20088 10606 20116 28086
rect 20180 24070 20208 28358
rect 20364 28257 20392 29566
rect 20350 28248 20406 28257
rect 20350 28183 20406 28192
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 20272 25702 20300 28018
rect 20352 26036 20404 26042
rect 20352 25978 20404 25984
rect 20364 25838 20392 25978
rect 20352 25832 20404 25838
rect 20352 25774 20404 25780
rect 20260 25696 20312 25702
rect 20260 25638 20312 25644
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 20180 19854 20208 24006
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 20272 17218 20300 25638
rect 20456 22234 20484 31726
rect 20536 28620 20588 28626
rect 20536 28562 20588 28568
rect 20548 28422 20576 28562
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 20536 27872 20588 27878
rect 20536 27814 20588 27820
rect 20548 27674 20576 27814
rect 20536 27668 20588 27674
rect 20536 27610 20588 27616
rect 20640 23882 20668 31726
rect 20824 30870 20852 37266
rect 21548 35012 21600 35018
rect 21548 34954 21600 34960
rect 20996 33448 21048 33454
rect 20996 33390 21048 33396
rect 21008 31754 21036 33390
rect 21364 33380 21416 33386
rect 21364 33322 21416 33328
rect 21272 32836 21324 32842
rect 21272 32778 21324 32784
rect 21008 31726 21220 31754
rect 20812 30864 20864 30870
rect 20812 30806 20864 30812
rect 20812 28620 20864 28626
rect 20812 28562 20864 28568
rect 20720 26512 20772 26518
rect 20718 26480 20720 26489
rect 20772 26480 20774 26489
rect 20718 26415 20774 26424
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20548 23866 20668 23882
rect 20536 23860 20668 23866
rect 20588 23854 20668 23860
rect 20536 23802 20588 23808
rect 20628 23792 20680 23798
rect 20628 23734 20680 23740
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20180 17190 20300 17218
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 20088 10130 20116 10542
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 20180 7206 20208 17190
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20272 15026 20300 15098
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20272 8498 20300 14418
rect 20364 9654 20392 17682
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20456 13462 20484 15438
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20548 14929 20576 14962
rect 20534 14920 20590 14929
rect 20534 14855 20590 14864
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20548 13190 20576 14758
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20640 12434 20668 23734
rect 20732 18601 20760 24142
rect 20718 18592 20774 18601
rect 20718 18527 20774 18536
rect 20718 15192 20774 15201
rect 20718 15127 20774 15136
rect 20732 14822 20760 15127
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20548 12406 20668 12434
rect 20444 12368 20496 12374
rect 20444 12310 20496 12316
rect 20352 9648 20404 9654
rect 20352 9590 20404 9596
rect 20456 8634 20484 12310
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20260 6112 20312 6118
rect 20364 6089 20392 6190
rect 20260 6054 20312 6060
rect 20350 6080 20406 6089
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 18878 5264 18934 5273
rect 18878 5199 18934 5208
rect 18788 4004 18840 4010
rect 18788 3946 18840 3952
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 18800 800 18828 2926
rect 18892 2582 18920 5199
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 18984 800 19012 3878
rect 19168 3126 19196 3946
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 19076 2961 19104 3062
rect 19062 2952 19118 2961
rect 19062 2887 19118 2896
rect 19260 2774 19288 4014
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19352 3738 19380 3878
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19168 2746 19288 2774
rect 19168 800 19196 2746
rect 19352 800 19380 2926
rect 19444 1714 19472 3334
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19904 2394 19932 4626
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19996 2854 20024 4490
rect 20088 3602 20116 4694
rect 20166 3768 20222 3777
rect 20166 3703 20222 3712
rect 20180 3670 20208 3703
rect 20168 3664 20220 3670
rect 20168 3606 20220 3612
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 20180 2990 20208 3130
rect 20168 2984 20220 2990
rect 20074 2952 20130 2961
rect 20168 2926 20220 2932
rect 20074 2887 20130 2896
rect 20088 2854 20116 2887
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 20166 2680 20222 2689
rect 20166 2615 20222 2624
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19812 2366 19932 2394
rect 19444 1686 19656 1714
rect 19628 800 19656 1686
rect 19812 800 19840 2366
rect 19996 800 20024 2450
rect 20180 800 20208 2615
rect 16212 128 16264 134
rect 16212 70 16264 76
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19338 0 19394 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20272 202 20300 6054
rect 20350 6015 20406 6024
rect 20352 4004 20404 4010
rect 20352 3946 20404 3952
rect 20364 800 20392 3946
rect 20456 3194 20484 6938
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 20260 196 20312 202
rect 20260 138 20312 144
rect 20350 0 20406 800
rect 20456 678 20484 2858
rect 20548 2582 20576 12406
rect 20824 10130 20852 28562
rect 20996 28552 21048 28558
rect 20996 28494 21048 28500
rect 20904 25764 20956 25770
rect 20904 25706 20956 25712
rect 20916 25498 20944 25706
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 21008 16658 21036 28494
rect 21192 27849 21220 31726
rect 21284 31414 21312 32778
rect 21376 31754 21404 33322
rect 21376 31726 21496 31754
rect 21272 31408 21324 31414
rect 21272 31350 21324 31356
rect 21178 27840 21234 27849
rect 21178 27775 21234 27784
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 21100 26450 21128 26862
rect 21088 26444 21140 26450
rect 21088 26386 21140 26392
rect 21192 25430 21220 27775
rect 21364 27668 21416 27674
rect 21364 27610 21416 27616
rect 21272 26444 21324 26450
rect 21272 26386 21324 26392
rect 21284 26314 21312 26386
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 21180 25424 21232 25430
rect 21180 25366 21232 25372
rect 21088 22160 21140 22166
rect 21088 22102 21140 22108
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20640 9722 20668 9930
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20640 3738 20668 7278
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20626 3632 20682 3641
rect 20626 3567 20682 3576
rect 20640 3534 20668 3567
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20536 2576 20588 2582
rect 20536 2518 20588 2524
rect 20640 800 20668 2858
rect 20732 921 20760 6054
rect 20824 5914 20852 6054
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20718 912 20774 921
rect 20718 847 20774 856
rect 20824 800 20852 3402
rect 20916 3194 20944 7482
rect 21100 6390 21128 22102
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 21088 6384 21140 6390
rect 21088 6326 21140 6332
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21008 800 21036 4626
rect 21192 4622 21220 10066
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 21192 2689 21220 3538
rect 21284 3346 21312 8910
rect 21376 6186 21404 27610
rect 21468 15910 21496 31726
rect 21560 27674 21588 34954
rect 21640 34060 21692 34066
rect 21640 34002 21692 34008
rect 21652 31754 21680 34002
rect 21824 33992 21876 33998
rect 21824 33934 21876 33940
rect 21652 31726 21772 31754
rect 21548 27668 21600 27674
rect 21548 27610 21600 27616
rect 21640 27124 21692 27130
rect 21640 27066 21692 27072
rect 21548 27056 21600 27062
rect 21546 27024 21548 27033
rect 21600 27024 21602 27033
rect 21546 26959 21602 26968
rect 21548 26580 21600 26586
rect 21548 26522 21600 26528
rect 21560 26489 21588 26522
rect 21652 26518 21680 27066
rect 21640 26512 21692 26518
rect 21546 26480 21602 26489
rect 21640 26454 21692 26460
rect 21546 26415 21602 26424
rect 21744 25650 21772 31726
rect 21836 29306 21864 33934
rect 21928 32434 21956 39238
rect 22282 39200 22338 40000
rect 23110 39200 23166 40000
rect 24030 39200 24086 40000
rect 24858 39200 24914 40000
rect 25778 39200 25834 40000
rect 26698 39200 26754 40000
rect 27526 39200 27582 40000
rect 28446 39200 28502 40000
rect 29274 39200 29330 40000
rect 30194 39200 30250 40000
rect 31022 39200 31078 40000
rect 31942 39200 31998 40000
rect 32770 39200 32826 40000
rect 33690 39200 33746 40000
rect 34518 39200 34574 40000
rect 35438 39200 35494 40000
rect 36266 39200 36322 40000
rect 37186 39200 37242 40000
rect 37464 39636 37516 39642
rect 37464 39578 37516 39584
rect 22296 37466 22324 39200
rect 23020 37664 23072 37670
rect 23020 37606 23072 37612
rect 22284 37460 22336 37466
rect 22284 37402 22336 37408
rect 23032 37398 23060 37606
rect 23124 37482 23152 39200
rect 23940 38956 23992 38962
rect 23940 38898 23992 38904
rect 23296 38548 23348 38554
rect 23296 38490 23348 38496
rect 23124 37466 23244 37482
rect 23124 37460 23256 37466
rect 23124 37454 23204 37460
rect 23204 37402 23256 37408
rect 23020 37392 23072 37398
rect 23020 37334 23072 37340
rect 22100 37256 22152 37262
rect 22100 37198 22152 37204
rect 22112 36174 22140 37198
rect 22100 36168 22152 36174
rect 22100 36110 22152 36116
rect 22836 34128 22888 34134
rect 22836 34070 22888 34076
rect 22100 33380 22152 33386
rect 22100 33322 22152 33328
rect 22006 33008 22062 33017
rect 22006 32943 22008 32952
rect 22060 32943 22062 32952
rect 22008 32914 22060 32920
rect 21916 32428 21968 32434
rect 21916 32370 21968 32376
rect 22112 32366 22140 33322
rect 22192 33040 22244 33046
rect 22190 33008 22192 33017
rect 22244 33008 22246 33017
rect 22190 32943 22246 32952
rect 22376 32972 22428 32978
rect 22376 32914 22428 32920
rect 22388 32842 22416 32914
rect 22652 32904 22704 32910
rect 22652 32846 22704 32852
rect 22376 32836 22428 32842
rect 22376 32778 22428 32784
rect 22100 32360 22152 32366
rect 22100 32302 22152 32308
rect 22374 32328 22430 32337
rect 22374 32263 22376 32272
rect 22428 32263 22430 32272
rect 22468 32292 22520 32298
rect 22376 32234 22428 32240
rect 22468 32234 22520 32240
rect 22284 32224 22336 32230
rect 22284 32166 22336 32172
rect 22296 31822 22324 32166
rect 22284 31816 22336 31822
rect 22284 31758 22336 31764
rect 22480 31736 22508 32234
rect 22560 31748 22612 31754
rect 22480 31708 22560 31736
rect 22560 31690 22612 31696
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 21824 29300 21876 29306
rect 21824 29242 21876 29248
rect 22100 28484 22152 28490
rect 22100 28426 22152 28432
rect 22008 27464 22060 27470
rect 22008 27406 22060 27412
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 21836 26994 21864 27066
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 21928 26450 21956 27270
rect 22020 26994 22048 27406
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 21916 26444 21968 26450
rect 21916 26386 21968 26392
rect 21744 25622 21956 25650
rect 21744 25362 21772 25622
rect 21928 25498 21956 25622
rect 21824 25492 21876 25498
rect 21824 25434 21876 25440
rect 21916 25492 21968 25498
rect 21916 25434 21968 25440
rect 21732 25356 21784 25362
rect 21732 25298 21784 25304
rect 21836 25158 21864 25434
rect 22112 25362 22140 28426
rect 22100 25356 22152 25362
rect 22100 25298 22152 25304
rect 21824 25152 21876 25158
rect 21824 25094 21876 25100
rect 21916 25152 21968 25158
rect 21916 25094 21968 25100
rect 21836 24410 21864 25094
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21732 20868 21784 20874
rect 21732 20810 21784 20816
rect 21638 19272 21694 19281
rect 21638 19207 21640 19216
rect 21692 19207 21694 19216
rect 21640 19178 21692 19184
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21364 6180 21416 6186
rect 21364 6122 21416 6128
rect 21468 3482 21496 15846
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21560 3670 21588 12582
rect 21744 11218 21772 20810
rect 21928 19514 21956 25094
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 22112 18426 22140 23530
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 21822 17912 21878 17921
rect 21822 17847 21878 17856
rect 21836 17678 21864 17847
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 22112 12986 22140 13738
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22204 12434 22232 29446
rect 22572 28762 22600 31690
rect 22560 28756 22612 28762
rect 22560 28698 22612 28704
rect 22376 28008 22428 28014
rect 22376 27950 22428 27956
rect 22284 27056 22336 27062
rect 22282 27024 22284 27033
rect 22336 27024 22338 27033
rect 22282 26959 22338 26968
rect 22388 12986 22416 27950
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22480 22094 22508 25298
rect 22560 24608 22612 24614
rect 22560 24550 22612 24556
rect 22572 24274 22600 24550
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22480 22066 22600 22094
rect 22466 20632 22522 20641
rect 22466 20567 22468 20576
rect 22520 20567 22522 20576
rect 22468 20538 22520 20544
rect 22466 20496 22522 20505
rect 22466 20431 22468 20440
rect 22520 20431 22522 20440
rect 22468 20402 22520 20408
rect 22468 19168 22520 19174
rect 22466 19136 22468 19145
rect 22520 19136 22522 19145
rect 22466 19071 22522 19080
rect 22468 13456 22520 13462
rect 22466 13424 22468 13433
rect 22520 13424 22522 13433
rect 22466 13359 22522 13368
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22572 12782 22600 22066
rect 22664 18766 22692 32846
rect 22744 24676 22796 24682
rect 22744 24618 22796 24624
rect 22756 20602 22784 24618
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22742 19272 22798 19281
rect 22742 19207 22798 19216
rect 22756 19174 22784 19207
rect 22744 19168 22796 19174
rect 22744 19110 22796 19116
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22664 17864 22692 18702
rect 22664 17836 22784 17864
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22664 17202 22692 17682
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22756 13802 22784 17836
rect 22848 14958 22876 34070
rect 23020 32496 23072 32502
rect 23020 32438 23072 32444
rect 23032 27402 23060 32438
rect 23308 28014 23336 38490
rect 23480 37120 23532 37126
rect 23480 37062 23532 37068
rect 23492 36786 23520 37062
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23664 35148 23716 35154
rect 23664 35090 23716 35096
rect 23388 28484 23440 28490
rect 23388 28426 23440 28432
rect 23400 28218 23428 28426
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 23296 28008 23348 28014
rect 23296 27950 23348 27956
rect 23204 27668 23256 27674
rect 23204 27610 23256 27616
rect 23020 27396 23072 27402
rect 23020 27338 23072 27344
rect 23216 26858 23244 27610
rect 23676 27538 23704 35090
rect 23664 27532 23716 27538
rect 23664 27474 23716 27480
rect 23204 26852 23256 26858
rect 23204 26794 23256 26800
rect 22928 25832 22980 25838
rect 22928 25774 22980 25780
rect 22940 18154 22968 25774
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 23032 24070 23060 24142
rect 23020 24064 23072 24070
rect 23020 24006 23072 24012
rect 23018 20632 23074 20641
rect 23018 20567 23020 20576
rect 23072 20567 23074 20576
rect 23020 20538 23072 20544
rect 23018 20496 23074 20505
rect 23018 20431 23020 20440
rect 23072 20431 23074 20440
rect 23020 20402 23072 20408
rect 23020 19236 23072 19242
rect 23020 19178 23072 19184
rect 23032 19145 23060 19178
rect 23018 19136 23074 19145
rect 23018 19071 23074 19080
rect 23018 18592 23074 18601
rect 23018 18527 23074 18536
rect 22928 18148 22980 18154
rect 22928 18090 22980 18096
rect 23032 17814 23060 18527
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22744 13796 22796 13802
rect 22744 13738 22796 13744
rect 22560 12776 22612 12782
rect 22560 12718 22612 12724
rect 22112 12406 22232 12434
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 22112 8838 22140 12406
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21652 5778 21680 6122
rect 21640 5772 21692 5778
rect 21640 5714 21692 5720
rect 21744 5166 21772 8774
rect 21822 6760 21878 6769
rect 21822 6695 21878 6704
rect 21836 6390 21864 6695
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 21928 6390 21956 6598
rect 21824 6384 21876 6390
rect 21824 6326 21876 6332
rect 21916 6384 21968 6390
rect 21916 6326 21968 6332
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 21836 6089 21864 6190
rect 21822 6080 21878 6089
rect 21822 6015 21878 6024
rect 22020 5846 22048 6598
rect 22008 5840 22060 5846
rect 22008 5782 22060 5788
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 21548 3664 21600 3670
rect 21548 3606 21600 3612
rect 21744 3505 21772 4626
rect 21916 4208 21968 4214
rect 21916 4150 21968 4156
rect 21928 3754 21956 4150
rect 21928 3726 22048 3754
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 21730 3496 21786 3505
rect 21468 3454 21680 3482
rect 21652 3346 21680 3454
rect 21730 3431 21786 3440
rect 21836 3398 21864 3606
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21824 3392 21876 3398
rect 21284 3318 21588 3346
rect 21652 3318 21772 3346
rect 21824 3334 21876 3340
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21178 2680 21234 2689
rect 21178 2615 21234 2624
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21192 800 21220 2450
rect 21272 2372 21324 2378
rect 21272 2314 21324 2320
rect 21284 1970 21312 2314
rect 21272 1964 21324 1970
rect 21272 1906 21324 1912
rect 21376 800 21404 2790
rect 21560 1057 21588 3318
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21546 1048 21602 1057
rect 21546 983 21602 992
rect 21652 800 21680 3130
rect 21744 2582 21772 3318
rect 21928 3210 21956 3538
rect 22020 3466 22048 3726
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 22006 3360 22062 3369
rect 22006 3295 22062 3304
rect 21836 3194 21956 3210
rect 21824 3188 21956 3194
rect 21876 3182 21956 3188
rect 21824 3130 21876 3136
rect 21732 2576 21784 2582
rect 21732 2518 21784 2524
rect 21824 2372 21876 2378
rect 21824 2314 21876 2320
rect 21836 800 21864 2314
rect 22020 800 22048 3295
rect 22112 2990 22140 8774
rect 22848 5710 22876 14894
rect 22940 12434 22968 15438
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23032 12782 23060 12922
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 22940 12406 23060 12434
rect 23032 8430 23060 12406
rect 23020 8424 23072 8430
rect 23020 8366 23072 8372
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22282 3632 22338 3641
rect 22282 3567 22338 3576
rect 22296 3534 22324 3567
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22204 800 22232 2926
rect 22468 2304 22520 2310
rect 22468 2246 22520 2252
rect 22480 800 22508 2246
rect 22664 800 22692 4626
rect 22848 4554 22876 5646
rect 22940 5302 22968 7346
rect 22928 5296 22980 5302
rect 22928 5238 22980 5244
rect 22836 4548 22888 4554
rect 22836 4490 22888 4496
rect 23032 4078 23060 8366
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22848 800 22876 3538
rect 23124 2582 23152 24550
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23204 20256 23256 20262
rect 23204 20198 23256 20204
rect 23216 5234 23244 20198
rect 23308 17270 23336 24142
rect 23952 23730 23980 38898
rect 24044 37398 24072 39200
rect 24872 37466 24900 39200
rect 25688 39024 25740 39030
rect 25688 38966 25740 38972
rect 24952 38072 25004 38078
rect 24952 38014 25004 38020
rect 24860 37460 24912 37466
rect 24860 37402 24912 37408
rect 24032 37392 24084 37398
rect 24032 37334 24084 37340
rect 24124 37324 24176 37330
rect 24124 37266 24176 37272
rect 24032 31680 24084 31686
rect 24030 31648 24032 31657
rect 24084 31648 24086 31657
rect 24030 31583 24086 31592
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23296 17264 23348 17270
rect 23296 17206 23348 17212
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23400 9382 23428 10066
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23400 7546 23428 8298
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 23112 2576 23164 2582
rect 23112 2518 23164 2524
rect 23020 2372 23072 2378
rect 23020 2314 23072 2320
rect 23032 800 23060 2314
rect 23216 800 23244 4626
rect 23400 3942 23428 5850
rect 23492 4078 23520 16186
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23676 8634 23704 14350
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23480 4072 23532 4078
rect 23480 4014 23532 4020
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23492 800 23520 2926
rect 23768 2582 23796 22578
rect 24136 22030 24164 37266
rect 24492 36848 24544 36854
rect 24492 36790 24544 36796
rect 24308 36168 24360 36174
rect 24308 36110 24360 36116
rect 24320 35222 24348 36110
rect 24504 35834 24532 36790
rect 24964 36378 24992 38014
rect 25504 37732 25556 37738
rect 25504 37674 25556 37680
rect 24768 36372 24820 36378
rect 24768 36314 24820 36320
rect 24952 36372 25004 36378
rect 24952 36314 25004 36320
rect 24492 35828 24544 35834
rect 24492 35770 24544 35776
rect 24780 35630 24808 36314
rect 24676 35624 24728 35630
rect 24676 35566 24728 35572
rect 24768 35624 24820 35630
rect 24768 35566 24820 35572
rect 25228 35624 25280 35630
rect 25228 35566 25280 35572
rect 24688 35442 24716 35566
rect 24688 35414 24900 35442
rect 24308 35216 24360 35222
rect 24308 35158 24360 35164
rect 24400 34536 24452 34542
rect 24400 34478 24452 34484
rect 24308 31136 24360 31142
rect 24308 31078 24360 31084
rect 24320 29170 24348 31078
rect 24308 29164 24360 29170
rect 24308 29106 24360 29112
rect 24216 29096 24268 29102
rect 24216 29038 24268 29044
rect 24228 28082 24256 29038
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 24216 24200 24268 24206
rect 24216 24142 24268 24148
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24124 16584 24176 16590
rect 24122 16552 24124 16561
rect 24176 16552 24178 16561
rect 24122 16487 24178 16496
rect 24032 15564 24084 15570
rect 24032 15506 24084 15512
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24044 15162 24072 15506
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 24136 13938 24164 15506
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24228 12646 24256 24142
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 24136 7177 24164 7210
rect 24122 7168 24178 7177
rect 24122 7103 24178 7112
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 23756 2576 23808 2582
rect 23756 2518 23808 2524
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 23676 800 23704 2382
rect 23860 800 23888 4014
rect 23952 3398 23980 5578
rect 24320 5370 24348 23666
rect 24412 16250 24440 34478
rect 24872 34066 24900 35414
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 24768 33924 24820 33930
rect 24768 33866 24820 33872
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24492 33448 24544 33454
rect 24492 33390 24544 33396
rect 24504 25906 24532 33390
rect 24596 31142 24624 33798
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 24780 30546 24808 33866
rect 24780 30518 24900 30546
rect 24872 30274 24900 30518
rect 25240 30394 25268 35566
rect 25320 34536 25372 34542
rect 25320 34478 25372 34484
rect 25332 33386 25360 34478
rect 25320 33380 25372 33386
rect 25320 33322 25372 33328
rect 25412 32496 25464 32502
rect 25412 32438 25464 32444
rect 25228 30388 25280 30394
rect 25228 30330 25280 30336
rect 24596 30246 24900 30274
rect 24492 25900 24544 25906
rect 24492 25842 24544 25848
rect 24504 24818 24532 25842
rect 24492 24812 24544 24818
rect 24492 24754 24544 24760
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24412 15706 24440 16186
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 24596 14618 24624 30246
rect 24676 30116 24728 30122
rect 24676 30058 24728 30064
rect 24688 17921 24716 30058
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 24780 24206 24808 29106
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 25148 23798 25176 24346
rect 25320 24336 25372 24342
rect 25320 24278 25372 24284
rect 25332 24206 25360 24278
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 25240 23798 25268 24142
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25228 23792 25280 23798
rect 25228 23734 25280 23740
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 24952 23588 25004 23594
rect 24952 23530 25004 23536
rect 24964 22094 24992 23530
rect 24964 22066 25084 22094
rect 25056 19145 25084 22066
rect 25042 19136 25098 19145
rect 25042 19071 25098 19080
rect 24674 17912 24730 17921
rect 24674 17847 24730 17856
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 25056 12434 25084 19071
rect 24964 12406 25084 12434
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24872 7342 24900 9998
rect 24860 7336 24912 7342
rect 24766 7304 24822 7313
rect 24860 7278 24912 7284
rect 24766 7239 24822 7248
rect 24780 5574 24808 7239
rect 24768 5568 24820 5574
rect 24768 5510 24820 5516
rect 24308 5364 24360 5370
rect 24308 5306 24360 5312
rect 24964 4758 24992 12406
rect 25148 10305 25176 23598
rect 25228 23112 25280 23118
rect 25228 23054 25280 23060
rect 25240 22506 25268 23054
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25332 22953 25360 22986
rect 25318 22944 25374 22953
rect 25318 22879 25374 22888
rect 25228 22500 25280 22506
rect 25228 22442 25280 22448
rect 25424 21554 25452 32438
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 25240 18329 25268 18702
rect 25226 18320 25282 18329
rect 25226 18255 25282 18264
rect 25228 11620 25280 11626
rect 25228 11562 25280 11568
rect 25240 11014 25268 11562
rect 25228 11008 25280 11014
rect 25228 10950 25280 10956
rect 25134 10296 25190 10305
rect 25134 10231 25190 10240
rect 25148 10062 25176 10231
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25332 7698 25360 18702
rect 25516 11558 25544 37674
rect 25700 31754 25728 38966
rect 25792 37482 25820 39200
rect 26148 38072 26200 38078
rect 26148 38014 26200 38020
rect 25792 37466 25912 37482
rect 25792 37460 25924 37466
rect 25792 37454 25872 37460
rect 25872 37402 25924 37408
rect 26160 37330 26188 38014
rect 26516 37732 26568 37738
rect 26516 37674 26568 37680
rect 26528 37398 26556 37674
rect 26516 37392 26568 37398
rect 26516 37334 26568 37340
rect 26148 37324 26200 37330
rect 26148 37266 26200 37272
rect 26712 36718 26740 39200
rect 27068 37732 27120 37738
rect 27068 37674 27120 37680
rect 26700 36712 26752 36718
rect 26700 36654 26752 36660
rect 26700 36576 26752 36582
rect 26700 36518 26752 36524
rect 26056 32836 26108 32842
rect 26056 32778 26108 32784
rect 25700 31726 25820 31754
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 25596 23520 25648 23526
rect 25596 23462 25648 23468
rect 25608 22166 25636 23462
rect 25596 22160 25648 22166
rect 25596 22102 25648 22108
rect 25596 21956 25648 21962
rect 25596 21898 25648 21904
rect 25608 21418 25636 21898
rect 25596 21412 25648 21418
rect 25596 21354 25648 21360
rect 25700 18766 25728 23666
rect 25688 18760 25740 18766
rect 25688 18702 25740 18708
rect 25594 17368 25650 17377
rect 25594 17303 25650 17312
rect 25608 17270 25636 17303
rect 25596 17264 25648 17270
rect 25596 17206 25648 17212
rect 25688 17264 25740 17270
rect 25688 17206 25740 17212
rect 25596 17128 25648 17134
rect 25596 17070 25648 17076
rect 25608 16726 25636 17070
rect 25596 16720 25648 16726
rect 25596 16662 25648 16668
rect 25700 16658 25728 17206
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25688 16516 25740 16522
rect 25688 16458 25740 16464
rect 25700 16046 25728 16458
rect 25792 16250 25820 31726
rect 25964 30116 26016 30122
rect 25964 30058 26016 30064
rect 25872 25288 25924 25294
rect 25872 25230 25924 25236
rect 25884 24954 25912 25230
rect 25872 24948 25924 24954
rect 25872 24890 25924 24896
rect 25884 23322 25912 24890
rect 25872 23316 25924 23322
rect 25872 23258 25924 23264
rect 25976 23202 26004 30058
rect 25884 23174 26004 23202
rect 26068 23202 26096 32778
rect 26516 31136 26568 31142
rect 26516 31078 26568 31084
rect 26148 29708 26200 29714
rect 26148 29650 26200 29656
rect 26160 29238 26188 29650
rect 26148 29232 26200 29238
rect 26148 29174 26200 29180
rect 26332 29232 26384 29238
rect 26332 29174 26384 29180
rect 26240 28552 26292 28558
rect 26240 28494 26292 28500
rect 26252 28014 26280 28494
rect 26240 28008 26292 28014
rect 26240 27950 26292 27956
rect 26148 27600 26200 27606
rect 26148 27542 26200 27548
rect 26160 23322 26188 27542
rect 26344 26602 26372 29174
rect 26252 26574 26372 26602
rect 26148 23316 26200 23322
rect 26148 23258 26200 23264
rect 26068 23174 26188 23202
rect 25884 22094 25912 23174
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 25884 22066 26004 22094
rect 25872 21616 25924 21622
rect 25872 21558 25924 21564
rect 25884 21486 25912 21558
rect 25872 21480 25924 21486
rect 25872 21422 25924 21428
rect 25780 16244 25832 16250
rect 25780 16186 25832 16192
rect 25688 16040 25740 16046
rect 25688 15982 25740 15988
rect 25976 12434 26004 22066
rect 26068 21010 26096 23054
rect 26160 23050 26188 23174
rect 26148 23044 26200 23050
rect 26148 22986 26200 22992
rect 26252 22166 26280 26574
rect 26332 26444 26384 26450
rect 26332 26386 26384 26392
rect 26344 23186 26372 26386
rect 26528 23361 26556 31078
rect 26608 29096 26660 29102
rect 26608 29038 26660 29044
rect 26514 23352 26570 23361
rect 26514 23287 26570 23296
rect 26332 23180 26384 23186
rect 26332 23122 26384 23128
rect 26516 23180 26568 23186
rect 26516 23122 26568 23128
rect 26330 23080 26386 23089
rect 26330 23015 26386 23024
rect 26344 22778 26372 23015
rect 26332 22772 26384 22778
rect 26332 22714 26384 22720
rect 26240 22160 26292 22166
rect 26240 22102 26292 22108
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26332 21480 26384 21486
rect 26332 21422 26384 21428
rect 26160 21146 26188 21422
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26148 21140 26200 21146
rect 26148 21082 26200 21088
rect 26056 21004 26108 21010
rect 26056 20946 26108 20952
rect 26252 18358 26280 21286
rect 26240 18352 26292 18358
rect 26240 18294 26292 18300
rect 26128 16584 26180 16590
rect 26180 16532 26188 16572
rect 26128 16526 26188 16532
rect 25976 12406 26096 12434
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25240 7670 25360 7698
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 24952 4752 25004 4758
rect 24952 4694 25004 4700
rect 24492 4072 24544 4078
rect 24492 4014 24544 4020
rect 24032 3596 24084 3602
rect 24032 3538 24084 3544
rect 23940 3392 23992 3398
rect 23940 3334 23992 3340
rect 24044 800 24072 3538
rect 24216 2304 24268 2310
rect 24216 2246 24268 2252
rect 24228 800 24256 2246
rect 24504 800 24532 4014
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24688 800 24716 3538
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 24872 800 24900 2858
rect 25056 800 25084 5102
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 25148 2990 25176 4762
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 25240 2854 25268 7670
rect 25320 7336 25372 7342
rect 25516 7324 25544 11494
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 25792 9926 25820 10202
rect 25872 10056 25924 10062
rect 25872 9998 25924 10004
rect 25780 9920 25832 9926
rect 25780 9862 25832 9868
rect 25884 9382 25912 9998
rect 25872 9376 25924 9382
rect 25872 9318 25924 9324
rect 25976 8294 26004 10610
rect 25964 8288 26016 8294
rect 25964 8230 26016 8236
rect 25780 7948 25832 7954
rect 25780 7890 25832 7896
rect 25792 7478 25820 7890
rect 25780 7472 25832 7478
rect 25780 7414 25832 7420
rect 25792 7342 25820 7414
rect 25372 7296 25544 7324
rect 25688 7336 25740 7342
rect 25686 7304 25688 7313
rect 25780 7336 25832 7342
rect 25740 7304 25742 7313
rect 25320 7278 25372 7284
rect 25964 7336 26016 7342
rect 25780 7278 25832 7284
rect 25962 7304 25964 7313
rect 26016 7304 26018 7313
rect 25686 7239 25742 7248
rect 25962 7239 26018 7248
rect 25964 7200 26016 7206
rect 25962 7168 25964 7177
rect 26016 7168 26018 7177
rect 25962 7103 26018 7112
rect 25688 5160 25740 5166
rect 25688 5102 25740 5108
rect 25320 4752 25372 4758
rect 25320 4694 25372 4700
rect 25332 4010 25360 4694
rect 25320 4004 25372 4010
rect 25320 3946 25372 3952
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 25332 2666 25360 3538
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25608 2990 25636 3402
rect 25596 2984 25648 2990
rect 25596 2926 25648 2932
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 25594 2816 25650 2825
rect 25240 2638 25360 2666
rect 25240 800 25268 2638
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 25332 1902 25360 2450
rect 25320 1896 25372 1902
rect 25320 1838 25372 1844
rect 25516 800 25544 2790
rect 25594 2751 25650 2760
rect 20444 672 20496 678
rect 20444 614 20496 620
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25608 746 25636 2751
rect 25700 800 25728 5102
rect 26068 4842 26096 12406
rect 25976 4814 26096 4842
rect 25976 4758 26004 4814
rect 25964 4752 26016 4758
rect 25964 4694 26016 4700
rect 25872 4684 25924 4690
rect 25872 4626 25924 4632
rect 26056 4684 26108 4690
rect 26056 4626 26108 4632
rect 25780 4004 25832 4010
rect 25780 3946 25832 3952
rect 25792 1034 25820 3946
rect 25884 1222 25912 4626
rect 25964 4072 26016 4078
rect 25964 4014 26016 4020
rect 25872 1216 25924 1222
rect 25872 1158 25924 1164
rect 25792 1006 25912 1034
rect 25884 800 25912 1006
rect 25596 740 25648 746
rect 25596 682 25648 688
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 25976 338 26004 4014
rect 26068 1018 26096 4626
rect 26160 2961 26188 16526
rect 26344 12434 26372 21422
rect 26528 20074 26556 23122
rect 26620 20262 26648 29038
rect 26608 20256 26660 20262
rect 26608 20198 26660 20204
rect 26528 20046 26648 20074
rect 26424 19916 26476 19922
rect 26424 19858 26476 19864
rect 26436 15434 26464 19858
rect 26516 18760 26568 18766
rect 26516 18702 26568 18708
rect 26528 18358 26556 18702
rect 26516 18352 26568 18358
rect 26516 18294 26568 18300
rect 26516 16584 26568 16590
rect 26514 16552 26516 16561
rect 26568 16552 26570 16561
rect 26514 16487 26570 16496
rect 26424 15428 26476 15434
rect 26424 15370 26476 15376
rect 26516 14884 26568 14890
rect 26516 14826 26568 14832
rect 26252 12406 26372 12434
rect 26252 11014 26280 12406
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26332 11824 26384 11830
rect 26332 11766 26384 11772
rect 26344 11218 26372 11766
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26436 11150 26464 12174
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 26240 11008 26292 11014
rect 26240 10950 26292 10956
rect 26252 10266 26280 10950
rect 26330 10296 26386 10305
rect 26240 10260 26292 10266
rect 26330 10231 26332 10240
rect 26240 10202 26292 10208
rect 26384 10231 26386 10240
rect 26332 10202 26384 10208
rect 26436 10146 26464 11086
rect 26252 10118 26464 10146
rect 26252 9382 26280 10118
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26252 5710 26280 9318
rect 26528 5778 26556 14826
rect 26620 7342 26648 20046
rect 26712 16250 26740 36518
rect 26792 36372 26844 36378
rect 26792 36314 26844 36320
rect 26804 31754 26832 36314
rect 26884 32904 26936 32910
rect 26884 32846 26936 32852
rect 26896 32570 26924 32846
rect 26884 32564 26936 32570
rect 26884 32506 26936 32512
rect 26976 32564 27028 32570
rect 26976 32506 27028 32512
rect 26988 32337 27016 32506
rect 26974 32328 27030 32337
rect 26974 32263 27030 32272
rect 26804 31726 27016 31754
rect 26882 30832 26938 30841
rect 26882 30767 26938 30776
rect 26792 28756 26844 28762
rect 26792 28698 26844 28704
rect 26804 20942 26832 28698
rect 26896 26450 26924 30767
rect 26884 26444 26936 26450
rect 26884 26386 26936 26392
rect 26884 26036 26936 26042
rect 26884 25978 26936 25984
rect 26896 25702 26924 25978
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26884 24064 26936 24070
rect 26884 24006 26936 24012
rect 26896 23594 26924 24006
rect 26884 23588 26936 23594
rect 26884 23530 26936 23536
rect 26884 23112 26936 23118
rect 26882 23080 26884 23089
rect 26936 23080 26938 23089
rect 26882 23015 26938 23024
rect 26884 22976 26936 22982
rect 26884 22918 26936 22924
rect 26896 22234 26924 22918
rect 26884 22228 26936 22234
rect 26884 22170 26936 22176
rect 26884 21412 26936 21418
rect 26884 21354 26936 21360
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26700 16244 26752 16250
rect 26700 16186 26752 16192
rect 26804 13394 26832 20878
rect 26896 19922 26924 21354
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26988 19854 27016 31726
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 26884 18760 26936 18766
rect 26884 18702 26936 18708
rect 26896 18222 26924 18702
rect 26884 18216 26936 18222
rect 26884 18158 26936 18164
rect 26884 17740 26936 17746
rect 26884 17682 26936 17688
rect 26896 17649 26924 17682
rect 26882 17640 26938 17649
rect 26882 17575 26938 17584
rect 26988 16726 27016 19790
rect 26976 16720 27028 16726
rect 26976 16662 27028 16668
rect 26884 15904 26936 15910
rect 26884 15846 26936 15852
rect 26896 15434 26924 15846
rect 26884 15428 26936 15434
rect 26884 15370 26936 15376
rect 26884 14884 26936 14890
rect 26884 14826 26936 14832
rect 26896 14550 26924 14826
rect 26884 14544 26936 14550
rect 26884 14486 26936 14492
rect 27080 13394 27108 37674
rect 27540 37398 27568 39200
rect 27988 38616 28040 38622
rect 27988 38558 28040 38564
rect 27528 37392 27580 37398
rect 27528 37334 27580 37340
rect 27160 37324 27212 37330
rect 27160 37266 27212 37272
rect 27172 29238 27200 37266
rect 27436 36576 27488 36582
rect 27436 36518 27488 36524
rect 27448 36242 27476 36518
rect 27436 36236 27488 36242
rect 27436 36178 27488 36184
rect 27804 36236 27856 36242
rect 27804 36178 27856 36184
rect 27252 31884 27304 31890
rect 27252 31826 27304 31832
rect 27160 29232 27212 29238
rect 27160 29174 27212 29180
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27172 28422 27200 28494
rect 27160 28416 27212 28422
rect 27160 28358 27212 28364
rect 27158 27432 27214 27441
rect 27158 27367 27160 27376
rect 27212 27367 27214 27376
rect 27160 27338 27212 27344
rect 27160 26444 27212 26450
rect 27160 26386 27212 26392
rect 27172 22710 27200 26386
rect 27160 22704 27212 22710
rect 27160 22646 27212 22652
rect 27264 20262 27292 31826
rect 27448 31754 27476 36178
rect 27816 34542 27844 36178
rect 28000 34746 28028 38558
rect 28460 37466 28488 39200
rect 28448 37460 28500 37466
rect 28448 37402 28500 37408
rect 28356 37324 28408 37330
rect 28356 37266 28408 37272
rect 28264 36644 28316 36650
rect 28264 36586 28316 36592
rect 28276 36310 28304 36586
rect 28264 36304 28316 36310
rect 28264 36246 28316 36252
rect 28080 36168 28132 36174
rect 28080 36110 28132 36116
rect 27988 34740 28040 34746
rect 27988 34682 28040 34688
rect 27804 34536 27856 34542
rect 27804 34478 27856 34484
rect 28092 34406 28120 36110
rect 27988 34400 28040 34406
rect 27988 34342 28040 34348
rect 28080 34400 28132 34406
rect 28080 34342 28132 34348
rect 27804 33584 27856 33590
rect 27804 33526 27856 33532
rect 27712 31884 27764 31890
rect 27712 31826 27764 31832
rect 27356 31726 27476 31754
rect 27528 31748 27580 31754
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 27252 20256 27304 20262
rect 27252 20198 27304 20204
rect 27172 19718 27200 20198
rect 27264 19922 27292 20198
rect 27252 19916 27304 19922
rect 27252 19858 27304 19864
rect 27160 19712 27212 19718
rect 27160 19654 27212 19660
rect 26792 13388 26844 13394
rect 26792 13330 26844 13336
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 27172 11830 27200 19654
rect 27356 19310 27384 31726
rect 27528 31690 27580 31696
rect 27540 31657 27568 31690
rect 27526 31648 27582 31657
rect 27526 31583 27582 31592
rect 27620 31408 27672 31414
rect 27526 31376 27582 31385
rect 27620 31350 27672 31356
rect 27526 31311 27582 31320
rect 27540 31142 27568 31311
rect 27528 31136 27580 31142
rect 27528 31078 27580 31084
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27540 26858 27568 27406
rect 27528 26852 27580 26858
rect 27528 26794 27580 26800
rect 27528 19916 27580 19922
rect 27528 19858 27580 19864
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 27356 16182 27384 16390
rect 27344 16176 27396 16182
rect 27344 16118 27396 16124
rect 27344 13796 27396 13802
rect 27344 13738 27396 13744
rect 27252 13388 27304 13394
rect 27356 13376 27384 13738
rect 27304 13348 27384 13376
rect 27252 13330 27304 13336
rect 27160 11824 27212 11830
rect 27160 11766 27212 11772
rect 26792 11280 26844 11286
rect 26844 11228 27016 11234
rect 26792 11222 27016 11228
rect 26804 11206 27016 11222
rect 26988 11200 27016 11206
rect 27252 11212 27304 11218
rect 26988 11172 27252 11200
rect 27252 11154 27304 11160
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26896 9602 26924 11086
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27264 10266 27292 10542
rect 27252 10260 27304 10266
rect 27252 10202 27304 10208
rect 27068 10124 27120 10130
rect 27068 10066 27120 10072
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26804 9574 26924 9602
rect 26804 7546 26832 9574
rect 26884 9512 26936 9518
rect 26884 9454 26936 9460
rect 26896 8906 26924 9454
rect 26884 8900 26936 8906
rect 26884 8842 26936 8848
rect 26792 7540 26844 7546
rect 26792 7482 26844 7488
rect 26608 7336 26660 7342
rect 26608 7278 26660 7284
rect 26516 5772 26568 5778
rect 26516 5714 26568 5720
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 26332 5160 26384 5166
rect 26332 5102 26384 5108
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26146 2952 26202 2961
rect 26252 2922 26280 3334
rect 26146 2887 26202 2896
rect 26240 2916 26292 2922
rect 26240 2858 26292 2864
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 26056 1012 26108 1018
rect 26056 954 26108 960
rect 26160 898 26188 2790
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 26252 1970 26280 2450
rect 26240 1964 26292 1970
rect 26240 1906 26292 1912
rect 26068 870 26188 898
rect 26068 800 26096 870
rect 26344 800 26372 5102
rect 26884 4684 26936 4690
rect 26988 4672 27016 9998
rect 27080 9926 27108 10066
rect 27068 9920 27120 9926
rect 27068 9862 27120 9868
rect 27356 8022 27384 13348
rect 27540 11694 27568 19858
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27344 8016 27396 8022
rect 27344 7958 27396 7964
rect 27436 4752 27488 4758
rect 27436 4694 27488 4700
rect 26936 4644 27016 4672
rect 27068 4684 27120 4690
rect 26884 4626 26936 4632
rect 27068 4626 27120 4632
rect 26516 4072 26568 4078
rect 26516 4014 26568 4020
rect 26424 4004 26476 4010
rect 26424 3946 26476 3952
rect 26436 3777 26464 3946
rect 26422 3768 26478 3777
rect 26422 3703 26478 3712
rect 26528 800 26556 4014
rect 26884 3936 26936 3942
rect 26884 3878 26936 3884
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26700 3392 26752 3398
rect 26700 3334 26752 3340
rect 26712 800 26740 3334
rect 26804 1970 26832 3538
rect 26792 1964 26844 1970
rect 26792 1906 26844 1912
rect 26896 800 26924 3878
rect 26976 2984 27028 2990
rect 26976 2926 27028 2932
rect 26988 2582 27016 2926
rect 26976 2576 27028 2582
rect 26976 2518 27028 2524
rect 27080 800 27108 4626
rect 27344 2916 27396 2922
rect 27344 2858 27396 2864
rect 27252 2508 27304 2514
rect 27252 2450 27304 2456
rect 27264 2038 27292 2450
rect 27252 2032 27304 2038
rect 27252 1974 27304 1980
rect 27356 800 27384 2858
rect 25964 332 26016 338
rect 25964 274 26016 280
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27448 513 27476 4694
rect 27528 3732 27580 3738
rect 27528 3674 27580 3680
rect 27540 800 27568 3674
rect 27632 2990 27660 31350
rect 27724 29510 27752 31826
rect 27712 29504 27764 29510
rect 27712 29446 27764 29452
rect 27816 27538 27844 33526
rect 28000 33386 28028 34342
rect 28092 34202 28120 34342
rect 28080 34196 28132 34202
rect 28080 34138 28132 34144
rect 27988 33380 28040 33386
rect 27988 33322 28040 33328
rect 27896 32360 27948 32366
rect 27896 32302 27948 32308
rect 27908 31754 27936 32302
rect 28368 31754 28396 37266
rect 28540 37188 28592 37194
rect 28540 37130 28592 37136
rect 28552 31754 28580 37130
rect 29288 36718 29316 39200
rect 30104 39160 30156 39166
rect 30104 39102 30156 39108
rect 29644 37324 29696 37330
rect 29644 37266 29696 37272
rect 29656 37126 29684 37266
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 28632 36712 28684 36718
rect 28632 36654 28684 36660
rect 29276 36712 29328 36718
rect 29276 36654 29328 36660
rect 28644 35834 28672 36654
rect 29000 36644 29052 36650
rect 29000 36586 29052 36592
rect 28724 36168 28776 36174
rect 28722 36136 28724 36145
rect 28776 36136 28778 36145
rect 28722 36071 28778 36080
rect 28632 35828 28684 35834
rect 28632 35770 28684 35776
rect 29012 35494 29040 36586
rect 29000 35488 29052 35494
rect 29000 35430 29052 35436
rect 29012 34474 29040 35430
rect 29000 34468 29052 34474
rect 29000 34410 29052 34416
rect 29368 34060 29420 34066
rect 29368 34002 29420 34008
rect 28816 33380 28868 33386
rect 28816 33322 28868 33328
rect 27908 31726 28028 31754
rect 28368 31726 28488 31754
rect 28552 31726 28764 31754
rect 27894 28248 27950 28257
rect 27894 28183 27950 28192
rect 27908 27538 27936 28183
rect 27804 27532 27856 27538
rect 27804 27474 27856 27480
rect 27896 27532 27948 27538
rect 27896 27474 27948 27480
rect 27802 26888 27858 26897
rect 27802 26823 27858 26832
rect 27712 25152 27764 25158
rect 27712 25094 27764 25100
rect 27724 24954 27752 25094
rect 27712 24948 27764 24954
rect 27712 24890 27764 24896
rect 27816 21418 27844 26823
rect 27804 21412 27856 21418
rect 27804 21354 27856 21360
rect 28000 16658 28028 31726
rect 28080 31408 28132 31414
rect 28356 31408 28408 31414
rect 28080 31350 28132 31356
rect 28354 31376 28356 31385
rect 28408 31376 28410 31385
rect 28092 31249 28120 31350
rect 28354 31311 28410 31320
rect 28078 31240 28134 31249
rect 28078 31175 28134 31184
rect 28172 31204 28224 31210
rect 28172 31146 28224 31152
rect 28184 31113 28212 31146
rect 28170 31104 28226 31113
rect 28170 31039 28226 31048
rect 28356 30864 28408 30870
rect 28354 30832 28356 30841
rect 28408 30832 28410 30841
rect 28354 30767 28410 30776
rect 28080 28756 28132 28762
rect 28080 28698 28132 28704
rect 28092 24682 28120 28698
rect 28080 24676 28132 24682
rect 28080 24618 28132 24624
rect 28356 17672 28408 17678
rect 28092 17632 28356 17660
rect 27988 16652 28040 16658
rect 27988 16594 28040 16600
rect 27712 13456 27764 13462
rect 27710 13424 27712 13433
rect 27764 13424 27766 13433
rect 27710 13359 27766 13368
rect 28000 10130 28028 16594
rect 28092 12434 28120 17632
rect 28356 17614 28408 17620
rect 28092 12406 28212 12434
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 28092 10266 28120 11698
rect 28080 10260 28132 10266
rect 28080 10202 28132 10208
rect 27988 10124 28040 10130
rect 27988 10066 28040 10072
rect 27804 5160 27856 5166
rect 27804 5102 27856 5108
rect 27816 3942 27844 5102
rect 28080 4072 28132 4078
rect 28080 4014 28132 4020
rect 27804 3936 27856 3942
rect 27804 3878 27856 3884
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 27724 800 27752 3538
rect 27896 2372 27948 2378
rect 27896 2314 27948 2320
rect 27908 800 27936 2314
rect 28092 800 28120 4014
rect 28184 2446 28212 12406
rect 28356 11552 28408 11558
rect 28356 11494 28408 11500
rect 28368 11286 28396 11494
rect 28356 11280 28408 11286
rect 28356 11222 28408 11228
rect 28460 10962 28488 31726
rect 28632 27396 28684 27402
rect 28632 27338 28684 27344
rect 28644 27130 28672 27338
rect 28632 27124 28684 27130
rect 28632 27066 28684 27072
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28368 10934 28488 10962
rect 28368 6662 28396 10934
rect 28448 10804 28500 10810
rect 28448 10746 28500 10752
rect 28460 10062 28488 10746
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28356 6656 28408 6662
rect 28356 6598 28408 6604
rect 28368 2922 28488 2938
rect 28368 2916 28500 2922
rect 28368 2910 28448 2916
rect 28172 2440 28224 2446
rect 28172 2382 28224 2388
rect 28368 800 28396 2910
rect 28448 2858 28500 2864
rect 28552 2774 28580 24006
rect 28632 17672 28684 17678
rect 28630 17640 28632 17649
rect 28684 17640 28686 17649
rect 28630 17575 28686 17584
rect 28632 13184 28684 13190
rect 28632 13126 28684 13132
rect 28644 12918 28672 13126
rect 28632 12912 28684 12918
rect 28632 12854 28684 12860
rect 28644 11762 28672 12854
rect 28736 12434 28764 31726
rect 28828 16726 28856 33322
rect 29380 32842 29408 34002
rect 29368 32836 29420 32842
rect 29368 32778 29420 32784
rect 28908 27668 28960 27674
rect 28908 27610 28960 27616
rect 29092 27668 29144 27674
rect 29092 27610 29144 27616
rect 28920 27538 28948 27610
rect 28908 27532 28960 27538
rect 28908 27474 28960 27480
rect 29000 27328 29052 27334
rect 29000 27270 29052 27276
rect 28908 27124 28960 27130
rect 28908 27066 28960 27072
rect 28920 21622 28948 27066
rect 29012 26994 29040 27270
rect 29000 26988 29052 26994
rect 29000 26930 29052 26936
rect 29104 23322 29132 27610
rect 29092 23316 29144 23322
rect 29092 23258 29144 23264
rect 29000 21956 29052 21962
rect 29000 21898 29052 21904
rect 28908 21616 28960 21622
rect 28908 21558 28960 21564
rect 29012 20942 29040 21898
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 28908 17332 28960 17338
rect 28908 17274 28960 17280
rect 28920 16726 28948 17274
rect 28816 16720 28868 16726
rect 28816 16662 28868 16668
rect 28908 16720 28960 16726
rect 28908 16662 28960 16668
rect 28736 12406 28856 12434
rect 28632 11756 28684 11762
rect 28632 11698 28684 11704
rect 28632 11008 28684 11014
rect 28632 10950 28684 10956
rect 28644 10810 28672 10950
rect 28632 10804 28684 10810
rect 28632 10746 28684 10752
rect 28632 4480 28684 4486
rect 28632 4422 28684 4428
rect 28460 2746 28580 2774
rect 28460 2582 28488 2746
rect 28644 2650 28672 4422
rect 28724 4072 28776 4078
rect 28724 4014 28776 4020
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 28448 2576 28500 2582
rect 28448 2518 28500 2524
rect 28540 2304 28592 2310
rect 28540 2246 28592 2252
rect 28552 800 28580 2246
rect 28736 800 28764 4014
rect 28828 2990 28856 12406
rect 29012 6254 29040 20878
rect 29092 20800 29144 20806
rect 29092 20742 29144 20748
rect 29104 19854 29132 20742
rect 29092 19848 29144 19854
rect 29092 19790 29144 19796
rect 29104 18057 29132 19790
rect 29090 18048 29146 18057
rect 29090 17983 29146 17992
rect 29090 17912 29146 17921
rect 29090 17847 29146 17856
rect 29104 17270 29132 17847
rect 29092 17264 29144 17270
rect 29092 17206 29144 17212
rect 29656 16250 29684 37062
rect 29828 34536 29880 34542
rect 29828 34478 29880 34484
rect 29840 32298 29868 34478
rect 30010 33416 30066 33425
rect 30010 33351 30012 33360
rect 30064 33351 30066 33360
rect 30012 33322 30064 33328
rect 29828 32292 29880 32298
rect 29828 32234 29880 32240
rect 29840 29510 29868 32234
rect 29920 32224 29972 32230
rect 29920 32166 29972 32172
rect 29828 29504 29880 29510
rect 29828 29446 29880 29452
rect 29932 26994 29960 32166
rect 30010 28656 30066 28665
rect 30010 28591 30066 28600
rect 30024 28218 30052 28591
rect 30012 28212 30064 28218
rect 30012 28154 30064 28160
rect 29920 26988 29972 26994
rect 29920 26930 29972 26936
rect 29920 23316 29972 23322
rect 29920 23258 29972 23264
rect 29932 22234 29960 23258
rect 29920 22228 29972 22234
rect 29920 22170 29972 22176
rect 29644 16244 29696 16250
rect 29644 16186 29696 16192
rect 29000 6248 29052 6254
rect 29000 6190 29052 6196
rect 29276 6248 29328 6254
rect 29276 6190 29328 6196
rect 29288 5302 29316 6190
rect 29736 5840 29788 5846
rect 29736 5782 29788 5788
rect 29276 5296 29328 5302
rect 29276 5238 29328 5244
rect 29092 4684 29144 4690
rect 29092 4626 29144 4632
rect 29104 3738 29132 4626
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 29092 3732 29144 3738
rect 29092 3674 29144 3680
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28816 2984 28868 2990
rect 28816 2926 28868 2932
rect 28920 800 28948 3538
rect 29092 2372 29144 2378
rect 29092 2314 29144 2320
rect 29104 800 29132 2314
rect 29380 800 29408 4014
rect 29552 2984 29604 2990
rect 29552 2926 29604 2932
rect 29564 800 29592 2926
rect 29748 2514 29776 5782
rect 29932 4010 29960 22170
rect 30116 20942 30144 39102
rect 30208 37466 30236 39200
rect 30564 38072 30616 38078
rect 30564 38014 30616 38020
rect 30196 37460 30248 37466
rect 30196 37402 30248 37408
rect 30288 36576 30340 36582
rect 30288 36518 30340 36524
rect 30194 33688 30250 33697
rect 30194 33623 30250 33632
rect 30208 33590 30236 33623
rect 30196 33584 30248 33590
rect 30196 33526 30248 33532
rect 30300 33454 30328 36518
rect 30472 34196 30524 34202
rect 30472 34138 30524 34144
rect 30380 34060 30432 34066
rect 30380 34002 30432 34008
rect 30196 33448 30248 33454
rect 30196 33390 30248 33396
rect 30288 33448 30340 33454
rect 30288 33390 30340 33396
rect 30208 22098 30236 33390
rect 30392 32570 30420 34002
rect 30484 33454 30512 34138
rect 30472 33448 30524 33454
rect 30472 33390 30524 33396
rect 30472 33312 30524 33318
rect 30470 33280 30472 33289
rect 30524 33280 30526 33289
rect 30470 33215 30526 33224
rect 30380 32564 30432 32570
rect 30380 32506 30432 32512
rect 30288 30388 30340 30394
rect 30288 30330 30340 30336
rect 30380 30388 30432 30394
rect 30380 30330 30432 30336
rect 30300 28422 30328 30330
rect 30392 30122 30420 30330
rect 30380 30116 30432 30122
rect 30380 30058 30432 30064
rect 30288 28416 30340 28422
rect 30288 28358 30340 28364
rect 30380 28212 30432 28218
rect 30380 28154 30432 28160
rect 30392 27538 30420 28154
rect 30380 27532 30432 27538
rect 30380 27474 30432 27480
rect 30472 27532 30524 27538
rect 30472 27474 30524 27480
rect 30484 27441 30512 27474
rect 30470 27432 30526 27441
rect 30470 27367 30526 27376
rect 30470 27024 30526 27033
rect 30288 26988 30340 26994
rect 30470 26959 30526 26968
rect 30288 26930 30340 26936
rect 30196 22092 30248 22098
rect 30196 22034 30248 22040
rect 30104 20936 30156 20942
rect 30104 20878 30156 20884
rect 30208 15570 30236 22034
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 30300 8362 30328 26930
rect 30378 26616 30434 26625
rect 30378 26551 30380 26560
rect 30432 26551 30434 26560
rect 30380 26522 30432 26528
rect 30484 26450 30512 26959
rect 30576 26586 30604 38014
rect 30932 37392 30984 37398
rect 31036 37380 31064 39200
rect 31576 38072 31628 38078
rect 31576 38014 31628 38020
rect 31208 37732 31260 37738
rect 31208 37674 31260 37680
rect 31392 37732 31444 37738
rect 31392 37674 31444 37680
rect 31220 37466 31248 37674
rect 31208 37460 31260 37466
rect 31208 37402 31260 37408
rect 31404 37398 31432 37674
rect 30984 37352 31064 37380
rect 31392 37392 31444 37398
rect 30932 37334 30984 37340
rect 31392 37334 31444 37340
rect 31484 37324 31536 37330
rect 31484 37266 31536 37272
rect 31496 34202 31524 37266
rect 31484 34196 31536 34202
rect 31484 34138 31536 34144
rect 30932 33516 30984 33522
rect 30932 33458 30984 33464
rect 30944 33425 30972 33458
rect 30930 33416 30986 33425
rect 30930 33351 30986 33360
rect 30748 33312 30800 33318
rect 30748 33254 30800 33260
rect 30656 29504 30708 29510
rect 30656 29446 30708 29452
rect 30564 26580 30616 26586
rect 30564 26522 30616 26528
rect 30472 26444 30524 26450
rect 30472 26386 30524 26392
rect 30472 25220 30524 25226
rect 30472 25162 30524 25168
rect 30380 24608 30432 24614
rect 30378 24576 30380 24585
rect 30432 24576 30434 24585
rect 30378 24511 30434 24520
rect 30380 18216 30432 18222
rect 30380 18158 30432 18164
rect 30392 16640 30420 18158
rect 30484 17678 30512 25162
rect 30472 17672 30524 17678
rect 30472 17614 30524 17620
rect 30576 16658 30604 26522
rect 30668 26450 30696 29446
rect 30656 26444 30708 26450
rect 30656 26386 30708 26392
rect 30472 16652 30524 16658
rect 30392 16612 30472 16640
rect 30472 16594 30524 16600
rect 30564 16652 30616 16658
rect 30564 16594 30616 16600
rect 30484 14482 30512 16594
rect 30472 14476 30524 14482
rect 30472 14418 30524 14424
rect 30380 12980 30432 12986
rect 30380 12922 30432 12928
rect 30392 11558 30420 12922
rect 30484 12238 30512 14418
rect 30472 12232 30524 12238
rect 30472 12174 30524 12180
rect 30668 12170 30696 26386
rect 30760 12306 30788 33254
rect 31588 31754 31616 38014
rect 31956 37398 31984 39200
rect 32588 38344 32640 38350
rect 32588 38286 32640 38292
rect 31944 37392 31996 37398
rect 31944 37334 31996 37340
rect 31668 36712 31720 36718
rect 31668 36654 31720 36660
rect 31680 36174 31708 36654
rect 31668 36168 31720 36174
rect 31668 36110 31720 36116
rect 31668 34740 31720 34746
rect 31668 34682 31720 34688
rect 31680 32570 31708 34682
rect 32496 33380 32548 33386
rect 32496 33322 32548 33328
rect 32404 32768 32456 32774
rect 32404 32710 32456 32716
rect 31668 32564 31720 32570
rect 31668 32506 31720 32512
rect 31588 31726 31708 31754
rect 31298 30696 31354 30705
rect 31298 30631 31354 30640
rect 31024 27328 31076 27334
rect 31024 27270 31076 27276
rect 30840 26852 30892 26858
rect 30840 26794 30892 26800
rect 30932 26852 30984 26858
rect 30932 26794 30984 26800
rect 30852 26586 30880 26794
rect 30840 26580 30892 26586
rect 30840 26522 30892 26528
rect 30944 26450 30972 26794
rect 31036 26450 31064 27270
rect 30932 26444 30984 26450
rect 30932 26386 30984 26392
rect 31024 26444 31076 26450
rect 31024 26386 31076 26392
rect 30932 25356 30984 25362
rect 30932 25298 30984 25304
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 30852 19174 30880 24550
rect 30840 19168 30892 19174
rect 30840 19110 30892 19116
rect 30748 12300 30800 12306
rect 30748 12242 30800 12248
rect 30656 12164 30708 12170
rect 30656 12106 30708 12112
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 30380 9988 30432 9994
rect 30380 9930 30432 9936
rect 30392 9178 30420 9930
rect 30380 9172 30432 9178
rect 30380 9114 30432 9120
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 29920 4004 29972 4010
rect 29920 3946 29972 3952
rect 29920 3596 29972 3602
rect 29920 3538 29972 3544
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 29736 2304 29788 2310
rect 29736 2246 29788 2252
rect 29748 800 29776 2246
rect 29932 800 29960 3538
rect 30104 2984 30156 2990
rect 30104 2926 30156 2932
rect 30116 800 30144 2926
rect 30300 1358 30328 8298
rect 30944 8294 30972 25298
rect 31116 18148 31168 18154
rect 31116 18090 31168 18096
rect 31024 16040 31076 16046
rect 31022 16008 31024 16017
rect 31076 16008 31078 16017
rect 31022 15943 31078 15952
rect 31024 12708 31076 12714
rect 31024 12650 31076 12656
rect 31036 12102 31064 12650
rect 31024 12096 31076 12102
rect 31024 12038 31076 12044
rect 30932 8288 30984 8294
rect 30932 8230 30984 8236
rect 31024 7540 31076 7546
rect 31024 7482 31076 7488
rect 30564 3596 30616 3602
rect 30564 3538 30616 3544
rect 30380 2372 30432 2378
rect 30380 2314 30432 2320
rect 30288 1352 30340 1358
rect 30288 1294 30340 1300
rect 30392 800 30420 2314
rect 30576 800 30604 3538
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 30760 800 30788 2926
rect 31036 2582 31064 7482
rect 31128 5574 31156 18090
rect 31208 15972 31260 15978
rect 31208 15914 31260 15920
rect 31220 15745 31248 15914
rect 31206 15736 31262 15745
rect 31206 15671 31262 15680
rect 31208 14068 31260 14074
rect 31208 14010 31260 14016
rect 31220 9994 31248 14010
rect 31208 9988 31260 9994
rect 31208 9930 31260 9936
rect 31116 5568 31168 5574
rect 31116 5510 31168 5516
rect 31208 4072 31260 4078
rect 31208 4014 31260 4020
rect 31024 2576 31076 2582
rect 31024 2518 31076 2524
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 30944 800 30972 2382
rect 31220 800 31248 4014
rect 31312 2038 31340 30631
rect 31484 18148 31536 18154
rect 31484 18090 31536 18096
rect 31390 16280 31446 16289
rect 31390 16215 31392 16224
rect 31444 16215 31446 16224
rect 31392 16186 31444 16192
rect 31390 16144 31446 16153
rect 31390 16079 31392 16088
rect 31444 16079 31446 16088
rect 31392 16050 31444 16056
rect 31496 15994 31524 18090
rect 31576 16108 31628 16114
rect 31576 16050 31628 16056
rect 31404 15978 31524 15994
rect 31392 15972 31524 15978
rect 31444 15966 31524 15972
rect 31392 15914 31444 15920
rect 31404 13802 31432 15914
rect 31482 15464 31538 15473
rect 31482 15399 31538 15408
rect 31496 15366 31524 15399
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31484 15088 31536 15094
rect 31484 15030 31536 15036
rect 31392 13796 31444 13802
rect 31392 13738 31444 13744
rect 31392 12912 31444 12918
rect 31392 12854 31444 12860
rect 31404 5234 31432 12854
rect 31392 5228 31444 5234
rect 31392 5170 31444 5176
rect 31392 2984 31444 2990
rect 31392 2926 31444 2932
rect 31300 2032 31352 2038
rect 31300 1974 31352 1980
rect 31404 800 31432 2926
rect 31496 1834 31524 15030
rect 31588 9586 31616 16050
rect 31576 9580 31628 9586
rect 31576 9522 31628 9528
rect 31680 5098 31708 31726
rect 31760 28484 31812 28490
rect 31760 28426 31812 28432
rect 31772 28121 31800 28426
rect 31758 28112 31814 28121
rect 31758 28047 31814 28056
rect 32128 28008 32180 28014
rect 32128 27950 32180 27956
rect 31852 25968 31904 25974
rect 31852 25910 31904 25916
rect 31760 17672 31812 17678
rect 31760 17614 31812 17620
rect 31772 17542 31800 17614
rect 31760 17536 31812 17542
rect 31760 17478 31812 17484
rect 31760 16448 31812 16454
rect 31758 16416 31760 16425
rect 31812 16416 31814 16425
rect 31758 16351 31814 16360
rect 31758 16280 31814 16289
rect 31758 16215 31814 16224
rect 31772 16182 31800 16215
rect 31760 16176 31812 16182
rect 31760 16118 31812 16124
rect 31758 16008 31814 16017
rect 31758 15943 31814 15952
rect 31772 15910 31800 15943
rect 31760 15904 31812 15910
rect 31760 15846 31812 15852
rect 31864 14618 31892 25910
rect 32140 25430 32168 27950
rect 32128 25424 32180 25430
rect 32128 25366 32180 25372
rect 32220 21548 32272 21554
rect 32220 21490 32272 21496
rect 31944 17536 31996 17542
rect 31944 17478 31996 17484
rect 31956 17202 31984 17478
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 32036 17196 32088 17202
rect 32036 17138 32088 17144
rect 32048 17066 32076 17138
rect 32036 17060 32088 17066
rect 32036 17002 32088 17008
rect 31944 16448 31996 16454
rect 31944 16390 31996 16396
rect 31956 15094 31984 16390
rect 32034 16144 32090 16153
rect 32034 16079 32036 16088
rect 32088 16079 32090 16088
rect 32036 16050 32088 16056
rect 32128 16040 32180 16046
rect 32128 15982 32180 15988
rect 32036 15972 32088 15978
rect 32036 15914 32088 15920
rect 32048 15745 32076 15914
rect 32034 15736 32090 15745
rect 32034 15671 32090 15680
rect 32140 15570 32168 15982
rect 32128 15564 32180 15570
rect 32128 15506 32180 15512
rect 32034 15464 32090 15473
rect 32034 15399 32090 15408
rect 32048 15366 32076 15399
rect 32036 15360 32088 15366
rect 32036 15302 32088 15308
rect 31944 15088 31996 15094
rect 31944 15030 31996 15036
rect 31852 14612 31904 14618
rect 31852 14554 31904 14560
rect 31864 8498 31892 14554
rect 32036 12232 32088 12238
rect 32036 12174 32088 12180
rect 32048 11558 32076 12174
rect 32036 11552 32088 11558
rect 32036 11494 32088 11500
rect 31852 8492 31904 8498
rect 31852 8434 31904 8440
rect 32048 7954 32076 11494
rect 32232 7954 32260 21490
rect 31852 7948 31904 7954
rect 31852 7890 31904 7896
rect 32036 7948 32088 7954
rect 32036 7890 32088 7896
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 31864 7342 31892 7890
rect 31852 7336 31904 7342
rect 31852 7278 31904 7284
rect 32416 5778 32444 32710
rect 32508 22273 32536 33322
rect 32600 32774 32628 38286
rect 32784 37466 32812 39200
rect 32864 39092 32916 39098
rect 32864 39034 32916 39040
rect 32772 37460 32824 37466
rect 32772 37402 32824 37408
rect 32876 37210 32904 39034
rect 32784 37182 32904 37210
rect 32588 32768 32640 32774
rect 32588 32710 32640 32716
rect 32494 22264 32550 22273
rect 32494 22199 32550 22208
rect 32508 18154 32536 22199
rect 32496 18148 32548 18154
rect 32496 18090 32548 18096
rect 32600 17218 32628 32710
rect 32680 27464 32732 27470
rect 32680 27406 32732 27412
rect 32692 17354 32720 27406
rect 32784 17490 32812 37182
rect 32864 37120 32916 37126
rect 32864 37062 32916 37068
rect 32876 21622 32904 37062
rect 33704 36854 33732 39200
rect 34532 37398 34560 39200
rect 34704 37800 34756 37806
rect 34704 37742 34756 37748
rect 34716 37466 34744 37742
rect 35452 37466 35480 39200
rect 36176 37664 36228 37670
rect 36176 37606 36228 37612
rect 34704 37460 34756 37466
rect 34704 37402 34756 37408
rect 35440 37460 35492 37466
rect 35440 37402 35492 37408
rect 34520 37392 34572 37398
rect 34520 37334 34572 37340
rect 34060 37324 34112 37330
rect 34060 37266 34112 37272
rect 36084 37324 36136 37330
rect 36084 37266 36136 37272
rect 33692 36848 33744 36854
rect 33692 36790 33744 36796
rect 33968 36644 34020 36650
rect 33968 36586 34020 36592
rect 33416 36304 33468 36310
rect 33416 36246 33468 36252
rect 33428 36038 33456 36246
rect 33692 36236 33744 36242
rect 33520 36196 33692 36224
rect 33324 36032 33376 36038
rect 33324 35974 33376 35980
rect 33416 36032 33468 36038
rect 33416 35974 33468 35980
rect 33336 35894 33364 35974
rect 33520 35894 33548 36196
rect 33692 36178 33744 36184
rect 33336 35866 33548 35894
rect 33508 35828 33560 35834
rect 33508 35770 33560 35776
rect 33520 35714 33548 35770
rect 33876 35760 33928 35766
rect 33520 35708 33876 35714
rect 33520 35702 33928 35708
rect 33520 35686 33916 35702
rect 33980 34626 34008 36586
rect 33796 34598 34008 34626
rect 33692 32292 33744 32298
rect 33692 32234 33744 32240
rect 33704 31890 33732 32234
rect 33692 31884 33744 31890
rect 33692 31826 33744 31832
rect 33232 30184 33284 30190
rect 33232 30126 33284 30132
rect 33140 28008 33192 28014
rect 33140 27950 33192 27956
rect 33152 23186 33180 27950
rect 33140 23180 33192 23186
rect 33140 23122 33192 23128
rect 33140 22976 33192 22982
rect 33140 22918 33192 22924
rect 33048 22160 33100 22166
rect 33046 22128 33048 22137
rect 33100 22128 33102 22137
rect 33046 22063 33102 22072
rect 32864 21616 32916 21622
rect 32864 21558 32916 21564
rect 33046 18320 33102 18329
rect 33046 18255 33102 18264
rect 33060 18154 33088 18255
rect 33048 18148 33100 18154
rect 33048 18090 33100 18096
rect 32784 17462 32996 17490
rect 32692 17326 32812 17354
rect 32600 17190 32720 17218
rect 32496 16176 32548 16182
rect 32496 16118 32548 16124
rect 32508 14006 32536 16118
rect 32588 15088 32640 15094
rect 32588 15030 32640 15036
rect 32496 14000 32548 14006
rect 32496 13942 32548 13948
rect 32496 12096 32548 12102
rect 32496 12038 32548 12044
rect 32404 5772 32456 5778
rect 32404 5714 32456 5720
rect 31668 5092 31720 5098
rect 31668 5034 31720 5040
rect 31944 3596 31996 3602
rect 31944 3538 31996 3544
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 31760 2508 31812 2514
rect 31760 2450 31812 2456
rect 31576 2304 31628 2310
rect 31772 2258 31800 2450
rect 31576 2246 31628 2252
rect 31484 1828 31536 1834
rect 31484 1770 31536 1776
rect 31588 800 31616 2246
rect 31680 2230 31800 2258
rect 31680 2038 31708 2230
rect 31760 2100 31812 2106
rect 31760 2042 31812 2048
rect 31668 2032 31720 2038
rect 31668 1974 31720 1980
rect 31772 1358 31800 2042
rect 31760 1352 31812 1358
rect 31760 1294 31812 1300
rect 31864 1204 31892 3470
rect 31772 1176 31892 1204
rect 31772 800 31800 1176
rect 31956 800 31984 3538
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 32232 800 32260 2314
rect 32416 800 32444 3334
rect 32508 2582 32536 12038
rect 32600 7478 32628 15030
rect 32692 7886 32720 17190
rect 32784 16250 32812 17326
rect 32772 16244 32824 16250
rect 32772 16186 32824 16192
rect 32772 10736 32824 10742
rect 32772 10678 32824 10684
rect 32784 10266 32812 10678
rect 32772 10260 32824 10266
rect 32772 10202 32824 10208
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 32588 7472 32640 7478
rect 32588 7414 32640 7420
rect 32968 4826 32996 17462
rect 33152 14958 33180 22918
rect 33244 14958 33272 30126
rect 33416 29096 33468 29102
rect 33416 29038 33468 29044
rect 33324 27600 33376 27606
rect 33324 27542 33376 27548
rect 33336 26761 33364 27542
rect 33322 26752 33378 26761
rect 33322 26687 33378 26696
rect 33428 26586 33456 29038
rect 33508 28620 33560 28626
rect 33508 28562 33560 28568
rect 33520 27674 33548 28562
rect 33600 27940 33652 27946
rect 33600 27882 33652 27888
rect 33612 27849 33640 27882
rect 33598 27840 33654 27849
rect 33598 27775 33654 27784
rect 33508 27668 33560 27674
rect 33508 27610 33560 27616
rect 33416 26580 33468 26586
rect 33416 26522 33468 26528
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 33140 14952 33192 14958
rect 33140 14894 33192 14900
rect 33232 14952 33284 14958
rect 33232 14894 33284 14900
rect 33232 10600 33284 10606
rect 33232 10542 33284 10548
rect 33244 10169 33272 10542
rect 33230 10160 33286 10169
rect 33230 10095 33286 10104
rect 33336 8090 33364 26386
rect 33428 22710 33456 26522
rect 33692 26512 33744 26518
rect 33690 26480 33692 26489
rect 33744 26480 33746 26489
rect 33690 26415 33746 26424
rect 33692 26376 33744 26382
rect 33690 26344 33692 26353
rect 33744 26344 33746 26353
rect 33690 26279 33746 26288
rect 33416 22704 33468 22710
rect 33416 22646 33468 22652
rect 33598 22672 33654 22681
rect 33598 22607 33600 22616
rect 33652 22607 33654 22616
rect 33600 22578 33652 22584
rect 33416 22432 33468 22438
rect 33416 22374 33468 22380
rect 33428 22234 33456 22374
rect 33416 22228 33468 22234
rect 33416 22170 33468 22176
rect 33796 21418 33824 34598
rect 33874 34504 33930 34513
rect 33874 34439 33930 34448
rect 33888 34406 33916 34439
rect 33876 34400 33928 34406
rect 33876 34342 33928 34348
rect 33968 34400 34020 34406
rect 33968 34342 34020 34348
rect 33980 33998 34008 34342
rect 33968 33992 34020 33998
rect 33968 33934 34020 33940
rect 33876 32224 33928 32230
rect 33876 32166 33928 32172
rect 33888 31890 33916 32166
rect 33876 31884 33928 31890
rect 33876 31826 33928 31832
rect 33968 31884 34020 31890
rect 33968 31826 34020 31832
rect 33980 31686 34008 31826
rect 33968 31680 34020 31686
rect 33968 31622 34020 31628
rect 33874 30832 33930 30841
rect 33874 30767 33930 30776
rect 33888 30734 33916 30767
rect 33980 30734 34008 31622
rect 33876 30728 33928 30734
rect 33876 30670 33928 30676
rect 33968 30728 34020 30734
rect 33968 30670 34020 30676
rect 34072 28994 34100 37266
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34152 36304 34204 36310
rect 34152 36246 34204 36252
rect 34164 34542 34192 36246
rect 35256 36100 35308 36106
rect 35256 36042 35308 36048
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34152 34536 34204 34542
rect 34152 34478 34204 34484
rect 34520 34536 34572 34542
rect 34520 34478 34572 34484
rect 34152 33992 34204 33998
rect 34152 33934 34204 33940
rect 34164 33658 34192 33934
rect 34242 33688 34298 33697
rect 34152 33652 34204 33658
rect 34242 33623 34244 33632
rect 34152 33594 34204 33600
rect 34296 33623 34298 33632
rect 34244 33594 34296 33600
rect 34428 29640 34480 29646
rect 34428 29582 34480 29588
rect 33980 28966 34100 28994
rect 33876 28416 33928 28422
rect 33876 28358 33928 28364
rect 33888 27334 33916 28358
rect 33876 27328 33928 27334
rect 33876 27270 33928 27276
rect 33874 22672 33930 22681
rect 33874 22607 33876 22616
rect 33928 22607 33930 22616
rect 33876 22578 33928 22584
rect 33980 22409 34008 28966
rect 34336 27600 34388 27606
rect 34336 27542 34388 27548
rect 34348 26450 34376 27542
rect 34336 26444 34388 26450
rect 34336 26386 34388 26392
rect 34244 24676 34296 24682
rect 34244 24618 34296 24624
rect 33966 22400 34022 22409
rect 33966 22335 34022 22344
rect 33784 21412 33836 21418
rect 33784 21354 33836 21360
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33704 20369 33732 20402
rect 33690 20360 33746 20369
rect 33690 20295 33746 20304
rect 33690 20088 33746 20097
rect 33690 20023 33746 20032
rect 33704 19990 33732 20023
rect 33692 19984 33744 19990
rect 33692 19926 33744 19932
rect 33690 19408 33746 19417
rect 33690 19343 33692 19352
rect 33744 19343 33746 19352
rect 33692 19314 33744 19320
rect 33598 18864 33654 18873
rect 33598 18799 33600 18808
rect 33652 18799 33654 18808
rect 33692 18828 33744 18834
rect 33600 18770 33652 18776
rect 33692 18770 33744 18776
rect 33414 18728 33470 18737
rect 33414 18663 33470 18672
rect 33428 18086 33456 18663
rect 33506 18456 33562 18465
rect 33506 18391 33562 18400
rect 33600 18420 33652 18426
rect 33520 18290 33548 18391
rect 33600 18362 33652 18368
rect 33612 18329 33640 18362
rect 33704 18358 33732 18770
rect 33692 18352 33744 18358
rect 33598 18320 33654 18329
rect 33508 18284 33560 18290
rect 33692 18294 33744 18300
rect 33598 18255 33654 18264
rect 33508 18226 33560 18232
rect 33416 18080 33468 18086
rect 33416 18022 33468 18028
rect 33506 17232 33562 17241
rect 33506 17167 33562 17176
rect 33416 10600 33468 10606
rect 33416 10542 33468 10548
rect 33428 10062 33456 10542
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33416 8628 33468 8634
rect 33416 8570 33468 8576
rect 33428 8430 33456 8570
rect 33416 8424 33468 8430
rect 33416 8366 33468 8372
rect 33324 8084 33376 8090
rect 33324 8026 33376 8032
rect 33048 7880 33100 7886
rect 33048 7822 33100 7828
rect 32956 4820 33008 4826
rect 32956 4762 33008 4768
rect 32968 4690 32996 4762
rect 32956 4684 33008 4690
rect 32956 4626 33008 4632
rect 33060 4486 33088 7822
rect 33520 5166 33548 17167
rect 33692 15020 33744 15026
rect 33692 14962 33744 14968
rect 33704 14929 33732 14962
rect 33690 14920 33746 14929
rect 33690 14855 33746 14864
rect 33796 13394 33824 21354
rect 33980 19334 34008 22335
rect 34060 21616 34112 21622
rect 34060 21558 34112 21564
rect 34072 20330 34100 21558
rect 34060 20324 34112 20330
rect 34060 20266 34112 20272
rect 34152 20256 34204 20262
rect 34152 20198 34204 20204
rect 34164 20058 34192 20198
rect 34060 20052 34112 20058
rect 34060 19994 34112 20000
rect 34152 20052 34204 20058
rect 34152 19994 34204 20000
rect 34072 19961 34100 19994
rect 34058 19952 34114 19961
rect 34058 19887 34114 19896
rect 33888 19306 34008 19334
rect 33784 13388 33836 13394
rect 33784 13330 33836 13336
rect 33692 8832 33744 8838
rect 33692 8774 33744 8780
rect 33704 8430 33732 8774
rect 33692 8424 33744 8430
rect 33692 8366 33744 8372
rect 33692 8084 33744 8090
rect 33692 8026 33744 8032
rect 33508 5160 33560 5166
rect 33508 5102 33560 5108
rect 33324 4820 33376 4826
rect 33324 4762 33376 4768
rect 33048 4480 33100 4486
rect 33048 4422 33100 4428
rect 33140 4208 33192 4214
rect 33140 4150 33192 4156
rect 32956 4072 33008 4078
rect 32956 4014 33008 4020
rect 32864 3596 32916 3602
rect 32864 3538 32916 3544
rect 32876 3398 32904 3538
rect 32864 3392 32916 3398
rect 32864 3334 32916 3340
rect 32588 2984 32640 2990
rect 32588 2926 32640 2932
rect 32496 2576 32548 2582
rect 32496 2518 32548 2524
rect 32600 800 32628 2926
rect 32772 1420 32824 1426
rect 32772 1362 32824 1368
rect 32784 800 32812 1362
rect 32968 800 32996 4014
rect 33152 2650 33180 4150
rect 33232 2984 33284 2990
rect 33232 2926 33284 2932
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 33048 2032 33100 2038
rect 33048 1974 33100 1980
rect 27434 504 27490 513
rect 27434 439 27490 448
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33060 649 33088 1974
rect 33244 800 33272 2926
rect 33336 1766 33364 4762
rect 33508 4276 33560 4282
rect 33508 4218 33560 4224
rect 33416 2644 33468 2650
rect 33416 2586 33468 2592
rect 33324 1760 33376 1766
rect 33324 1702 33376 1708
rect 33428 800 33456 2586
rect 33520 1902 33548 4218
rect 33600 4072 33652 4078
rect 33600 4014 33652 4020
rect 33508 1896 33560 1902
rect 33508 1838 33560 1844
rect 33612 800 33640 4014
rect 33704 2582 33732 8026
rect 33888 6798 33916 19306
rect 34256 19009 34284 24618
rect 34440 23730 34468 29582
rect 34428 23724 34480 23730
rect 34428 23666 34480 23672
rect 34336 23588 34388 23594
rect 34336 23530 34388 23536
rect 34242 19000 34298 19009
rect 34242 18935 34298 18944
rect 34150 18456 34206 18465
rect 34150 18391 34206 18400
rect 34164 18290 34192 18391
rect 34152 18284 34204 18290
rect 34152 18226 34204 18232
rect 34256 17626 34284 18935
rect 34164 17598 34284 17626
rect 33968 17264 34020 17270
rect 33968 17206 34020 17212
rect 33980 14074 34008 17206
rect 34164 16538 34192 17598
rect 34244 16992 34296 16998
rect 34244 16934 34296 16940
rect 34256 16658 34284 16934
rect 34244 16652 34296 16658
rect 34244 16594 34296 16600
rect 34164 16510 34284 16538
rect 34060 16176 34112 16182
rect 34058 16144 34060 16153
rect 34112 16144 34114 16153
rect 34058 16079 34114 16088
rect 33968 14068 34020 14074
rect 33968 14010 34020 14016
rect 33980 12434 34008 14010
rect 33980 12406 34192 12434
rect 33968 10124 34020 10130
rect 33968 10066 34020 10072
rect 33980 9926 34008 10066
rect 33968 9920 34020 9926
rect 33968 9862 34020 9868
rect 33980 8838 34008 9862
rect 33968 8832 34020 8838
rect 33968 8774 34020 8780
rect 33876 6792 33928 6798
rect 33876 6734 33928 6740
rect 33876 6180 33928 6186
rect 33876 6122 33928 6128
rect 33784 2984 33836 2990
rect 33784 2926 33836 2932
rect 33692 2576 33744 2582
rect 33692 2518 33744 2524
rect 33796 800 33824 2926
rect 33888 950 33916 6122
rect 34060 5568 34112 5574
rect 34060 5510 34112 5516
rect 34072 2582 34100 5510
rect 34164 5166 34192 12406
rect 34256 8242 34284 16510
rect 34348 8498 34376 23530
rect 34426 19136 34482 19145
rect 34426 19071 34482 19080
rect 34440 18222 34468 19071
rect 34428 18216 34480 18222
rect 34428 18158 34480 18164
rect 34428 17128 34480 17134
rect 34426 17096 34428 17105
rect 34480 17096 34482 17105
rect 34426 17031 34482 17040
rect 34336 8492 34388 8498
rect 34336 8434 34388 8440
rect 34532 8378 34560 34478
rect 35268 34202 35296 36042
rect 35992 35556 36044 35562
rect 35992 35498 36044 35504
rect 36004 35465 36032 35498
rect 35990 35456 36046 35465
rect 35990 35391 36046 35400
rect 34796 34196 34848 34202
rect 34796 34138 34848 34144
rect 35256 34196 35308 34202
rect 35256 34138 35308 34144
rect 34808 33318 34836 34138
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34796 33312 34848 33318
rect 34796 33254 34848 33260
rect 35440 32904 35492 32910
rect 35440 32846 35492 32852
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 35348 30728 35400 30734
rect 35348 30670 35400 30676
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 34796 28008 34848 28014
rect 34796 27950 34848 27956
rect 34612 25696 34664 25702
rect 34612 25638 34664 25644
rect 34624 8498 34652 25638
rect 34808 21554 34836 27950
rect 35256 27464 35308 27470
rect 35256 27406 35308 27412
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 35268 27130 35296 27406
rect 35256 27124 35308 27130
rect 35256 27066 35308 27072
rect 35268 26586 35296 27066
rect 35256 26580 35308 26586
rect 35256 26522 35308 26528
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35256 22432 35308 22438
rect 35256 22374 35308 22380
rect 35268 22234 35296 22374
rect 35256 22228 35308 22234
rect 35256 22170 35308 22176
rect 35360 22094 35388 30670
rect 35268 22066 35388 22094
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 35268 21350 35296 22066
rect 35348 21548 35400 21554
rect 35348 21490 35400 21496
rect 35256 21344 35308 21350
rect 35256 21286 35308 21292
rect 35256 20936 35308 20942
rect 35256 20878 35308 20884
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34702 20360 34758 20369
rect 34702 20295 34704 20304
rect 34756 20295 34758 20304
rect 34704 20266 34756 20272
rect 34796 19712 34848 19718
rect 34796 19654 34848 19660
rect 34808 19446 34836 19654
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 34796 19440 34848 19446
rect 34796 19382 34848 19388
rect 34888 19440 34940 19446
rect 34888 19382 34940 19388
rect 34900 19334 34928 19382
rect 34808 19306 34928 19334
rect 34704 19236 34756 19242
rect 34704 19178 34756 19184
rect 34716 19145 34744 19178
rect 34702 19136 34758 19145
rect 34702 19071 34758 19080
rect 34808 17134 34836 19306
rect 35268 18834 35296 20878
rect 35256 18828 35308 18834
rect 35256 18770 35308 18776
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 35268 18358 35296 18770
rect 35360 18426 35388 21490
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 35256 18352 35308 18358
rect 35162 18320 35218 18329
rect 35256 18294 35308 18300
rect 35346 18320 35402 18329
rect 35162 18255 35218 18264
rect 35346 18255 35402 18264
rect 35176 18086 35204 18255
rect 35164 18080 35216 18086
rect 35164 18022 35216 18028
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35164 17264 35216 17270
rect 35162 17232 35164 17241
rect 35216 17232 35218 17241
rect 35162 17167 35218 17176
rect 34796 17128 34848 17134
rect 35256 17128 35308 17134
rect 34796 17070 34848 17076
rect 35084 17076 35256 17082
rect 35084 17070 35308 17076
rect 34702 16416 34758 16425
rect 34702 16351 34758 16360
rect 34716 16046 34744 16351
rect 34704 16040 34756 16046
rect 34704 15982 34756 15988
rect 34704 14612 34756 14618
rect 34704 14554 34756 14560
rect 34612 8492 34664 8498
rect 34612 8434 34664 8440
rect 34428 8356 34480 8362
rect 34532 8350 34652 8378
rect 34428 8298 34480 8304
rect 34440 8242 34468 8298
rect 34256 8214 34376 8242
rect 34440 8214 34560 8242
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 34256 7002 34284 7346
rect 34244 6996 34296 7002
rect 34244 6938 34296 6944
rect 34152 5160 34204 5166
rect 34152 5102 34204 5108
rect 34244 4684 34296 4690
rect 34244 4626 34296 4632
rect 34060 2576 34112 2582
rect 34060 2518 34112 2524
rect 33968 2304 34020 2310
rect 33968 2246 34020 2252
rect 33980 1426 34008 2246
rect 33968 1420 34020 1426
rect 33968 1362 34020 1368
rect 34060 1420 34112 1426
rect 34060 1362 34112 1368
rect 34072 1204 34100 1362
rect 33980 1176 34100 1204
rect 33876 944 33928 950
rect 33876 886 33928 892
rect 33980 800 34008 1176
rect 34256 800 34284 4626
rect 34348 4078 34376 8214
rect 34428 6928 34480 6934
rect 34428 6870 34480 6876
rect 34440 6254 34468 6870
rect 34428 6248 34480 6254
rect 34428 6190 34480 6196
rect 34336 4072 34388 4078
rect 34336 4014 34388 4020
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34440 800 34468 3538
rect 34532 814 34560 8214
rect 34624 5302 34652 8350
rect 34716 7478 34744 14554
rect 34808 11529 34836 17070
rect 35084 17054 35296 17070
rect 35084 16998 35112 17054
rect 35072 16992 35124 16998
rect 35072 16934 35124 16940
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35360 15366 35388 18255
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35256 14340 35308 14346
rect 35256 14282 35308 14288
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34794 11520 34850 11529
rect 34794 11455 34850 11464
rect 34704 7472 34756 7478
rect 34704 7414 34756 7420
rect 34808 5710 34836 11455
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34796 5704 34848 5710
rect 34796 5646 34848 5652
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34612 5296 34664 5302
rect 34612 5238 34664 5244
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34796 4072 34848 4078
rect 34796 4014 34848 4020
rect 34704 3732 34756 3738
rect 34704 3674 34756 3680
rect 34716 3058 34744 3674
rect 34704 3052 34756 3058
rect 34704 2994 34756 3000
rect 34612 2916 34664 2922
rect 34612 2858 34664 2864
rect 34520 808 34572 814
rect 33046 640 33102 649
rect 33046 575 33102 584
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34624 800 34652 2858
rect 34704 2372 34756 2378
rect 34704 2314 34756 2320
rect 34716 1426 34744 2314
rect 34704 1420 34756 1426
rect 34704 1362 34756 1368
rect 34808 800 34836 4014
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35268 2582 35296 14282
rect 35360 12481 35388 15302
rect 35346 12472 35402 12481
rect 35346 12407 35402 12416
rect 35348 12368 35400 12374
rect 35348 12310 35400 12316
rect 35360 2990 35388 12310
rect 35452 6798 35480 32846
rect 35624 30116 35676 30122
rect 35624 30058 35676 30064
rect 35532 29640 35584 29646
rect 35532 29582 35584 29588
rect 35544 23866 35572 29582
rect 35636 29102 35664 30058
rect 35716 29572 35768 29578
rect 35716 29514 35768 29520
rect 35728 29481 35756 29514
rect 35714 29472 35770 29481
rect 35714 29407 35770 29416
rect 35624 29096 35676 29102
rect 35624 29038 35676 29044
rect 35900 27600 35952 27606
rect 35898 27568 35900 27577
rect 35992 27600 36044 27606
rect 35952 27568 35954 27577
rect 35992 27542 36044 27548
rect 35898 27503 35954 27512
rect 36004 26926 36032 27542
rect 35992 26920 36044 26926
rect 36096 26897 36124 37266
rect 36188 28257 36216 37606
rect 36280 36854 36308 39200
rect 36636 38616 36688 38622
rect 36636 38558 36688 38564
rect 36648 37330 36676 38558
rect 37096 37800 37148 37806
rect 37096 37742 37148 37748
rect 36636 37324 36688 37330
rect 36636 37266 36688 37272
rect 36268 36848 36320 36854
rect 36268 36790 36320 36796
rect 36636 36848 36688 36854
rect 36636 36790 36688 36796
rect 36648 36718 36676 36790
rect 36636 36712 36688 36718
rect 36636 36654 36688 36660
rect 36728 36712 36780 36718
rect 36728 36654 36780 36660
rect 36268 36644 36320 36650
rect 36268 36586 36320 36592
rect 36280 33300 36308 36586
rect 36740 36242 36768 36654
rect 36728 36236 36780 36242
rect 36728 36178 36780 36184
rect 36360 35556 36412 35562
rect 36360 35498 36412 35504
rect 36372 35222 36400 35498
rect 36452 35488 36504 35494
rect 36452 35430 36504 35436
rect 36544 35488 36596 35494
rect 36544 35430 36596 35436
rect 36464 35222 36492 35430
rect 36360 35216 36412 35222
rect 36360 35158 36412 35164
rect 36452 35216 36504 35222
rect 36452 35158 36504 35164
rect 36556 35034 36584 35430
rect 36464 35006 36584 35034
rect 36464 34678 36492 35006
rect 36452 34672 36504 34678
rect 36452 34614 36504 34620
rect 36372 34202 36676 34218
rect 36360 34196 36676 34202
rect 36412 34190 36676 34196
rect 36360 34138 36412 34144
rect 36544 34128 36596 34134
rect 36544 34070 36596 34076
rect 36452 34060 36504 34066
rect 36452 34002 36504 34008
rect 36464 33454 36492 34002
rect 36556 33930 36584 34070
rect 36648 34066 36676 34190
rect 36636 34060 36688 34066
rect 36636 34002 36688 34008
rect 36544 33924 36596 33930
rect 36544 33866 36596 33872
rect 36452 33448 36504 33454
rect 36452 33390 36504 33396
rect 36280 33272 36676 33300
rect 36648 32366 36676 33272
rect 36636 32360 36688 32366
rect 36636 32302 36688 32308
rect 36268 31748 36320 31754
rect 36268 31690 36320 31696
rect 36280 30841 36308 31690
rect 36648 30870 36676 32302
rect 36740 31754 36768 36178
rect 36820 35148 36872 35154
rect 36820 35090 36872 35096
rect 36912 35148 36964 35154
rect 36912 35090 36964 35096
rect 36832 34746 36860 35090
rect 36820 34740 36872 34746
rect 36820 34682 36872 34688
rect 36924 34542 36952 35090
rect 36912 34536 36964 34542
rect 36912 34478 36964 34484
rect 37004 32224 37056 32230
rect 37004 32166 37056 32172
rect 36740 31726 36860 31754
rect 36636 30864 36688 30870
rect 36266 30832 36322 30841
rect 36636 30806 36688 30812
rect 36266 30767 36322 30776
rect 36544 30796 36596 30802
rect 36174 28248 36230 28257
rect 36174 28183 36230 28192
rect 36188 26994 36216 28183
rect 36176 26988 36228 26994
rect 36176 26930 36228 26936
rect 35992 26862 36044 26868
rect 36082 26888 36138 26897
rect 36082 26823 36138 26832
rect 35808 26444 35860 26450
rect 35808 26386 35860 26392
rect 35992 26444 36044 26450
rect 35992 26386 36044 26392
rect 35820 26330 35848 26386
rect 35820 26302 35940 26330
rect 35806 25800 35862 25809
rect 35806 25735 35862 25744
rect 35820 25702 35848 25735
rect 35808 25696 35860 25702
rect 35808 25638 35860 25644
rect 35532 23860 35584 23866
rect 35532 23802 35584 23808
rect 35808 23860 35860 23866
rect 35808 23802 35860 23808
rect 35544 14958 35572 23802
rect 35624 23180 35676 23186
rect 35624 23122 35676 23128
rect 35636 16658 35664 23122
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 35624 16652 35676 16658
rect 35624 16594 35676 16600
rect 35532 14952 35584 14958
rect 35532 14894 35584 14900
rect 35530 12336 35586 12345
rect 35530 12271 35586 12280
rect 35440 6792 35492 6798
rect 35440 6734 35492 6740
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 35348 2984 35400 2990
rect 35348 2926 35400 2932
rect 35256 2576 35308 2582
rect 35256 2518 35308 2524
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35452 1850 35480 3538
rect 35544 3058 35572 12271
rect 35636 4146 35664 16594
rect 35728 16574 35756 21286
rect 35820 19242 35848 23802
rect 35912 20806 35940 26302
rect 36004 25702 36032 26386
rect 36096 26382 36124 26823
rect 36084 26376 36136 26382
rect 36084 26318 36136 26324
rect 35992 25696 36044 25702
rect 35992 25638 36044 25644
rect 35992 24812 36044 24818
rect 35992 24754 36044 24760
rect 36004 24070 36032 24754
rect 35992 24064 36044 24070
rect 35992 24006 36044 24012
rect 35992 23316 36044 23322
rect 35992 23258 36044 23264
rect 35900 20800 35952 20806
rect 35900 20742 35952 20748
rect 35900 19304 35952 19310
rect 35900 19246 35952 19252
rect 35808 19236 35860 19242
rect 35808 19178 35860 19184
rect 35808 18964 35860 18970
rect 35808 18906 35860 18912
rect 35820 18834 35848 18906
rect 35808 18828 35860 18834
rect 35808 18770 35860 18776
rect 35912 18426 35940 19246
rect 35900 18420 35952 18426
rect 35900 18362 35952 18368
rect 35808 18352 35860 18358
rect 35808 18294 35860 18300
rect 35820 16726 35848 18294
rect 35900 17196 35952 17202
rect 35900 17138 35952 17144
rect 35912 17105 35940 17138
rect 35898 17096 35954 17105
rect 35898 17031 35954 17040
rect 35808 16720 35860 16726
rect 35808 16662 35860 16668
rect 35900 16720 35952 16726
rect 35900 16662 35952 16668
rect 35912 16574 35940 16662
rect 35728 16546 35940 16574
rect 35728 9042 35756 16546
rect 35808 16176 35860 16182
rect 35808 16118 35860 16124
rect 35820 14958 35848 16118
rect 36004 14958 36032 23258
rect 36280 22094 36308 30767
rect 36544 30738 36596 30744
rect 36360 30116 36412 30122
rect 36360 30058 36412 30064
rect 36372 29578 36400 30058
rect 36360 29572 36412 29578
rect 36360 29514 36412 29520
rect 36358 27024 36414 27033
rect 36358 26959 36414 26968
rect 36372 26858 36400 26959
rect 36360 26852 36412 26858
rect 36360 26794 36412 26800
rect 36450 26616 36506 26625
rect 36450 26551 36506 26560
rect 36464 26450 36492 26551
rect 36360 26444 36412 26450
rect 36360 26386 36412 26392
rect 36452 26444 36504 26450
rect 36452 26386 36504 26392
rect 36188 22066 36308 22094
rect 36084 19304 36136 19310
rect 36082 19272 36084 19281
rect 36136 19272 36138 19281
rect 36082 19207 36138 19216
rect 36096 18358 36124 19207
rect 36084 18352 36136 18358
rect 36084 18294 36136 18300
rect 36084 15700 36136 15706
rect 36084 15642 36136 15648
rect 36096 15502 36124 15642
rect 36084 15496 36136 15502
rect 36084 15438 36136 15444
rect 35808 14952 35860 14958
rect 35808 14894 35860 14900
rect 35992 14952 36044 14958
rect 35992 14894 36044 14900
rect 35820 14618 35848 14894
rect 35808 14612 35860 14618
rect 35808 14554 35860 14560
rect 36188 12434 36216 22066
rect 36268 19780 36320 19786
rect 36268 19722 36320 19728
rect 36280 19446 36308 19722
rect 36268 19440 36320 19446
rect 36268 19382 36320 19388
rect 36372 19394 36400 26386
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 36464 23730 36492 24006
rect 36452 23724 36504 23730
rect 36452 23666 36504 23672
rect 36556 23322 36584 30738
rect 36728 30728 36780 30734
rect 36728 30670 36780 30676
rect 36740 29034 36768 30670
rect 36728 29028 36780 29034
rect 36728 28970 36780 28976
rect 36636 26988 36688 26994
rect 36636 26930 36688 26936
rect 36544 23316 36596 23322
rect 36544 23258 36596 23264
rect 36452 22704 36504 22710
rect 36452 22646 36504 22652
rect 36464 22166 36492 22646
rect 36452 22160 36504 22166
rect 36452 22102 36504 22108
rect 36648 22094 36676 26930
rect 36728 26512 36780 26518
rect 36726 26480 36728 26489
rect 36780 26480 36782 26489
rect 36726 26415 36782 26424
rect 36728 26376 36780 26382
rect 36726 26344 36728 26353
rect 36780 26344 36782 26353
rect 36726 26279 36782 26288
rect 36556 22066 36676 22094
rect 36372 19366 36492 19394
rect 36360 19304 36412 19310
rect 36360 19246 36412 19252
rect 36372 17338 36400 19246
rect 36464 18850 36492 19366
rect 36556 19310 36584 22066
rect 36634 19408 36690 19417
rect 36634 19343 36636 19352
rect 36688 19343 36690 19352
rect 36636 19314 36688 19320
rect 36544 19304 36596 19310
rect 36544 19246 36596 19252
rect 36726 19272 36782 19281
rect 36726 19207 36728 19216
rect 36780 19207 36782 19216
rect 36728 19178 36780 19184
rect 36636 19168 36688 19174
rect 36636 19110 36688 19116
rect 36726 19136 36782 19145
rect 36464 18822 36584 18850
rect 36452 18760 36504 18766
rect 36452 18702 36504 18708
rect 36464 18358 36492 18702
rect 36452 18352 36504 18358
rect 36452 18294 36504 18300
rect 36360 17332 36412 17338
rect 36360 17274 36412 17280
rect 36268 16516 36320 16522
rect 36268 16458 36320 16464
rect 36280 15706 36308 16458
rect 36268 15700 36320 15706
rect 36268 15642 36320 15648
rect 36268 15020 36320 15026
rect 36268 14962 36320 14968
rect 36280 14929 36308 14962
rect 36266 14920 36322 14929
rect 36266 14855 36322 14864
rect 36188 12406 36308 12434
rect 35900 12300 35952 12306
rect 35900 12242 35952 12248
rect 35808 11008 35860 11014
rect 35808 10950 35860 10956
rect 35820 9586 35848 10950
rect 35808 9580 35860 9586
rect 35808 9522 35860 9528
rect 35716 9036 35768 9042
rect 35716 8978 35768 8984
rect 35728 8430 35756 8978
rect 35912 8974 35940 12242
rect 35990 9616 36046 9625
rect 35990 9551 36046 9560
rect 36004 9518 36032 9551
rect 36280 9518 36308 12406
rect 36372 11762 36400 17274
rect 36556 14958 36584 18822
rect 36648 18737 36676 19110
rect 36726 19071 36782 19080
rect 36740 18970 36768 19071
rect 36728 18964 36780 18970
rect 36728 18906 36780 18912
rect 36728 18828 36780 18834
rect 36728 18770 36780 18776
rect 36634 18728 36690 18737
rect 36634 18663 36690 18672
rect 36740 18057 36768 18770
rect 36726 18048 36782 18057
rect 36726 17983 36782 17992
rect 36544 14952 36596 14958
rect 36544 14894 36596 14900
rect 36556 12434 36584 14894
rect 36728 13388 36780 13394
rect 36728 13330 36780 13336
rect 36740 13190 36768 13330
rect 36728 13184 36780 13190
rect 36728 13126 36780 13132
rect 36556 12406 36676 12434
rect 36452 12300 36504 12306
rect 36452 12242 36504 12248
rect 36360 11756 36412 11762
rect 36360 11698 36412 11704
rect 36464 11218 36492 12242
rect 36544 12164 36596 12170
rect 36544 12106 36596 12112
rect 36556 11354 36584 12106
rect 36544 11348 36596 11354
rect 36544 11290 36596 11296
rect 36452 11212 36504 11218
rect 36452 11154 36504 11160
rect 36544 10736 36596 10742
rect 36544 10678 36596 10684
rect 36452 10600 36504 10606
rect 36452 10542 36504 10548
rect 36464 10441 36492 10542
rect 36450 10432 36506 10441
rect 36450 10367 36506 10376
rect 36556 10198 36584 10678
rect 36544 10192 36596 10198
rect 36544 10134 36596 10140
rect 36648 9602 36676 12406
rect 36372 9574 36676 9602
rect 35992 9512 36044 9518
rect 35992 9454 36044 9460
rect 36268 9512 36320 9518
rect 36268 9454 36320 9460
rect 35900 8968 35952 8974
rect 35900 8910 35952 8916
rect 35716 8424 35768 8430
rect 35716 8366 35768 8372
rect 35992 5772 36044 5778
rect 35992 5714 36044 5720
rect 35624 4140 35676 4146
rect 35624 4082 35676 4088
rect 35716 4072 35768 4078
rect 35716 4014 35768 4020
rect 35624 3528 35676 3534
rect 35624 3470 35676 3476
rect 35532 3052 35584 3058
rect 35532 2994 35584 3000
rect 35532 2848 35584 2854
rect 35532 2790 35584 2796
rect 35084 1822 35480 1850
rect 35084 800 35112 1822
rect 35544 1714 35572 2790
rect 35452 1686 35572 1714
rect 35256 1488 35308 1494
rect 35256 1430 35308 1436
rect 35268 800 35296 1430
rect 35452 800 35480 1686
rect 35636 800 35664 3470
rect 35728 2854 35756 4014
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 35820 3194 35848 3334
rect 35808 3188 35860 3194
rect 35808 3130 35860 3136
rect 35716 2848 35768 2854
rect 35716 2790 35768 2796
rect 35808 2848 35860 2854
rect 35808 2790 35860 2796
rect 35820 800 35848 2790
rect 36004 2582 36032 5714
rect 36084 4684 36136 4690
rect 36084 4626 36136 4632
rect 35992 2576 36044 2582
rect 35992 2518 36044 2524
rect 36096 800 36124 4626
rect 36372 3942 36400 9574
rect 36544 9512 36596 9518
rect 36596 9460 36676 9466
rect 36544 9454 36676 9460
rect 36556 9438 36676 9454
rect 36648 5846 36676 9438
rect 36636 5840 36688 5846
rect 36636 5782 36688 5788
rect 36544 5568 36596 5574
rect 36544 5510 36596 5516
rect 36452 5024 36504 5030
rect 36452 4966 36504 4972
rect 36464 4622 36492 4966
rect 36556 4758 36584 5510
rect 36832 5166 36860 31726
rect 37016 30870 37044 32166
rect 37004 30864 37056 30870
rect 37004 30806 37056 30812
rect 37016 29238 37044 30806
rect 37004 29232 37056 29238
rect 37004 29174 37056 29180
rect 37004 28620 37056 28626
rect 37004 28562 37056 28568
rect 37016 28529 37044 28562
rect 37002 28520 37058 28529
rect 37002 28455 37058 28464
rect 37004 28416 37056 28422
rect 37004 28358 37056 28364
rect 37016 25974 37044 28358
rect 37108 26586 37136 37742
rect 37200 37330 37228 39200
rect 37372 37868 37424 37874
rect 37372 37810 37424 37816
rect 37384 37466 37412 37810
rect 37372 37460 37424 37466
rect 37372 37402 37424 37408
rect 37188 37324 37240 37330
rect 37188 37266 37240 37272
rect 37476 36394 37504 39578
rect 38106 39200 38162 40000
rect 38934 39200 38990 40000
rect 39854 39200 39910 40000
rect 40682 39200 40738 40000
rect 40776 39432 40828 39438
rect 40776 39374 40828 39380
rect 38120 37466 38148 39200
rect 38476 38888 38528 38894
rect 38476 38830 38528 38836
rect 38108 37460 38160 37466
rect 38108 37402 38160 37408
rect 38108 36576 38160 36582
rect 38108 36518 38160 36524
rect 37384 36366 37504 36394
rect 37278 35456 37334 35465
rect 37278 35391 37334 35400
rect 37292 34542 37320 35391
rect 37280 34536 37332 34542
rect 37280 34478 37332 34484
rect 37188 31816 37240 31822
rect 37188 31758 37240 31764
rect 37200 30802 37228 31758
rect 37188 30796 37240 30802
rect 37188 30738 37240 30744
rect 37188 29504 37240 29510
rect 37188 29446 37240 29452
rect 37200 29238 37228 29446
rect 37188 29232 37240 29238
rect 37188 29174 37240 29180
rect 37384 28762 37412 36366
rect 37464 36236 37516 36242
rect 37464 36178 37516 36184
rect 37476 31754 37504 36178
rect 37832 34060 37884 34066
rect 37832 34002 37884 34008
rect 37740 33924 37792 33930
rect 37740 33866 37792 33872
rect 37464 31748 37516 31754
rect 37464 31690 37516 31696
rect 37648 30252 37700 30258
rect 37648 30194 37700 30200
rect 37372 28756 37424 28762
rect 37372 28698 37424 28704
rect 37554 28656 37610 28665
rect 37280 28620 37332 28626
rect 37332 28580 37412 28608
rect 37554 28591 37556 28600
rect 37280 28562 37332 28568
rect 37188 26920 37240 26926
rect 37188 26862 37240 26868
rect 37280 26920 37332 26926
rect 37280 26862 37332 26868
rect 37200 26586 37228 26862
rect 37096 26580 37148 26586
rect 37096 26522 37148 26528
rect 37188 26580 37240 26586
rect 37188 26522 37240 26528
rect 37004 25968 37056 25974
rect 37004 25910 37056 25916
rect 36912 24880 36964 24886
rect 36912 24822 36964 24828
rect 37096 24880 37148 24886
rect 37096 24822 37148 24828
rect 36924 24750 36952 24822
rect 36912 24744 36964 24750
rect 36912 24686 36964 24692
rect 37004 24676 37056 24682
rect 37004 24618 37056 24624
rect 37016 24585 37044 24618
rect 37002 24576 37058 24585
rect 37002 24511 37058 24520
rect 37108 21622 37136 24822
rect 37096 21616 37148 21622
rect 37096 21558 37148 21564
rect 37004 20800 37056 20806
rect 37004 20742 37056 20748
rect 36912 19304 36964 19310
rect 36912 19246 36964 19252
rect 36924 18222 36952 19246
rect 36912 18216 36964 18222
rect 36912 18158 36964 18164
rect 36912 13796 36964 13802
rect 36912 13738 36964 13744
rect 36924 12434 36952 13738
rect 37016 13190 37044 20742
rect 37292 18222 37320 26862
rect 37384 25498 37412 28580
rect 37608 28591 37610 28600
rect 37556 28562 37608 28568
rect 37660 28370 37688 30194
rect 37752 28694 37780 33866
rect 37740 28688 37792 28694
rect 37740 28630 37792 28636
rect 37740 28552 37792 28558
rect 37738 28520 37740 28529
rect 37792 28520 37794 28529
rect 37738 28455 37794 28464
rect 37660 28342 37780 28370
rect 37648 27328 37700 27334
rect 37648 27270 37700 27276
rect 37660 27130 37688 27270
rect 37648 27124 37700 27130
rect 37648 27066 37700 27072
rect 37464 25968 37516 25974
rect 37464 25910 37516 25916
rect 37372 25492 37424 25498
rect 37372 25434 37424 25440
rect 37384 21622 37412 25434
rect 37372 21616 37424 21622
rect 37372 21558 37424 21564
rect 37280 18216 37332 18222
rect 37280 18158 37332 18164
rect 37280 16040 37332 16046
rect 37280 15982 37332 15988
rect 37004 13184 37056 13190
rect 37004 13126 37056 13132
rect 36924 12406 37044 12434
rect 36912 9648 36964 9654
rect 36912 9590 36964 9596
rect 36924 9178 36952 9590
rect 36912 9172 36964 9178
rect 36912 9114 36964 9120
rect 37016 9110 37044 12406
rect 37292 11218 37320 15982
rect 37280 11212 37332 11218
rect 37280 11154 37332 11160
rect 37186 10432 37242 10441
rect 37186 10367 37242 10376
rect 37004 9104 37056 9110
rect 37004 9046 37056 9052
rect 36912 6792 36964 6798
rect 36912 6734 36964 6740
rect 36636 5160 36688 5166
rect 36636 5102 36688 5108
rect 36820 5160 36872 5166
rect 36820 5102 36872 5108
rect 36648 4842 36676 5102
rect 36820 5024 36872 5030
rect 36820 4966 36872 4972
rect 36648 4814 36768 4842
rect 36544 4752 36596 4758
rect 36544 4694 36596 4700
rect 36636 4684 36688 4690
rect 36636 4626 36688 4632
rect 36452 4616 36504 4622
rect 36452 4558 36504 4564
rect 36360 3936 36412 3942
rect 36360 3878 36412 3884
rect 36544 3936 36596 3942
rect 36544 3878 36596 3884
rect 36556 3670 36584 3878
rect 36544 3664 36596 3670
rect 36544 3606 36596 3612
rect 36176 2916 36228 2922
rect 36176 2858 36228 2864
rect 36268 2916 36320 2922
rect 36268 2858 36320 2864
rect 36188 2582 36216 2858
rect 36176 2576 36228 2582
rect 36176 2518 36228 2524
rect 36280 800 36308 2858
rect 36452 2508 36504 2514
rect 36452 2450 36504 2456
rect 36464 2310 36492 2450
rect 36452 2304 36504 2310
rect 36452 2246 36504 2252
rect 36452 1420 36504 1426
rect 36452 1362 36504 1368
rect 36464 800 36492 1362
rect 36648 800 36676 4626
rect 36740 1222 36768 4814
rect 36832 4486 36860 4966
rect 36820 4480 36872 4486
rect 36820 4422 36872 4428
rect 36820 4072 36872 4078
rect 36820 4014 36872 4020
rect 36728 1216 36780 1222
rect 36728 1158 36780 1164
rect 36832 800 36860 4014
rect 36924 2514 36952 6734
rect 37200 5166 37228 10367
rect 37278 9616 37334 9625
rect 37278 9551 37334 9560
rect 37372 9580 37424 9586
rect 37292 9518 37320 9551
rect 37372 9522 37424 9528
rect 37280 9512 37332 9518
rect 37280 9454 37332 9460
rect 37280 9104 37332 9110
rect 37280 9046 37332 9052
rect 37292 8922 37320 9046
rect 37384 9042 37412 9522
rect 37372 9036 37424 9042
rect 37372 8978 37424 8984
rect 37292 8894 37412 8922
rect 37280 7948 37332 7954
rect 37280 7890 37332 7896
rect 37292 7478 37320 7890
rect 37280 7472 37332 7478
rect 37280 7414 37332 7420
rect 37188 5160 37240 5166
rect 37188 5102 37240 5108
rect 37384 4826 37412 8894
rect 37372 4820 37424 4826
rect 37372 4762 37424 4768
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 36912 2508 36964 2514
rect 36912 2450 36964 2456
rect 37188 2372 37240 2378
rect 37188 2314 37240 2320
rect 37096 2304 37148 2310
rect 37096 2246 37148 2252
rect 37108 800 37136 2246
rect 37200 1494 37228 2314
rect 37188 1488 37240 1494
rect 37188 1430 37240 1436
rect 37292 800 37320 4082
rect 37476 3738 37504 25910
rect 37752 23798 37780 28342
rect 37844 26625 37872 34002
rect 37924 33312 37976 33318
rect 38016 33312 38068 33318
rect 37924 33254 37976 33260
rect 38014 33280 38016 33289
rect 38068 33280 38070 33289
rect 37936 26926 37964 33254
rect 38014 33215 38070 33224
rect 38120 31754 38148 36518
rect 38200 34536 38252 34542
rect 38200 34478 38252 34484
rect 38212 34241 38240 34478
rect 38198 34232 38254 34241
rect 38198 34167 38254 34176
rect 38028 31726 38148 31754
rect 38028 27674 38056 31726
rect 38108 29096 38160 29102
rect 38108 29038 38160 29044
rect 38016 27668 38068 27674
rect 38016 27610 38068 27616
rect 38016 27464 38068 27470
rect 38016 27406 38068 27412
rect 38028 27334 38056 27406
rect 38016 27328 38068 27334
rect 38016 27270 38068 27276
rect 37924 26920 37976 26926
rect 37924 26862 37976 26868
rect 37830 26616 37886 26625
rect 37830 26551 37886 26560
rect 38016 25696 38068 25702
rect 38016 25638 38068 25644
rect 37740 23792 37792 23798
rect 37740 23734 37792 23740
rect 37924 23316 37976 23322
rect 37924 23258 37976 23264
rect 37740 22976 37792 22982
rect 37740 22918 37792 22924
rect 37752 22778 37780 22918
rect 37740 22772 37792 22778
rect 37740 22714 37792 22720
rect 37660 22166 37688 22197
rect 37648 22160 37700 22166
rect 37646 22128 37648 22137
rect 37700 22128 37702 22137
rect 37646 22063 37702 22072
rect 37660 14618 37688 22063
rect 37936 21894 37964 23258
rect 37924 21888 37976 21894
rect 37924 21830 37976 21836
rect 37830 21584 37886 21593
rect 37830 21519 37886 21528
rect 37738 19952 37794 19961
rect 37738 19887 37794 19896
rect 37648 14612 37700 14618
rect 37648 14554 37700 14560
rect 37556 12232 37608 12238
rect 37556 12174 37608 12180
rect 37568 11558 37596 12174
rect 37556 11552 37608 11558
rect 37556 11494 37608 11500
rect 37648 11552 37700 11558
rect 37648 11494 37700 11500
rect 37568 9994 37596 11494
rect 37556 9988 37608 9994
rect 37556 9930 37608 9936
rect 37568 8922 37596 9930
rect 37660 9110 37688 11494
rect 37648 9104 37700 9110
rect 37648 9046 37700 9052
rect 37752 9042 37780 19887
rect 37844 9450 37872 21519
rect 37936 21350 37964 21830
rect 37924 21344 37976 21350
rect 37924 21286 37976 21292
rect 37924 20800 37976 20806
rect 37924 20742 37976 20748
rect 37936 15094 37964 20742
rect 38028 15366 38056 25638
rect 38120 19334 38148 29038
rect 38212 25974 38240 34167
rect 38292 32972 38344 32978
rect 38292 32914 38344 32920
rect 38304 31822 38332 32914
rect 38292 31816 38344 31822
rect 38292 31758 38344 31764
rect 38292 29776 38344 29782
rect 38344 29724 38424 29730
rect 38292 29718 38424 29724
rect 38304 29702 38424 29718
rect 38292 29640 38344 29646
rect 38292 29582 38344 29588
rect 38304 29102 38332 29582
rect 38292 29096 38344 29102
rect 38292 29038 38344 29044
rect 38292 28416 38344 28422
rect 38292 28358 38344 28364
rect 38304 28218 38332 28358
rect 38292 28212 38344 28218
rect 38292 28154 38344 28160
rect 38200 25968 38252 25974
rect 38200 25910 38252 25916
rect 38292 25968 38344 25974
rect 38292 25910 38344 25916
rect 38304 24954 38332 25910
rect 38292 24948 38344 24954
rect 38292 24890 38344 24896
rect 38396 22386 38424 29702
rect 38488 29578 38516 38830
rect 38948 37670 38976 39200
rect 39120 37936 39172 37942
rect 39120 37878 39172 37884
rect 38936 37664 38988 37670
rect 38936 37606 38988 37612
rect 38660 37324 38712 37330
rect 38660 37266 38712 37272
rect 38672 34513 38700 37266
rect 39028 35760 39080 35766
rect 39028 35702 39080 35708
rect 38658 34504 38714 34513
rect 38658 34439 38714 34448
rect 38672 34066 38700 34439
rect 38660 34060 38712 34066
rect 38660 34002 38712 34008
rect 38934 33144 38990 33153
rect 38934 33079 38990 33088
rect 38948 33046 38976 33079
rect 38936 33040 38988 33046
rect 38936 32982 38988 32988
rect 38752 32972 38804 32978
rect 38752 32914 38804 32920
rect 38660 32768 38712 32774
rect 38658 32736 38660 32745
rect 38712 32736 38714 32745
rect 38658 32671 38714 32680
rect 38476 29572 38528 29578
rect 38476 29514 38528 29520
rect 38568 29572 38620 29578
rect 38568 29514 38620 29520
rect 38488 29102 38516 29514
rect 38580 29481 38608 29514
rect 38566 29472 38622 29481
rect 38566 29407 38622 29416
rect 38476 29096 38528 29102
rect 38476 29038 38528 29044
rect 38764 28994 38792 32914
rect 38844 32904 38896 32910
rect 38844 32846 38896 32852
rect 38856 32774 38884 32846
rect 38844 32768 38896 32774
rect 38844 32710 38896 32716
rect 38856 31686 38884 32710
rect 39040 31686 39068 35702
rect 38844 31680 38896 31686
rect 38844 31622 38896 31628
rect 39028 31680 39080 31686
rect 39028 31622 39080 31628
rect 39132 29782 39160 37878
rect 39868 37330 39896 39200
rect 40316 37868 40368 37874
rect 40316 37810 40368 37816
rect 40040 37732 40092 37738
rect 40040 37674 40092 37680
rect 40052 37466 40080 37674
rect 40040 37460 40092 37466
rect 40040 37402 40092 37408
rect 39856 37324 39908 37330
rect 39856 37266 39908 37272
rect 39948 36712 40000 36718
rect 39948 36654 40000 36660
rect 39960 36553 39988 36654
rect 39946 36544 40002 36553
rect 39946 36479 40002 36488
rect 39670 35728 39726 35737
rect 39488 35692 39540 35698
rect 39488 35634 39540 35640
rect 39580 35692 39632 35698
rect 39670 35663 39726 35672
rect 40040 35692 40092 35698
rect 39580 35634 39632 35640
rect 39304 35624 39356 35630
rect 39302 35592 39304 35601
rect 39396 35624 39448 35630
rect 39356 35592 39358 35601
rect 39396 35566 39448 35572
rect 39302 35527 39358 35536
rect 39408 35494 39436 35566
rect 39396 35488 39448 35494
rect 39396 35430 39448 35436
rect 39500 35193 39528 35634
rect 39486 35184 39542 35193
rect 39486 35119 39542 35128
rect 39592 34728 39620 35634
rect 39684 35562 39712 35663
rect 40040 35634 40092 35640
rect 39672 35556 39724 35562
rect 39672 35498 39724 35504
rect 39408 34700 39620 34728
rect 39408 34542 39436 34700
rect 39500 34598 39988 34626
rect 39500 34542 39528 34598
rect 39960 34542 39988 34598
rect 39396 34536 39448 34542
rect 39396 34478 39448 34484
rect 39488 34536 39540 34542
rect 39488 34478 39540 34484
rect 39672 34536 39724 34542
rect 39672 34478 39724 34484
rect 39948 34536 40000 34542
rect 39948 34478 40000 34484
rect 39578 33008 39634 33017
rect 39488 32972 39540 32978
rect 39578 32943 39634 32952
rect 39488 32914 39540 32920
rect 39396 32904 39448 32910
rect 39394 32872 39396 32881
rect 39448 32872 39450 32881
rect 39394 32807 39450 32816
rect 39120 29776 39172 29782
rect 39120 29718 39172 29724
rect 38764 28966 39160 28994
rect 38936 28008 38988 28014
rect 38936 27950 38988 27956
rect 38568 27600 38620 27606
rect 38752 27600 38804 27606
rect 38620 27548 38700 27554
rect 38568 27542 38700 27548
rect 38752 27542 38804 27548
rect 38580 27526 38700 27542
rect 38672 26926 38700 27526
rect 38660 26920 38712 26926
rect 38660 26862 38712 26868
rect 38568 25492 38620 25498
rect 38568 25434 38620 25440
rect 38580 24954 38608 25434
rect 38660 25356 38712 25362
rect 38660 25298 38712 25304
rect 38568 24948 38620 24954
rect 38568 24890 38620 24896
rect 38672 24834 38700 25298
rect 38580 24806 38700 24834
rect 38580 23746 38608 24806
rect 38580 23718 38700 23746
rect 38304 22358 38424 22386
rect 38566 22400 38622 22409
rect 38200 22092 38252 22098
rect 38200 22034 38252 22040
rect 38212 21894 38240 22034
rect 38200 21888 38252 21894
rect 38200 21830 38252 21836
rect 38304 20806 38332 22358
rect 38566 22335 38622 22344
rect 38474 22264 38530 22273
rect 38580 22234 38608 22335
rect 38474 22199 38530 22208
rect 38568 22228 38620 22234
rect 38488 22098 38516 22199
rect 38568 22170 38620 22176
rect 38476 22092 38528 22098
rect 38476 22034 38528 22040
rect 38384 21956 38436 21962
rect 38384 21898 38436 21904
rect 38396 20874 38424 21898
rect 38566 21584 38622 21593
rect 38566 21519 38622 21528
rect 38580 21486 38608 21519
rect 38568 21480 38620 21486
rect 38568 21422 38620 21428
rect 38476 21344 38528 21350
rect 38476 21286 38528 21292
rect 38384 20868 38436 20874
rect 38384 20810 38436 20816
rect 38292 20800 38344 20806
rect 38292 20742 38344 20748
rect 38120 19306 38240 19334
rect 38212 19145 38240 19306
rect 38198 19136 38254 19145
rect 38198 19071 38254 19080
rect 38108 18216 38160 18222
rect 38108 18158 38160 18164
rect 38016 15360 38068 15366
rect 38016 15302 38068 15308
rect 37924 15088 37976 15094
rect 37924 15030 37976 15036
rect 38016 14476 38068 14482
rect 38016 14418 38068 14424
rect 38028 12374 38056 14418
rect 37924 12368 37976 12374
rect 37924 12310 37976 12316
rect 38016 12368 38068 12374
rect 38016 12310 38068 12316
rect 37936 12209 37964 12310
rect 37922 12200 37978 12209
rect 37922 12135 37978 12144
rect 37924 11688 37976 11694
rect 37924 11630 37976 11636
rect 37936 10985 37964 11630
rect 38028 11558 38056 12310
rect 38016 11552 38068 11558
rect 38016 11494 38068 11500
rect 38014 11384 38070 11393
rect 38014 11319 38070 11328
rect 37922 10976 37978 10985
rect 37922 10911 37978 10920
rect 37924 10532 37976 10538
rect 37924 10474 37976 10480
rect 37936 10062 37964 10474
rect 37924 10056 37976 10062
rect 37924 9998 37976 10004
rect 37832 9444 37884 9450
rect 37832 9386 37884 9392
rect 37740 9036 37792 9042
rect 37740 8978 37792 8984
rect 37648 8968 37700 8974
rect 37568 8916 37648 8922
rect 37700 8916 37780 8922
rect 37568 8894 37780 8916
rect 37556 8832 37608 8838
rect 37556 8774 37608 8780
rect 37568 8294 37596 8774
rect 37556 8288 37608 8294
rect 37556 8230 37608 8236
rect 37648 8288 37700 8294
rect 37648 8230 37700 8236
rect 37660 8090 37688 8230
rect 37648 8084 37700 8090
rect 37648 8026 37700 8032
rect 37556 7880 37608 7886
rect 37556 7822 37608 7828
rect 37464 3732 37516 3738
rect 37464 3674 37516 3680
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 37476 800 37504 2926
rect 34520 750 34572 756
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36450 0 36506 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37568 66 37596 7822
rect 37648 5636 37700 5642
rect 37648 5578 37700 5584
rect 37660 4690 37688 5578
rect 37648 4684 37700 4690
rect 37648 4626 37700 4632
rect 37752 4622 37780 8894
rect 38028 7954 38056 11319
rect 38016 7948 38068 7954
rect 38016 7890 38068 7896
rect 38120 7886 38148 18158
rect 38212 16182 38240 19071
rect 38292 18420 38344 18426
rect 38292 18362 38344 18368
rect 38200 16176 38252 16182
rect 38200 16118 38252 16124
rect 38200 12436 38252 12442
rect 38200 12378 38252 12384
rect 38212 11354 38240 12378
rect 38304 11676 38332 18362
rect 38381 11688 38433 11694
rect 38304 11648 38381 11676
rect 38200 11348 38252 11354
rect 38200 11290 38252 11296
rect 38198 10160 38254 10169
rect 38198 10095 38254 10104
rect 38108 7880 38160 7886
rect 38108 7822 38160 7828
rect 38016 5296 38068 5302
rect 38016 5238 38068 5244
rect 37740 4616 37792 4622
rect 37740 4558 37792 4564
rect 37832 3732 37884 3738
rect 37832 3674 37884 3680
rect 37740 3596 37792 3602
rect 37740 3538 37792 3544
rect 37648 2916 37700 2922
rect 37648 2858 37700 2864
rect 37660 800 37688 2858
rect 37556 60 37608 66
rect 37556 2 37608 8
rect 37646 0 37702 800
rect 37752 610 37780 3538
rect 37844 800 37872 3674
rect 38028 3194 38056 5238
rect 38108 3596 38160 3602
rect 38108 3538 38160 3544
rect 38016 3188 38068 3194
rect 38016 3130 38068 3136
rect 38028 2854 38056 3130
rect 38016 2848 38068 2854
rect 38016 2790 38068 2796
rect 37924 2440 37976 2446
rect 37924 2382 37976 2388
rect 37936 1426 37964 2382
rect 37924 1420 37976 1426
rect 37924 1362 37976 1368
rect 38120 800 38148 3538
rect 38212 3194 38240 10095
rect 38304 7342 38332 11648
rect 38381 11630 38433 11636
rect 38488 11506 38516 21286
rect 38672 20244 38700 23718
rect 38764 21486 38792 27542
rect 38844 27464 38896 27470
rect 38844 27406 38896 27412
rect 38752 21480 38804 21486
rect 38752 21422 38804 21428
rect 38752 21344 38804 21350
rect 38752 21286 38804 21292
rect 38764 20806 38792 21286
rect 38752 20800 38804 20806
rect 38752 20742 38804 20748
rect 38856 20398 38884 27406
rect 38948 26994 38976 27950
rect 39028 27532 39080 27538
rect 39028 27474 39080 27480
rect 38936 26988 38988 26994
rect 38936 26930 38988 26936
rect 38934 26752 38990 26761
rect 38934 26687 38990 26696
rect 38844 20392 38896 20398
rect 38844 20334 38896 20340
rect 38672 20216 38884 20244
rect 38566 20088 38622 20097
rect 38566 20023 38568 20032
rect 38620 20023 38622 20032
rect 38568 19994 38620 20000
rect 38752 19916 38804 19922
rect 38752 19858 38804 19864
rect 38658 19816 38714 19825
rect 38658 19751 38660 19760
rect 38712 19751 38714 19760
rect 38660 19722 38712 19728
rect 38764 19689 38792 19858
rect 38750 19680 38806 19689
rect 38750 19615 38806 19624
rect 38568 18216 38620 18222
rect 38568 18158 38620 18164
rect 38580 17921 38608 18158
rect 38566 17912 38622 17921
rect 38566 17847 38622 17856
rect 38660 15564 38712 15570
rect 38660 15506 38712 15512
rect 38568 12436 38620 12442
rect 38568 12378 38620 12384
rect 38580 11694 38608 12378
rect 38672 12345 38700 15506
rect 38658 12336 38714 12345
rect 38658 12271 38714 12280
rect 38856 11937 38884 20216
rect 38842 11928 38898 11937
rect 38672 11898 38792 11914
rect 38660 11892 38792 11898
rect 38712 11886 38792 11892
rect 38660 11834 38712 11840
rect 38764 11812 38792 11886
rect 38842 11863 38898 11872
rect 38844 11824 38896 11830
rect 38764 11784 38844 11812
rect 38844 11766 38896 11772
rect 38568 11688 38620 11694
rect 38568 11630 38620 11636
rect 38660 11688 38712 11694
rect 38712 11648 38792 11676
rect 38660 11630 38712 11636
rect 38764 11558 38792 11648
rect 38752 11552 38804 11558
rect 38396 11478 38516 11506
rect 38566 11520 38622 11529
rect 38396 11354 38424 11478
rect 38622 11500 38752 11506
rect 38948 11540 38976 26687
rect 39040 25294 39068 27474
rect 39028 25288 39080 25294
rect 39028 25230 39080 25236
rect 39028 20392 39080 20398
rect 39028 20334 39080 20340
rect 39040 19786 39068 20334
rect 39132 19825 39160 28966
rect 39304 28144 39356 28150
rect 39304 28086 39356 28092
rect 39396 28144 39448 28150
rect 39396 28086 39448 28092
rect 39316 27713 39344 28086
rect 39302 27704 39358 27713
rect 39302 27639 39358 27648
rect 39304 27464 39356 27470
rect 39304 27406 39356 27412
rect 39212 25832 39264 25838
rect 39212 25774 39264 25780
rect 39224 23254 39252 25774
rect 39316 24750 39344 27406
rect 39408 26926 39436 28086
rect 39396 26920 39448 26926
rect 39396 26862 39448 26868
rect 39396 25832 39448 25838
rect 39396 25774 39448 25780
rect 39408 25498 39436 25774
rect 39396 25492 39448 25498
rect 39396 25434 39448 25440
rect 39500 24954 39528 32914
rect 39592 32842 39620 32943
rect 39580 32836 39632 32842
rect 39580 32778 39632 32784
rect 39684 28694 39712 34478
rect 39948 34060 40000 34066
rect 39948 34002 40000 34008
rect 39960 33697 39988 34002
rect 39946 33688 40002 33697
rect 39946 33623 40002 33632
rect 40052 33454 40080 35634
rect 40132 33584 40184 33590
rect 40132 33526 40184 33532
rect 40040 33448 40092 33454
rect 40144 33425 40172 33526
rect 40040 33390 40092 33396
rect 40130 33416 40186 33425
rect 39948 32768 40000 32774
rect 39948 32710 40000 32716
rect 39960 32502 39988 32710
rect 39948 32496 40000 32502
rect 39948 32438 40000 32444
rect 40052 32366 40080 33390
rect 40130 33351 40186 33360
rect 39948 32360 40000 32366
rect 39946 32328 39948 32337
rect 40040 32360 40092 32366
rect 40000 32328 40002 32337
rect 40040 32302 40092 32308
rect 39946 32263 40002 32272
rect 40052 30122 40080 32302
rect 40040 30116 40092 30122
rect 40040 30058 40092 30064
rect 40132 29640 40184 29646
rect 39960 29588 40132 29594
rect 39960 29582 40184 29588
rect 39960 29566 40172 29582
rect 39960 29510 39988 29566
rect 39948 29504 40000 29510
rect 39948 29446 40000 29452
rect 39672 28688 39724 28694
rect 39672 28630 39724 28636
rect 40038 27840 40094 27849
rect 40038 27775 40094 27784
rect 40052 27674 40080 27775
rect 40040 27668 40092 27674
rect 40040 27610 40092 27616
rect 39578 27568 39634 27577
rect 39578 27503 39580 27512
rect 39632 27503 39634 27512
rect 39580 27474 39632 27480
rect 39672 27464 39724 27470
rect 39672 27406 39724 27412
rect 39684 26994 39712 27406
rect 39672 26988 39724 26994
rect 39672 26930 39724 26936
rect 39854 25936 39910 25945
rect 39854 25871 39910 25880
rect 39868 25838 39896 25871
rect 39580 25832 39632 25838
rect 39580 25774 39632 25780
rect 39856 25832 39908 25838
rect 39856 25774 39908 25780
rect 39592 25702 39620 25774
rect 39580 25696 39632 25702
rect 39580 25638 39632 25644
rect 39868 25226 39896 25774
rect 39856 25220 39908 25226
rect 39856 25162 39908 25168
rect 39488 24948 39540 24954
rect 39488 24890 39540 24896
rect 39304 24744 39356 24750
rect 39304 24686 39356 24692
rect 39212 23248 39264 23254
rect 39212 23190 39264 23196
rect 39396 21480 39448 21486
rect 39396 21422 39448 21428
rect 39118 19816 39174 19825
rect 39028 19780 39080 19786
rect 39118 19751 39174 19760
rect 39028 19722 39080 19728
rect 39040 18970 39068 19722
rect 39028 18964 39080 18970
rect 39028 18906 39080 18912
rect 39304 18216 39356 18222
rect 39132 18164 39304 18170
rect 39132 18158 39356 18164
rect 39132 18142 39344 18158
rect 39028 13456 39080 13462
rect 39028 13398 39080 13404
rect 39040 11762 39068 13398
rect 39132 12850 39160 18142
rect 39212 18080 39264 18086
rect 39316 18057 39344 18142
rect 39212 18022 39264 18028
rect 39302 18048 39358 18057
rect 39120 12844 39172 12850
rect 39120 12786 39172 12792
rect 39120 12640 39172 12646
rect 39120 12582 39172 12588
rect 39028 11756 39080 11762
rect 39028 11698 39080 11704
rect 38622 11494 38804 11500
rect 38856 11512 38976 11540
rect 38622 11478 38792 11494
rect 38566 11455 38622 11464
rect 38474 11384 38530 11393
rect 38384 11348 38436 11354
rect 38658 11384 38714 11393
rect 38530 11354 38608 11370
rect 38530 11348 38620 11354
rect 38530 11342 38568 11348
rect 38474 11319 38530 11328
rect 38384 11290 38436 11296
rect 38658 11319 38714 11328
rect 38568 11290 38620 11296
rect 38568 11212 38620 11218
rect 38568 11154 38620 11160
rect 38580 7886 38608 11154
rect 38672 8362 38700 11319
rect 38856 11286 38884 11512
rect 38934 11384 38990 11393
rect 38934 11319 38990 11328
rect 38844 11280 38896 11286
rect 38844 11222 38896 11228
rect 38750 11112 38806 11121
rect 38750 11047 38806 11056
rect 38764 8430 38792 11047
rect 38752 8424 38804 8430
rect 38752 8366 38804 8372
rect 38660 8356 38712 8362
rect 38660 8298 38712 8304
rect 38842 8120 38898 8129
rect 38842 8055 38898 8064
rect 38856 8022 38884 8055
rect 38844 8016 38896 8022
rect 38844 7958 38896 7964
rect 38568 7880 38620 7886
rect 38568 7822 38620 7828
rect 38660 7880 38712 7886
rect 38660 7822 38712 7828
rect 38292 7336 38344 7342
rect 38292 7278 38344 7284
rect 38476 7336 38528 7342
rect 38476 7278 38528 7284
rect 38488 7154 38516 7278
rect 38672 7274 38700 7822
rect 38660 7268 38712 7274
rect 38660 7210 38712 7216
rect 38752 7268 38804 7274
rect 38752 7210 38804 7216
rect 38764 7154 38792 7210
rect 38488 7126 38792 7154
rect 38752 5160 38804 5166
rect 38752 5102 38804 5108
rect 38660 4072 38712 4078
rect 38660 4014 38712 4020
rect 38568 4004 38620 4010
rect 38568 3946 38620 3952
rect 38200 3188 38252 3194
rect 38200 3130 38252 3136
rect 38580 2666 38608 3946
rect 38292 2644 38344 2650
rect 38292 2586 38344 2592
rect 38488 2638 38608 2666
rect 38304 800 38332 2586
rect 38488 800 38516 2638
rect 38568 2032 38620 2038
rect 38568 1974 38620 1980
rect 38580 1290 38608 1974
rect 38568 1284 38620 1290
rect 38568 1226 38620 1232
rect 38672 800 38700 4014
rect 38764 2582 38792 5102
rect 38948 3398 38976 11319
rect 39028 8424 39080 8430
rect 39028 8366 39080 8372
rect 39040 7410 39068 8366
rect 39028 7404 39080 7410
rect 39028 7346 39080 7352
rect 38936 3392 38988 3398
rect 38936 3334 38988 3340
rect 39132 2582 39160 12582
rect 39224 10198 39252 18022
rect 39302 17983 39358 17992
rect 39304 16244 39356 16250
rect 39304 16186 39356 16192
rect 39212 10192 39264 10198
rect 39212 10134 39264 10140
rect 39212 7948 39264 7954
rect 39212 7890 39264 7896
rect 39224 7002 39252 7890
rect 39316 7410 39344 16186
rect 39408 13394 39436 21422
rect 39396 13388 39448 13394
rect 39396 13330 39448 13336
rect 39394 12200 39450 12209
rect 39394 12135 39450 12144
rect 39408 11830 39436 12135
rect 39396 11824 39448 11830
rect 39396 11766 39448 11772
rect 39500 11506 39528 24890
rect 40040 22092 40092 22098
rect 40040 22034 40092 22040
rect 40052 21622 40080 22034
rect 40040 21616 40092 21622
rect 40040 21558 40092 21564
rect 39854 19000 39910 19009
rect 39854 18935 39910 18944
rect 40038 19000 40094 19009
rect 40038 18935 40094 18944
rect 39762 18592 39818 18601
rect 39762 18527 39818 18536
rect 39776 18290 39804 18527
rect 39868 18426 39896 18935
rect 40052 18766 40080 18935
rect 40040 18760 40092 18766
rect 40040 18702 40092 18708
rect 39856 18420 39908 18426
rect 39856 18362 39908 18368
rect 39764 18284 39816 18290
rect 39592 18244 39764 18272
rect 39592 12782 39620 18244
rect 39764 18226 39816 18232
rect 40132 17808 40184 17814
rect 40132 17750 40184 17756
rect 40040 16720 40092 16726
rect 40038 16688 40040 16697
rect 40092 16688 40094 16697
rect 40038 16623 40094 16632
rect 39764 13388 39816 13394
rect 39764 13330 39816 13336
rect 39672 12844 39724 12850
rect 39672 12786 39724 12792
rect 39580 12776 39632 12782
rect 39580 12718 39632 12724
rect 39580 12096 39632 12102
rect 39580 12038 39632 12044
rect 39592 11626 39620 12038
rect 39580 11620 39632 11626
rect 39580 11562 39632 11568
rect 39408 11478 39528 11506
rect 39408 11393 39436 11478
rect 39394 11384 39450 11393
rect 39394 11319 39450 11328
rect 39578 10976 39634 10985
rect 39578 10911 39634 10920
rect 39396 8628 39448 8634
rect 39396 8570 39448 8576
rect 39408 8430 39436 8570
rect 39396 8424 39448 8430
rect 39396 8366 39448 8372
rect 39592 8294 39620 10911
rect 39684 10538 39712 12786
rect 39776 12782 39804 13330
rect 39764 12776 39816 12782
rect 39764 12718 39816 12724
rect 40144 12434 40172 17750
rect 40224 16788 40276 16794
rect 40224 16730 40276 16736
rect 40236 16250 40264 16730
rect 40224 16244 40276 16250
rect 40224 16186 40276 16192
rect 40328 15638 40356 37810
rect 40696 37466 40724 39200
rect 40684 37460 40736 37466
rect 40684 37402 40736 37408
rect 40500 34536 40552 34542
rect 40500 34478 40552 34484
rect 40512 34202 40540 34478
rect 40500 34196 40552 34202
rect 40500 34138 40552 34144
rect 40408 34060 40460 34066
rect 40408 34002 40460 34008
rect 40420 32366 40448 34002
rect 40500 32904 40552 32910
rect 40500 32846 40552 32852
rect 40408 32360 40460 32366
rect 40408 32302 40460 32308
rect 40512 31754 40540 32846
rect 40682 32736 40738 32745
rect 40682 32671 40738 32680
rect 40696 32366 40724 32671
rect 40684 32360 40736 32366
rect 40684 32302 40736 32308
rect 40500 31748 40552 31754
rect 40500 31690 40552 31696
rect 40684 30116 40736 30122
rect 40684 30058 40736 30064
rect 40590 28112 40646 28121
rect 40590 28047 40646 28056
rect 40500 27396 40552 27402
rect 40500 27338 40552 27344
rect 40512 27305 40540 27338
rect 40498 27296 40554 27305
rect 40498 27231 40554 27240
rect 40408 26988 40460 26994
rect 40408 26930 40460 26936
rect 40420 21350 40448 26930
rect 40500 26512 40552 26518
rect 40498 26480 40500 26489
rect 40552 26480 40554 26489
rect 40498 26415 40554 26424
rect 40498 25528 40554 25537
rect 40498 25463 40554 25472
rect 40512 25362 40540 25463
rect 40500 25356 40552 25362
rect 40500 25298 40552 25304
rect 40500 24744 40552 24750
rect 40498 24712 40500 24721
rect 40552 24712 40554 24721
rect 40498 24647 40554 24656
rect 40500 22092 40552 22098
rect 40500 22034 40552 22040
rect 40408 21344 40460 21350
rect 40408 21286 40460 21292
rect 40408 17332 40460 17338
rect 40408 17274 40460 17280
rect 40420 16658 40448 17274
rect 40408 16652 40460 16658
rect 40408 16594 40460 16600
rect 40224 15632 40276 15638
rect 40316 15632 40368 15638
rect 40224 15574 40276 15580
rect 40314 15600 40316 15609
rect 40368 15600 40370 15609
rect 39960 12406 40172 12434
rect 39764 11756 39816 11762
rect 39764 11698 39816 11704
rect 39672 10532 39724 10538
rect 39672 10474 39724 10480
rect 39684 9926 39712 10474
rect 39672 9920 39724 9926
rect 39672 9862 39724 9868
rect 39776 9110 39804 11698
rect 39856 9920 39908 9926
rect 39856 9862 39908 9868
rect 39764 9104 39816 9110
rect 39764 9046 39816 9052
rect 39592 8266 39804 8294
rect 39486 8120 39542 8129
rect 39486 8055 39542 8064
rect 39500 7954 39528 8055
rect 39488 7948 39540 7954
rect 39488 7890 39540 7896
rect 39304 7404 39356 7410
rect 39304 7346 39356 7352
rect 39212 6996 39264 7002
rect 39212 6938 39264 6944
rect 39212 5160 39264 5166
rect 39212 5102 39264 5108
rect 39224 4010 39252 5102
rect 39488 4684 39540 4690
rect 39488 4626 39540 4632
rect 39396 4140 39448 4146
rect 39396 4082 39448 4088
rect 39212 4004 39264 4010
rect 39212 3946 39264 3952
rect 39408 3754 39436 4082
rect 39224 3726 39436 3754
rect 39500 3738 39528 4626
rect 39672 4004 39724 4010
rect 39672 3946 39724 3952
rect 39488 3732 39540 3738
rect 38752 2576 38804 2582
rect 38752 2518 38804 2524
rect 39120 2576 39172 2582
rect 39120 2518 39172 2524
rect 39028 2372 39080 2378
rect 39028 2314 39080 2320
rect 39040 1170 39068 2314
rect 39224 2122 39252 3726
rect 39488 3674 39540 3680
rect 39304 3596 39356 3602
rect 39304 3538 39356 3544
rect 38856 1142 39068 1170
rect 39132 2094 39252 2122
rect 38856 800 38884 1142
rect 39132 800 39160 2094
rect 39316 800 39344 3538
rect 39488 3188 39540 3194
rect 39488 3130 39540 3136
rect 39580 3188 39632 3194
rect 39580 3130 39632 3136
rect 39500 2990 39528 3130
rect 39488 2984 39540 2990
rect 39488 2926 39540 2932
rect 39592 2666 39620 3130
rect 39408 2638 39620 2666
rect 39408 2514 39436 2638
rect 39396 2508 39448 2514
rect 39396 2450 39448 2456
rect 39488 2508 39540 2514
rect 39488 2450 39540 2456
rect 39500 800 39528 2450
rect 39684 800 39712 3946
rect 37740 604 37792 610
rect 37740 546 37792 552
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38384 468 38436 474
rect 38384 410 38436 416
rect 38396 66 38424 410
rect 38384 60 38436 66
rect 38384 2 38436 8
rect 38474 0 38530 800
rect 38568 604 38620 610
rect 38568 546 38620 552
rect 38580 377 38608 546
rect 38566 368 38622 377
rect 38566 303 38622 312
rect 38658 0 38714 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39776 66 39804 8266
rect 39868 7698 39896 9862
rect 39960 8634 39988 12406
rect 39948 8628 40000 8634
rect 39948 8570 40000 8576
rect 40236 8090 40264 15574
rect 40314 15535 40370 15544
rect 40408 15496 40460 15502
rect 40408 15438 40460 15444
rect 40420 14385 40448 15438
rect 40406 14376 40462 14385
rect 40406 14311 40462 14320
rect 40408 14068 40460 14074
rect 40408 14010 40460 14016
rect 40420 13938 40448 14010
rect 40408 13932 40460 13938
rect 40408 13874 40460 13880
rect 40406 13832 40462 13841
rect 40406 13767 40408 13776
rect 40460 13767 40462 13776
rect 40408 13738 40460 13744
rect 40408 12980 40460 12986
rect 40408 12922 40460 12928
rect 40316 12708 40368 12714
rect 40316 12650 40368 12656
rect 40328 9042 40356 12650
rect 40316 9036 40368 9042
rect 40316 8978 40368 8984
rect 40420 8566 40448 12922
rect 40512 12102 40540 22034
rect 40500 12096 40552 12102
rect 40500 12038 40552 12044
rect 40512 9450 40540 12038
rect 40500 9444 40552 9450
rect 40500 9386 40552 9392
rect 40408 8560 40460 8566
rect 40408 8502 40460 8508
rect 40224 8084 40276 8090
rect 40224 8026 40276 8032
rect 40040 8016 40092 8022
rect 40040 7958 40092 7964
rect 39868 7670 39988 7698
rect 39856 7404 39908 7410
rect 39856 7346 39908 7352
rect 39868 2582 39896 7346
rect 39960 4758 39988 7670
rect 40052 7410 40080 7958
rect 40040 7404 40092 7410
rect 40040 7346 40092 7352
rect 39948 4752 40000 4758
rect 39948 4694 40000 4700
rect 40316 4684 40368 4690
rect 40316 4626 40368 4632
rect 39948 4072 40000 4078
rect 39948 4014 40000 4020
rect 39856 2576 39908 2582
rect 39856 2518 39908 2524
rect 39960 800 39988 4014
rect 40132 2848 40184 2854
rect 40132 2790 40184 2796
rect 40144 800 40172 2790
rect 40328 800 40356 4626
rect 40500 3596 40552 3602
rect 40500 3538 40552 3544
rect 40512 800 40540 3538
rect 40604 2582 40632 28047
rect 40696 25226 40724 30058
rect 40684 25220 40736 25226
rect 40684 25162 40736 25168
rect 40696 24750 40724 25162
rect 40684 24744 40736 24750
rect 40684 24686 40736 24692
rect 40788 22094 40816 39374
rect 41602 39200 41658 40000
rect 41972 39228 42024 39234
rect 41616 37398 41644 39200
rect 42430 39200 42486 40000
rect 43350 39200 43406 40000
rect 44178 39200 44234 40000
rect 44732 39364 44784 39370
rect 44732 39306 44784 39312
rect 41972 39170 42024 39176
rect 41696 37800 41748 37806
rect 41696 37742 41748 37748
rect 41328 37392 41380 37398
rect 41328 37334 41380 37340
rect 41604 37392 41656 37398
rect 41604 37334 41656 37340
rect 41052 37256 41104 37262
rect 40880 37204 41052 37210
rect 40880 37198 41104 37204
rect 40880 37182 41092 37198
rect 40880 37126 40908 37182
rect 40868 37120 40920 37126
rect 40868 37062 40920 37068
rect 41144 35624 41196 35630
rect 41144 35566 41196 35572
rect 41052 35556 41104 35562
rect 41052 35498 41104 35504
rect 40960 35488 41012 35494
rect 40960 35430 41012 35436
rect 40868 34672 40920 34678
rect 40868 34614 40920 34620
rect 40880 33833 40908 34614
rect 40972 34202 41000 35430
rect 40960 34196 41012 34202
rect 40960 34138 41012 34144
rect 40866 33824 40922 33833
rect 40866 33759 40922 33768
rect 40868 31816 40920 31822
rect 40868 31758 40920 31764
rect 40880 26994 40908 31758
rect 40972 31482 41000 34138
rect 40960 31476 41012 31482
rect 40960 31418 41012 31424
rect 40960 27328 41012 27334
rect 40960 27270 41012 27276
rect 40972 26994 41000 27270
rect 40868 26988 40920 26994
rect 40868 26930 40920 26936
rect 40960 26988 41012 26994
rect 40960 26930 41012 26936
rect 41064 26874 41092 35498
rect 41156 34082 41184 35566
rect 41340 35494 41368 37334
rect 41708 37330 41736 37742
rect 41696 37324 41748 37330
rect 41696 37266 41748 37272
rect 41510 36544 41566 36553
rect 41510 36479 41566 36488
rect 41418 36272 41474 36281
rect 41418 36207 41474 36216
rect 41432 36174 41460 36207
rect 41524 36174 41552 36479
rect 41420 36168 41472 36174
rect 41420 36110 41472 36116
rect 41512 36168 41564 36174
rect 41512 36110 41564 36116
rect 41418 35592 41474 35601
rect 41418 35527 41474 35536
rect 41328 35488 41380 35494
rect 41328 35430 41380 35436
rect 41326 35320 41382 35329
rect 41326 35255 41382 35264
rect 41340 35154 41368 35255
rect 41432 35154 41460 35527
rect 41328 35148 41380 35154
rect 41328 35090 41380 35096
rect 41420 35148 41472 35154
rect 41420 35090 41472 35096
rect 41326 35048 41382 35057
rect 41326 34983 41382 34992
rect 41340 34406 41368 34983
rect 41512 34672 41564 34678
rect 41512 34614 41564 34620
rect 41524 34542 41552 34614
rect 41512 34536 41564 34542
rect 41512 34478 41564 34484
rect 41328 34400 41380 34406
rect 41696 34400 41748 34406
rect 41328 34342 41380 34348
rect 41432 34348 41696 34354
rect 41432 34342 41748 34348
rect 41432 34326 41736 34342
rect 41432 34202 41460 34326
rect 41510 34232 41566 34241
rect 41420 34196 41472 34202
rect 41510 34167 41512 34176
rect 41420 34138 41472 34144
rect 41564 34167 41566 34176
rect 41512 34138 41564 34144
rect 41156 34054 41276 34082
rect 41144 33924 41196 33930
rect 41144 33866 41196 33872
rect 41156 33658 41184 33866
rect 41144 33652 41196 33658
rect 41144 33594 41196 33600
rect 41248 33153 41276 34054
rect 41326 33688 41382 33697
rect 41326 33623 41382 33632
rect 41340 33522 41368 33623
rect 41328 33516 41380 33522
rect 41328 33458 41380 33464
rect 41696 33380 41748 33386
rect 41432 33340 41696 33368
rect 41234 33144 41290 33153
rect 41234 33079 41290 33088
rect 41432 31958 41460 33340
rect 41696 33322 41748 33328
rect 41984 32609 42012 39170
rect 42248 38004 42300 38010
rect 42248 37946 42300 37952
rect 42260 37074 42288 37946
rect 42340 37800 42392 37806
rect 42340 37742 42392 37748
rect 42352 37330 42380 37742
rect 42340 37324 42392 37330
rect 42340 37266 42392 37272
rect 42260 37046 42380 37074
rect 42154 36952 42210 36961
rect 42064 36916 42116 36922
rect 42154 36887 42210 36896
rect 42248 36916 42300 36922
rect 42064 36858 42116 36864
rect 42076 36156 42104 36858
rect 42168 36310 42196 36887
rect 42248 36858 42300 36864
rect 42260 36650 42288 36858
rect 42248 36644 42300 36650
rect 42248 36586 42300 36592
rect 42156 36304 42208 36310
rect 42156 36246 42208 36252
rect 42248 36304 42300 36310
rect 42248 36246 42300 36252
rect 42260 36156 42288 36246
rect 42076 36128 42288 36156
rect 42352 34082 42380 37046
rect 42444 36718 42472 39200
rect 42524 37664 42576 37670
rect 42524 37606 42576 37612
rect 43076 37664 43128 37670
rect 43076 37606 43128 37612
rect 42536 37466 42564 37606
rect 42524 37460 42576 37466
rect 42524 37402 42576 37408
rect 42892 37324 42944 37330
rect 42892 37266 42944 37272
rect 42432 36712 42484 36718
rect 42432 36654 42484 36660
rect 42352 34066 42472 34082
rect 42248 34060 42300 34066
rect 42076 34020 42248 34048
rect 42076 32978 42104 34020
rect 42352 34060 42484 34066
rect 42352 34054 42432 34060
rect 42248 34002 42300 34008
rect 42432 34002 42484 34008
rect 42616 34060 42668 34066
rect 42616 34002 42668 34008
rect 42444 33946 42472 34002
rect 42444 33918 42564 33946
rect 42154 33144 42210 33153
rect 42154 33079 42210 33088
rect 42168 33046 42196 33079
rect 42156 33040 42208 33046
rect 42432 33040 42484 33046
rect 42156 32982 42208 32988
rect 42260 33000 42432 33028
rect 42064 32972 42116 32978
rect 42064 32914 42116 32920
rect 41970 32600 42026 32609
rect 41970 32535 42026 32544
rect 41972 32428 42024 32434
rect 41972 32370 42024 32376
rect 41788 32292 41840 32298
rect 41788 32234 41840 32240
rect 41420 31952 41472 31958
rect 41420 31894 41472 31900
rect 41328 31884 41380 31890
rect 41328 31826 41380 31832
rect 41340 31754 41368 31826
rect 41800 31754 41828 32234
rect 41984 32230 42012 32370
rect 42076 32230 42104 32914
rect 41972 32224 42024 32230
rect 41972 32166 42024 32172
rect 42064 32224 42116 32230
rect 42064 32166 42116 32172
rect 41328 31748 41380 31754
rect 41328 31690 41380 31696
rect 41788 31748 41840 31754
rect 41788 31690 41840 31696
rect 41144 31680 41196 31686
rect 41144 31622 41196 31628
rect 40696 22066 40816 22094
rect 40880 26846 41092 26874
rect 40696 5642 40724 22066
rect 40776 17672 40828 17678
rect 40776 17614 40828 17620
rect 40788 14482 40816 17614
rect 40776 14476 40828 14482
rect 40776 14418 40828 14424
rect 40880 14074 40908 26846
rect 40960 26580 41012 26586
rect 40960 26522 41012 26528
rect 40972 26217 41000 26522
rect 41052 26444 41104 26450
rect 41052 26386 41104 26392
rect 41064 26353 41092 26386
rect 41050 26344 41106 26353
rect 41050 26279 41106 26288
rect 40958 26208 41014 26217
rect 40958 26143 41014 26152
rect 40960 24132 41012 24138
rect 40960 24074 41012 24080
rect 41052 24132 41104 24138
rect 41052 24074 41104 24080
rect 40972 24041 41000 24074
rect 40958 24032 41014 24041
rect 40958 23967 41014 23976
rect 40958 18728 41014 18737
rect 40958 18663 40960 18672
rect 41012 18663 41014 18672
rect 40960 18634 41012 18640
rect 40960 17672 41012 17678
rect 40960 17614 41012 17620
rect 40972 17270 41000 17614
rect 40960 17264 41012 17270
rect 40960 17206 41012 17212
rect 40960 16720 41012 16726
rect 40960 16662 41012 16668
rect 40868 14068 40920 14074
rect 40868 14010 40920 14016
rect 40972 7410 41000 16662
rect 41064 16658 41092 24074
rect 41156 16726 41184 31622
rect 41604 29504 41656 29510
rect 41604 29446 41656 29452
rect 41510 28248 41566 28257
rect 41510 28183 41566 28192
rect 41524 28014 41552 28183
rect 41512 28008 41564 28014
rect 41512 27950 41564 27956
rect 41236 27668 41288 27674
rect 41236 27610 41288 27616
rect 41420 27668 41472 27674
rect 41420 27610 41472 27616
rect 41248 22094 41276 27610
rect 41328 27328 41380 27334
rect 41328 27270 41380 27276
rect 41340 25362 41368 27270
rect 41432 27062 41460 27610
rect 41510 27568 41566 27577
rect 41510 27503 41512 27512
rect 41564 27503 41566 27512
rect 41512 27474 41564 27480
rect 41420 27056 41472 27062
rect 41420 26998 41472 27004
rect 41616 26926 41644 29446
rect 42064 29232 42116 29238
rect 42064 29174 42116 29180
rect 42076 28529 42104 29174
rect 42062 28520 42118 28529
rect 42062 28455 42118 28464
rect 42064 27532 42116 27538
rect 42064 27474 42116 27480
rect 41696 27464 41748 27470
rect 41696 27406 41748 27412
rect 41604 26920 41656 26926
rect 41604 26862 41656 26868
rect 41510 26752 41566 26761
rect 41510 26687 41566 26696
rect 41524 26586 41552 26687
rect 41512 26580 41564 26586
rect 41512 26522 41564 26528
rect 41420 26036 41472 26042
rect 41420 25978 41472 25984
rect 41512 26036 41564 26042
rect 41512 25978 41564 25984
rect 41328 25356 41380 25362
rect 41328 25298 41380 25304
rect 41432 25265 41460 25978
rect 41524 25537 41552 25978
rect 41510 25528 41566 25537
rect 41510 25463 41566 25472
rect 41512 25356 41564 25362
rect 41512 25298 41564 25304
rect 41418 25256 41474 25265
rect 41418 25191 41474 25200
rect 41420 24744 41472 24750
rect 41420 24686 41472 24692
rect 41248 22066 41368 22094
rect 41340 18834 41368 22066
rect 41432 21486 41460 24686
rect 41524 21894 41552 25298
rect 41512 21888 41564 21894
rect 41512 21830 41564 21836
rect 41420 21480 41472 21486
rect 41420 21422 41472 21428
rect 41510 21448 41566 21457
rect 41510 21383 41512 21392
rect 41564 21383 41566 21392
rect 41512 21354 41564 21360
rect 41328 18828 41380 18834
rect 41328 18770 41380 18776
rect 41418 18456 41474 18465
rect 41418 18391 41474 18400
rect 41432 18358 41460 18391
rect 41420 18352 41472 18358
rect 41420 18294 41472 18300
rect 41236 18080 41288 18086
rect 41236 18022 41288 18028
rect 41420 18080 41472 18086
rect 41420 18022 41472 18028
rect 41144 16720 41196 16726
rect 41144 16662 41196 16668
rect 41052 16652 41104 16658
rect 41052 16594 41104 16600
rect 41144 16244 41196 16250
rect 41144 16186 41196 16192
rect 41050 15736 41106 15745
rect 41050 15671 41052 15680
rect 41104 15671 41106 15680
rect 41052 15642 41104 15648
rect 41156 15094 41184 16186
rect 41052 15088 41104 15094
rect 41052 15030 41104 15036
rect 41144 15088 41196 15094
rect 41144 15030 41196 15036
rect 41064 14634 41092 15030
rect 41064 14618 41184 14634
rect 41064 14612 41196 14618
rect 41064 14606 41144 14612
rect 41144 14554 41196 14560
rect 41144 14000 41196 14006
rect 41142 13968 41144 13977
rect 41196 13968 41198 13977
rect 41142 13903 41198 13912
rect 41248 10826 41276 18022
rect 41432 17921 41460 18022
rect 41418 17912 41474 17921
rect 41418 17847 41474 17856
rect 41328 17264 41380 17270
rect 41328 17206 41380 17212
rect 41340 15706 41368 17206
rect 41328 15700 41380 15706
rect 41328 15642 41380 15648
rect 41510 15600 41566 15609
rect 41510 15535 41512 15544
rect 41564 15535 41566 15544
rect 41512 15506 41564 15512
rect 41616 11370 41644 26862
rect 41708 12209 41736 27406
rect 41788 27396 41840 27402
rect 41788 27338 41840 27344
rect 41800 24449 41828 27338
rect 41880 26920 41932 26926
rect 41880 26862 41932 26868
rect 41892 25362 41920 26862
rect 41880 25356 41932 25362
rect 41880 25298 41932 25304
rect 41786 24440 41842 24449
rect 41786 24375 41842 24384
rect 41788 18284 41840 18290
rect 41788 18226 41840 18232
rect 41800 18057 41828 18226
rect 41786 18048 41842 18057
rect 41786 17983 41842 17992
rect 41786 15736 41842 15745
rect 41786 15671 41788 15680
rect 41840 15671 41842 15680
rect 41788 15642 41840 15648
rect 41800 15366 41828 15642
rect 41788 15360 41840 15366
rect 41788 15302 41840 15308
rect 42076 12306 42104 27474
rect 42260 24274 42288 33000
rect 42432 32982 42484 32988
rect 42340 32836 42392 32842
rect 42340 32778 42392 32784
rect 42352 26353 42380 32778
rect 42536 28558 42564 33918
rect 42628 29510 42656 34002
rect 42708 33380 42760 33386
rect 42708 33322 42760 33328
rect 42720 32774 42748 33322
rect 42800 32904 42852 32910
rect 42800 32846 42852 32852
rect 42708 32768 42760 32774
rect 42708 32710 42760 32716
rect 42706 32600 42762 32609
rect 42706 32535 42762 32544
rect 42616 29504 42668 29510
rect 42616 29446 42668 29452
rect 42432 28552 42484 28558
rect 42432 28494 42484 28500
rect 42524 28552 42576 28558
rect 42524 28494 42576 28500
rect 42444 28393 42472 28494
rect 42430 28384 42486 28393
rect 42430 28319 42486 28328
rect 42614 27568 42670 27577
rect 42614 27503 42670 27512
rect 42524 27396 42576 27402
rect 42524 27338 42576 27344
rect 42536 27305 42564 27338
rect 42522 27296 42578 27305
rect 42522 27231 42578 27240
rect 42338 26344 42394 26353
rect 42394 26302 42472 26330
rect 42338 26279 42394 26288
rect 42340 25424 42392 25430
rect 42340 25366 42392 25372
rect 42248 24268 42300 24274
rect 42248 24210 42300 24216
rect 42156 22024 42208 22030
rect 42156 21966 42208 21972
rect 42064 12300 42116 12306
rect 42064 12242 42116 12248
rect 41694 12200 41750 12209
rect 41694 12135 41696 12144
rect 41748 12135 41750 12144
rect 41696 12106 41748 12112
rect 41708 12075 41736 12106
rect 42064 11892 42116 11898
rect 42064 11834 42116 11840
rect 42076 11762 42104 11834
rect 41972 11756 42024 11762
rect 41972 11698 42024 11704
rect 42064 11756 42116 11762
rect 42064 11698 42116 11704
rect 41616 11342 41736 11370
rect 41984 11354 42012 11698
rect 41604 11212 41656 11218
rect 41604 11154 41656 11160
rect 41248 10798 41368 10826
rect 41142 10704 41198 10713
rect 41142 10639 41144 10648
rect 41196 10639 41198 10648
rect 41144 10610 41196 10616
rect 41340 8634 41368 10798
rect 41512 9376 41564 9382
rect 41512 9318 41564 9324
rect 41328 8628 41380 8634
rect 41328 8570 41380 8576
rect 41524 8430 41552 9318
rect 41512 8424 41564 8430
rect 41512 8366 41564 8372
rect 40960 7404 41012 7410
rect 40960 7346 41012 7352
rect 40684 5636 40736 5642
rect 40684 5578 40736 5584
rect 41512 4684 41564 4690
rect 41512 4626 41564 4632
rect 40960 4004 41012 4010
rect 40960 3946 41012 3952
rect 40592 2576 40644 2582
rect 40592 2518 40644 2524
rect 40684 2440 40736 2446
rect 40684 2382 40736 2388
rect 40696 800 40724 2382
rect 40972 800 41000 3946
rect 41144 2984 41196 2990
rect 41144 2926 41196 2932
rect 41156 800 41184 2926
rect 41236 2848 41288 2854
rect 41288 2808 41368 2836
rect 41236 2790 41288 2796
rect 41340 800 41368 2808
rect 41524 800 41552 4626
rect 41616 2922 41644 11154
rect 41708 10713 41736 11342
rect 41972 11348 42024 11354
rect 41972 11290 42024 11296
rect 41694 10704 41750 10713
rect 41694 10639 41750 10648
rect 41708 10470 41736 10639
rect 41788 10600 41840 10606
rect 41786 10568 41788 10577
rect 41840 10568 41842 10577
rect 41786 10503 41842 10512
rect 41696 10464 41748 10470
rect 41696 10406 41748 10412
rect 42168 6934 42196 21966
rect 42248 21616 42300 21622
rect 42248 21558 42300 21564
rect 42260 12646 42288 21558
rect 42248 12640 42300 12646
rect 42248 12582 42300 12588
rect 42248 12300 42300 12306
rect 42248 12242 42300 12248
rect 42260 11898 42288 12242
rect 42248 11892 42300 11898
rect 42248 11834 42300 11840
rect 42156 6928 42208 6934
rect 42156 6870 42208 6876
rect 42156 4480 42208 4486
rect 42156 4422 42208 4428
rect 41696 3596 41748 3602
rect 41696 3538 41748 3544
rect 41604 2916 41656 2922
rect 41604 2858 41656 2864
rect 41708 800 41736 3538
rect 42168 3058 42196 4422
rect 42352 3942 42380 25366
rect 42444 16658 42472 26302
rect 42628 25430 42656 27503
rect 42616 25424 42668 25430
rect 42616 25366 42668 25372
rect 42616 17536 42668 17542
rect 42616 17478 42668 17484
rect 42432 16652 42484 16658
rect 42432 16594 42484 16600
rect 42524 13796 42576 13802
rect 42524 13738 42576 13744
rect 42432 12776 42484 12782
rect 42432 12718 42484 12724
rect 42444 12238 42472 12718
rect 42536 12306 42564 13738
rect 42524 12300 42576 12306
rect 42524 12242 42576 12248
rect 42432 12232 42484 12238
rect 42432 12174 42484 12180
rect 42432 10192 42484 10198
rect 42432 10134 42484 10140
rect 42340 3936 42392 3942
rect 42340 3878 42392 3884
rect 42340 3596 42392 3602
rect 42340 3538 42392 3544
rect 42248 3528 42300 3534
rect 42248 3470 42300 3476
rect 42156 3052 42208 3058
rect 42156 2994 42208 3000
rect 42260 2774 42288 3470
rect 42168 2746 42288 2774
rect 41972 2304 42024 2310
rect 41972 2246 42024 2252
rect 41984 800 42012 2246
rect 42168 800 42196 2746
rect 42248 2508 42300 2514
rect 42248 2450 42300 2456
rect 39764 60 39816 66
rect 39764 2 39816 8
rect 39946 0 40002 800
rect 40130 0 40186 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42260 678 42288 2450
rect 42352 800 42380 3538
rect 42444 3058 42472 10134
rect 42628 9110 42656 17478
rect 42720 12374 42748 32535
rect 42812 29238 42840 32846
rect 42904 31754 42932 37266
rect 42984 35148 43036 35154
rect 42984 35090 43036 35096
rect 42892 31748 42944 31754
rect 42892 31690 42944 31696
rect 42996 30122 43024 35090
rect 42984 30116 43036 30122
rect 42984 30058 43036 30064
rect 42800 29232 42852 29238
rect 42800 29174 42852 29180
rect 42800 27328 42852 27334
rect 42800 27270 42852 27276
rect 42812 24342 42840 27270
rect 42892 26376 42944 26382
rect 42890 26344 42892 26353
rect 42944 26344 42946 26353
rect 42890 26279 42946 26288
rect 42800 24336 42852 24342
rect 42800 24278 42852 24284
rect 42982 23760 43038 23769
rect 42982 23695 42984 23704
rect 43036 23695 43038 23704
rect 42984 23666 43036 23672
rect 42892 21344 42944 21350
rect 42892 21286 42944 21292
rect 42904 21146 42932 21286
rect 42800 21140 42852 21146
rect 42800 21082 42852 21088
rect 42892 21140 42944 21146
rect 42892 21082 42944 21088
rect 42812 20942 42840 21082
rect 42800 20936 42852 20942
rect 42800 20878 42852 20884
rect 42798 18728 42854 18737
rect 42798 18663 42854 18672
rect 42812 17814 42840 18663
rect 42800 17808 42852 17814
rect 42800 17750 42852 17756
rect 42892 15088 42944 15094
rect 42892 15030 42944 15036
rect 42800 13320 42852 13326
rect 42800 13262 42852 13268
rect 42812 12374 42840 13262
rect 42708 12368 42760 12374
rect 42708 12310 42760 12316
rect 42800 12368 42852 12374
rect 42800 12310 42852 12316
rect 42904 12306 42932 15030
rect 43088 14278 43116 37606
rect 43364 37398 43392 39200
rect 43352 37392 43404 37398
rect 43352 37334 43404 37340
rect 43536 36712 43588 36718
rect 43536 36654 43588 36660
rect 43812 36712 43864 36718
rect 43812 36654 43864 36660
rect 43350 36544 43406 36553
rect 43350 36479 43406 36488
rect 43364 36242 43392 36479
rect 43442 36408 43498 36417
rect 43442 36343 43498 36352
rect 43352 36236 43404 36242
rect 43352 36178 43404 36184
rect 43456 36038 43484 36343
rect 43548 36242 43576 36654
rect 43536 36236 43588 36242
rect 43588 36196 43668 36224
rect 43536 36178 43588 36184
rect 43444 36032 43496 36038
rect 43444 35974 43496 35980
rect 43536 35828 43588 35834
rect 43536 35770 43588 35776
rect 43548 35222 43576 35770
rect 43640 35698 43668 36196
rect 43628 35692 43680 35698
rect 43628 35634 43680 35640
rect 43824 35630 43852 36654
rect 44192 35834 44220 39200
rect 44364 37324 44416 37330
rect 44364 37266 44416 37272
rect 44180 35828 44232 35834
rect 44180 35770 44232 35776
rect 43812 35624 43864 35630
rect 43812 35566 43864 35572
rect 43904 35488 43956 35494
rect 43904 35430 43956 35436
rect 43352 35216 43404 35222
rect 43352 35158 43404 35164
rect 43536 35216 43588 35222
rect 43536 35158 43588 35164
rect 43626 35184 43682 35193
rect 43364 34921 43392 35158
rect 43916 35154 43944 35430
rect 44272 35216 44324 35222
rect 44272 35158 44324 35164
rect 43626 35119 43682 35128
rect 43720 35148 43772 35154
rect 43350 34912 43406 34921
rect 43350 34847 43406 34856
rect 43640 34678 43668 35119
rect 43720 35090 43772 35096
rect 43904 35148 43956 35154
rect 43904 35090 43956 35096
rect 43536 34672 43588 34678
rect 43536 34614 43588 34620
rect 43628 34672 43680 34678
rect 43628 34614 43680 34620
rect 43548 34542 43576 34614
rect 43536 34536 43588 34542
rect 43536 34478 43588 34484
rect 43732 33425 43760 35090
rect 43718 33416 43774 33425
rect 43718 33351 43774 33360
rect 43168 32768 43220 32774
rect 43168 32710 43220 32716
rect 43180 32570 43208 32710
rect 43168 32564 43220 32570
rect 43168 32506 43220 32512
rect 43536 31680 43588 31686
rect 43536 31622 43588 31628
rect 43548 31414 43576 31622
rect 43536 31408 43588 31414
rect 43536 31350 43588 31356
rect 43628 31408 43680 31414
rect 43628 31350 43680 31356
rect 43640 31210 43668 31350
rect 43628 31204 43680 31210
rect 43628 31146 43680 31152
rect 43534 30560 43590 30569
rect 43534 30495 43590 30504
rect 43444 30116 43496 30122
rect 43444 30058 43496 30064
rect 43350 30016 43406 30025
rect 43350 29951 43406 29960
rect 43364 29850 43392 29951
rect 43352 29844 43404 29850
rect 43352 29786 43404 29792
rect 43168 29776 43220 29782
rect 43168 29718 43220 29724
rect 43180 19009 43208 29718
rect 43352 29572 43404 29578
rect 43352 29514 43404 29520
rect 43364 29481 43392 29514
rect 43350 29472 43406 29481
rect 43350 29407 43406 29416
rect 43352 27056 43404 27062
rect 43352 26998 43404 27004
rect 43364 26625 43392 26998
rect 43350 26616 43406 26625
rect 43350 26551 43406 26560
rect 43260 26240 43312 26246
rect 43260 26182 43312 26188
rect 43352 26240 43404 26246
rect 43352 26182 43404 26188
rect 43272 25673 43300 26182
rect 43364 25770 43392 26182
rect 43352 25764 43404 25770
rect 43352 25706 43404 25712
rect 43258 25664 43314 25673
rect 43258 25599 43314 25608
rect 43352 25288 43404 25294
rect 43352 25230 43404 25236
rect 43260 24064 43312 24070
rect 43260 24006 43312 24012
rect 43272 23866 43300 24006
rect 43260 23860 43312 23866
rect 43260 23802 43312 23808
rect 43260 23724 43312 23730
rect 43260 23666 43312 23672
rect 43166 19000 43222 19009
rect 43166 18935 43222 18944
rect 43168 14476 43220 14482
rect 43168 14418 43220 14424
rect 43076 14272 43128 14278
rect 43076 14214 43128 14220
rect 42984 13864 43036 13870
rect 43036 13824 43116 13852
rect 42984 13806 43036 13812
rect 42892 12300 42944 12306
rect 42892 12242 42944 12248
rect 42708 12164 42760 12170
rect 42708 12106 42760 12112
rect 42616 9104 42668 9110
rect 42616 9046 42668 9052
rect 42720 7426 42748 12106
rect 42984 12096 43036 12102
rect 42984 12038 43036 12044
rect 42996 11286 43024 12038
rect 42984 11280 43036 11286
rect 42984 11222 43036 11228
rect 42892 10804 42944 10810
rect 42892 10746 42944 10752
rect 42800 10192 42852 10198
rect 42800 10134 42852 10140
rect 42812 9926 42840 10134
rect 42904 9926 42932 10746
rect 42800 9920 42852 9926
rect 42800 9862 42852 9868
rect 42892 9920 42944 9926
rect 42892 9862 42944 9868
rect 43088 8974 43116 13824
rect 43180 12850 43208 14418
rect 43168 12844 43220 12850
rect 43168 12786 43220 12792
rect 43076 8968 43128 8974
rect 43076 8910 43128 8916
rect 42536 7398 42748 7426
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 42536 2774 42564 7398
rect 42708 7336 42760 7342
rect 42708 7278 42760 7284
rect 42720 4214 42748 7278
rect 42800 6248 42852 6254
rect 42800 6190 42852 6196
rect 42812 6118 42840 6190
rect 42800 6112 42852 6118
rect 42800 6054 42852 6060
rect 42708 4208 42760 4214
rect 42708 4150 42760 4156
rect 42708 4072 42760 4078
rect 42708 4014 42760 4020
rect 42444 2746 42564 2774
rect 42444 2582 42472 2746
rect 42432 2576 42484 2582
rect 42432 2518 42484 2524
rect 42524 2508 42576 2514
rect 42524 2450 42576 2456
rect 42536 800 42564 2450
rect 42720 800 42748 4014
rect 42984 3596 43036 3602
rect 42984 3538 43036 3544
rect 42996 800 43024 3538
rect 43076 3460 43128 3466
rect 43076 3402 43128 3408
rect 43088 1290 43116 3402
rect 43168 2848 43220 2854
rect 43168 2790 43220 2796
rect 43076 1284 43128 1290
rect 43076 1226 43128 1232
rect 43180 800 43208 2790
rect 43272 1290 43300 23666
rect 43364 12434 43392 25230
rect 43456 24857 43484 30058
rect 43548 28665 43576 30495
rect 43732 30258 43760 33351
rect 43720 30252 43772 30258
rect 43720 30194 43772 30200
rect 43534 28656 43590 28665
rect 43590 28614 43852 28642
rect 43534 28591 43590 28600
rect 43536 25832 43588 25838
rect 43536 25774 43588 25780
rect 43548 24886 43576 25774
rect 43718 25664 43774 25673
rect 43718 25599 43774 25608
rect 43732 25430 43760 25599
rect 43720 25424 43772 25430
rect 43626 25392 43682 25401
rect 43720 25366 43772 25372
rect 43626 25327 43628 25336
rect 43680 25327 43682 25336
rect 43628 25298 43680 25304
rect 43640 25158 43668 25298
rect 43718 25256 43774 25265
rect 43718 25191 43774 25200
rect 43732 25158 43760 25191
rect 43628 25152 43680 25158
rect 43628 25094 43680 25100
rect 43720 25152 43772 25158
rect 43720 25094 43772 25100
rect 43536 24880 43588 24886
rect 43442 24848 43498 24857
rect 43824 24834 43852 28614
rect 43536 24822 43588 24828
rect 43442 24783 43498 24792
rect 43732 24806 43852 24834
rect 43456 22094 43484 24783
rect 43628 24676 43680 24682
rect 43628 24618 43680 24624
rect 43534 24576 43590 24585
rect 43534 24511 43590 24520
rect 43548 24410 43576 24511
rect 43536 24404 43588 24410
rect 43536 24346 43588 24352
rect 43640 24342 43668 24618
rect 43628 24336 43680 24342
rect 43628 24278 43680 24284
rect 43732 23610 43760 24806
rect 43812 24744 43864 24750
rect 43812 24686 43864 24692
rect 43824 23730 43852 24686
rect 43812 23724 43864 23730
rect 43812 23666 43864 23672
rect 43732 23582 43852 23610
rect 43824 22098 43852 23582
rect 43456 22066 43576 22094
rect 43444 19848 43496 19854
rect 43444 19790 43496 19796
rect 43456 19689 43484 19790
rect 43442 19680 43498 19689
rect 43442 19615 43498 19624
rect 43444 19236 43496 19242
rect 43444 19178 43496 19184
rect 43456 19145 43484 19178
rect 43442 19136 43498 19145
rect 43442 19071 43498 19080
rect 43444 18352 43496 18358
rect 43442 18320 43444 18329
rect 43496 18320 43498 18329
rect 43442 18255 43498 18264
rect 43548 17270 43576 22066
rect 43812 22092 43864 22098
rect 43812 22034 43864 22040
rect 43916 19802 43944 35090
rect 44284 35057 44312 35158
rect 44270 35048 44326 35057
rect 44270 34983 44326 34992
rect 44284 34066 44312 34983
rect 44272 34060 44324 34066
rect 44272 34002 44324 34008
rect 43994 33416 44050 33425
rect 43994 33351 44050 33360
rect 44008 30802 44036 33351
rect 44178 32328 44234 32337
rect 44178 32263 44234 32272
rect 44192 31822 44220 32263
rect 44180 31816 44232 31822
rect 44180 31758 44232 31764
rect 44272 31748 44324 31754
rect 44272 31690 44324 31696
rect 44284 31482 44312 31690
rect 44088 31476 44140 31482
rect 44088 31418 44140 31424
rect 44272 31476 44324 31482
rect 44272 31418 44324 31424
rect 43996 30796 44048 30802
rect 43996 30738 44048 30744
rect 44100 27169 44128 31418
rect 44086 27160 44142 27169
rect 44086 27095 44142 27104
rect 44088 25356 44140 25362
rect 44088 25298 44140 25304
rect 43996 24404 44048 24410
rect 43996 24346 44048 24352
rect 44008 24206 44036 24346
rect 43996 24200 44048 24206
rect 43996 24142 44048 24148
rect 44100 24070 44128 25298
rect 44272 25288 44324 25294
rect 44272 25230 44324 25236
rect 44284 24426 44312 25230
rect 44192 24398 44312 24426
rect 44088 24064 44140 24070
rect 44088 24006 44140 24012
rect 44192 23610 44220 24398
rect 44376 24274 44404 37266
rect 44456 33992 44508 33998
rect 44456 33934 44508 33940
rect 44364 24268 44416 24274
rect 44364 24210 44416 24216
rect 44192 23582 44404 23610
rect 44180 23180 44232 23186
rect 44180 23122 44232 23128
rect 43996 22568 44048 22574
rect 43996 22510 44048 22516
rect 44008 21622 44036 22510
rect 43996 21616 44048 21622
rect 43996 21558 44048 21564
rect 44088 21412 44140 21418
rect 44088 21354 44140 21360
rect 44100 20942 44128 21354
rect 44088 20936 44140 20942
rect 44088 20878 44140 20884
rect 44088 20596 44140 20602
rect 44088 20538 44140 20544
rect 44100 20058 44128 20538
rect 44088 20052 44140 20058
rect 44088 19994 44140 20000
rect 43824 19774 43944 19802
rect 43994 19816 44050 19825
rect 43628 18216 43680 18222
rect 43628 18158 43680 18164
rect 43640 17542 43668 18158
rect 43824 17814 43852 19774
rect 43994 19751 44050 19760
rect 44008 19718 44036 19751
rect 43904 19712 43956 19718
rect 43902 19680 43904 19689
rect 43996 19712 44048 19718
rect 43956 19680 43958 19689
rect 43996 19654 44048 19660
rect 43902 19615 43958 19624
rect 44086 19544 44142 19553
rect 44086 19479 44142 19488
rect 44100 19446 44128 19479
rect 44088 19440 44140 19446
rect 44088 19382 44140 19388
rect 44088 19168 44140 19174
rect 44088 19110 44140 19116
rect 43812 17808 43864 17814
rect 43812 17750 43864 17756
rect 43628 17536 43680 17542
rect 43628 17478 43680 17484
rect 43536 17264 43588 17270
rect 43536 17206 43588 17212
rect 43536 14408 43588 14414
rect 43536 14350 43588 14356
rect 43548 12782 43576 14350
rect 43640 13802 43668 17478
rect 44100 16114 44128 19110
rect 44088 16108 44140 16114
rect 44088 16050 44140 16056
rect 43812 14952 43864 14958
rect 43812 14894 43864 14900
rect 43720 14272 43772 14278
rect 43720 14214 43772 14220
rect 43732 13870 43760 14214
rect 43824 13938 43852 14894
rect 43904 14544 43956 14550
rect 43904 14486 43956 14492
rect 43916 14278 43944 14486
rect 43904 14272 43956 14278
rect 43904 14214 43956 14220
rect 44086 13968 44142 13977
rect 43812 13932 43864 13938
rect 44086 13903 44088 13912
rect 43812 13874 43864 13880
rect 44140 13903 44142 13912
rect 44088 13874 44140 13880
rect 43720 13864 43772 13870
rect 43720 13806 43772 13812
rect 43628 13796 43680 13802
rect 43628 13738 43680 13744
rect 43812 12844 43864 12850
rect 43812 12786 43864 12792
rect 43536 12776 43588 12782
rect 43534 12744 43536 12753
rect 43588 12744 43590 12753
rect 43534 12679 43590 12688
rect 43364 12406 43484 12434
rect 43352 6860 43404 6866
rect 43352 6802 43404 6808
rect 43364 6118 43392 6802
rect 43352 6112 43404 6118
rect 43352 6054 43404 6060
rect 43456 5234 43484 12406
rect 43824 6254 43852 12786
rect 44192 10606 44220 23122
rect 44272 16176 44324 16182
rect 44272 16118 44324 16124
rect 44284 13841 44312 16118
rect 44270 13832 44326 13841
rect 44270 13767 44326 13776
rect 44376 10742 44404 23582
rect 44364 10736 44416 10742
rect 44270 10704 44326 10713
rect 44364 10678 44416 10684
rect 44270 10639 44326 10648
rect 44284 10606 44312 10639
rect 44180 10600 44232 10606
rect 44180 10542 44232 10548
rect 44272 10600 44324 10606
rect 44272 10542 44324 10548
rect 44086 10432 44142 10441
rect 44086 10367 44142 10376
rect 43994 10024 44050 10033
rect 44100 9994 44128 10367
rect 43994 9959 43996 9968
rect 44048 9959 44050 9968
rect 44088 9988 44140 9994
rect 43996 9930 44048 9936
rect 44088 9930 44140 9936
rect 44192 9674 44220 10542
rect 44192 9646 44312 9674
rect 43812 6248 43864 6254
rect 43812 6190 43864 6196
rect 43444 5228 43496 5234
rect 43444 5170 43496 5176
rect 44088 5092 44140 5098
rect 44088 5034 44140 5040
rect 43996 4684 44048 4690
rect 43996 4626 44048 4632
rect 43352 4004 43404 4010
rect 43352 3946 43404 3952
rect 43260 1284 43312 1290
rect 43260 1226 43312 1232
rect 43364 800 43392 3946
rect 43536 2984 43588 2990
rect 43536 2926 43588 2932
rect 43548 800 43576 2926
rect 43628 2916 43680 2922
rect 43628 2858 43680 2864
rect 43640 1358 43668 2858
rect 43812 2372 43864 2378
rect 43812 2314 43864 2320
rect 43628 1352 43680 1358
rect 43628 1294 43680 1300
rect 43824 800 43852 2314
rect 44008 800 44036 4626
rect 44100 2582 44128 5034
rect 44180 2916 44232 2922
rect 44180 2858 44232 2864
rect 44088 2576 44140 2582
rect 44088 2518 44140 2524
rect 44192 800 44220 2858
rect 44284 950 44312 9646
rect 44364 2848 44416 2854
rect 44364 2790 44416 2796
rect 44272 944 44324 950
rect 44272 886 44324 892
rect 44376 800 44404 2790
rect 44468 2582 44496 33934
rect 44548 25356 44600 25362
rect 44548 25298 44600 25304
rect 44560 23186 44588 25298
rect 44640 24880 44692 24886
rect 44638 24848 44640 24857
rect 44692 24848 44694 24857
rect 44638 24783 44694 24792
rect 44744 24750 44772 39306
rect 45098 39200 45154 40000
rect 45926 39200 45982 40000
rect 46480 39364 46532 39370
rect 46480 39306 46532 39312
rect 45112 37330 45140 39200
rect 45284 38004 45336 38010
rect 45284 37946 45336 37952
rect 45296 37466 45324 37946
rect 45940 37466 45968 39200
rect 45284 37460 45336 37466
rect 45284 37402 45336 37408
rect 45928 37460 45980 37466
rect 45928 37402 45980 37408
rect 45100 37324 45152 37330
rect 45100 37266 45152 37272
rect 45100 36576 45152 36582
rect 45100 36518 45152 36524
rect 45112 35698 45140 36518
rect 45100 35692 45152 35698
rect 45100 35634 45152 35640
rect 46112 35624 46164 35630
rect 46164 35584 46428 35612
rect 46112 35566 46164 35572
rect 46400 35494 46428 35584
rect 46388 35488 46440 35494
rect 46388 35430 46440 35436
rect 46492 35306 46520 39306
rect 46846 39200 46902 40000
rect 47674 39200 47730 40000
rect 48594 39200 48650 40000
rect 49422 39200 49478 40000
rect 50342 39200 50398 40000
rect 51262 39200 51318 40000
rect 52090 39200 52146 40000
rect 53010 39200 53066 40000
rect 53838 39200 53894 40000
rect 54758 39200 54814 40000
rect 55496 39432 55548 39438
rect 55496 39374 55548 39380
rect 46860 36938 46888 39200
rect 47688 37398 47716 39200
rect 47860 38072 47912 38078
rect 47860 38014 47912 38020
rect 47872 37466 47900 38014
rect 48412 37868 48464 37874
rect 48412 37810 48464 37816
rect 47860 37460 47912 37466
rect 47860 37402 47912 37408
rect 47676 37392 47728 37398
rect 47676 37334 47728 37340
rect 47952 37324 48004 37330
rect 47952 37266 48004 37272
rect 46860 36922 46980 36938
rect 46860 36916 46992 36922
rect 46860 36910 46940 36916
rect 46940 36858 46992 36864
rect 47308 36780 47360 36786
rect 47308 36722 47360 36728
rect 46664 36576 46716 36582
rect 46664 36518 46716 36524
rect 46572 35692 46624 35698
rect 46572 35634 46624 35640
rect 46400 35278 46520 35306
rect 46584 35290 46612 35634
rect 46676 35630 46704 36518
rect 47320 36394 47348 36722
rect 47400 36712 47452 36718
rect 47400 36654 47452 36660
rect 47412 36417 47440 36654
rect 47766 36544 47822 36553
rect 47766 36479 47822 36488
rect 46952 36366 47348 36394
rect 47398 36408 47454 36417
rect 46952 36310 46980 36366
rect 47398 36343 47454 36352
rect 46940 36304 46992 36310
rect 46940 36246 46992 36252
rect 47044 36230 47624 36258
rect 47780 36242 47808 36479
rect 46940 36168 46992 36174
rect 47044 36156 47072 36230
rect 47596 36174 47624 36230
rect 47768 36236 47820 36242
rect 47768 36178 47820 36184
rect 46992 36128 47072 36156
rect 47400 36168 47452 36174
rect 46940 36110 46992 36116
rect 47400 36110 47452 36116
rect 47584 36168 47636 36174
rect 47584 36110 47636 36116
rect 47124 36100 47176 36106
rect 47124 36042 47176 36048
rect 47136 35850 47164 36042
rect 47412 35850 47440 36110
rect 47136 35822 47440 35850
rect 46756 35760 46808 35766
rect 46754 35728 46756 35737
rect 46808 35728 46810 35737
rect 46754 35663 46810 35672
rect 46664 35624 46716 35630
rect 46664 35566 46716 35572
rect 47306 35320 47362 35329
rect 46572 35284 46624 35290
rect 45466 34096 45522 34105
rect 45466 34031 45522 34040
rect 45480 33998 45508 34031
rect 45468 33992 45520 33998
rect 45468 33934 45520 33940
rect 45560 33992 45612 33998
rect 45560 33934 45612 33940
rect 45572 33522 45600 33934
rect 45560 33516 45612 33522
rect 45560 33458 45612 33464
rect 45652 33516 45704 33522
rect 45652 33458 45704 33464
rect 45466 33008 45522 33017
rect 45466 32943 45522 32952
rect 45100 30592 45152 30598
rect 45100 30534 45152 30540
rect 44732 24744 44784 24750
rect 44732 24686 44784 24692
rect 44916 24744 44968 24750
rect 44916 24686 44968 24692
rect 44732 24268 44784 24274
rect 44732 24210 44784 24216
rect 44548 23180 44600 23186
rect 44548 23122 44600 23128
rect 44548 21616 44600 21622
rect 44548 21558 44600 21564
rect 44560 21457 44588 21558
rect 44546 21448 44602 21457
rect 44546 21383 44602 21392
rect 44548 20936 44600 20942
rect 44548 20878 44600 20884
rect 44560 18970 44588 20878
rect 44640 20596 44692 20602
rect 44640 20538 44692 20544
rect 44652 20262 44680 20538
rect 44640 20256 44692 20262
rect 44640 20198 44692 20204
rect 44640 19168 44692 19174
rect 44640 19110 44692 19116
rect 44652 19009 44680 19110
rect 44638 19000 44694 19009
rect 44548 18964 44600 18970
rect 44638 18935 44694 18944
rect 44548 18906 44600 18912
rect 44560 18601 44588 18906
rect 44546 18592 44602 18601
rect 44546 18527 44602 18536
rect 44652 16810 44680 18935
rect 44744 18737 44772 24210
rect 44822 19544 44878 19553
rect 44822 19479 44878 19488
rect 44730 18728 44786 18737
rect 44730 18663 44786 18672
rect 44560 16782 44680 16810
rect 44560 9674 44588 16782
rect 44744 16708 44772 18663
rect 44652 16680 44772 16708
rect 44652 13258 44680 16680
rect 44836 16590 44864 19479
rect 44824 16584 44876 16590
rect 44824 16526 44876 16532
rect 44640 13252 44692 13258
rect 44640 13194 44692 13200
rect 44640 12640 44692 12646
rect 44640 12582 44692 12588
rect 44652 12306 44680 12582
rect 44640 12300 44692 12306
rect 44640 12242 44692 12248
rect 44824 12300 44876 12306
rect 44824 12242 44876 12248
rect 44640 10804 44692 10810
rect 44640 10746 44692 10752
rect 44652 10577 44680 10746
rect 44638 10568 44694 10577
rect 44638 10503 44694 10512
rect 44560 9646 44680 9674
rect 44548 4684 44600 4690
rect 44548 4626 44600 4632
rect 44456 2576 44508 2582
rect 44456 2518 44508 2524
rect 44560 800 44588 4626
rect 44652 3670 44680 9646
rect 44732 9036 44784 9042
rect 44732 8978 44784 8984
rect 44640 3664 44692 3670
rect 44640 3606 44692 3612
rect 44744 2650 44772 8978
rect 44836 6662 44864 12242
rect 44928 9518 44956 24686
rect 45008 23792 45060 23798
rect 45008 23734 45060 23740
rect 44916 9512 44968 9518
rect 44916 9454 44968 9460
rect 45020 8838 45048 23734
rect 45112 20262 45140 30534
rect 45284 30048 45336 30054
rect 45284 29990 45336 29996
rect 45192 23860 45244 23866
rect 45192 23802 45244 23808
rect 45100 20256 45152 20262
rect 45100 20198 45152 20204
rect 45100 19440 45152 19446
rect 45098 19408 45100 19417
rect 45152 19408 45154 19417
rect 45098 19343 45154 19352
rect 45100 17060 45152 17066
rect 45100 17002 45152 17008
rect 45112 10810 45140 17002
rect 45204 13802 45232 23802
rect 45296 20398 45324 29990
rect 45376 26376 45428 26382
rect 45376 26318 45428 26324
rect 45388 24206 45416 26318
rect 45480 24750 45508 32943
rect 45664 29782 45692 33458
rect 45836 31748 45888 31754
rect 45836 31690 45888 31696
rect 45848 30666 45876 31690
rect 46294 30832 46350 30841
rect 46020 30796 46072 30802
rect 46294 30767 46350 30776
rect 46020 30738 46072 30744
rect 45836 30660 45888 30666
rect 45836 30602 45888 30608
rect 45926 29880 45982 29889
rect 45926 29815 45982 29824
rect 45652 29776 45704 29782
rect 45652 29718 45704 29724
rect 45834 29744 45890 29753
rect 45744 29708 45796 29714
rect 45834 29679 45890 29688
rect 45744 29650 45796 29656
rect 45560 25968 45612 25974
rect 45560 25910 45612 25916
rect 45652 25968 45704 25974
rect 45652 25910 45704 25916
rect 45468 24744 45520 24750
rect 45468 24686 45520 24692
rect 45376 24200 45428 24206
rect 45376 24142 45428 24148
rect 45376 23792 45428 23798
rect 45374 23760 45376 23769
rect 45428 23760 45430 23769
rect 45374 23695 45430 23704
rect 45480 22094 45508 24686
rect 45388 22066 45508 22094
rect 45284 20392 45336 20398
rect 45284 20334 45336 20340
rect 45284 20256 45336 20262
rect 45284 20198 45336 20204
rect 45296 17270 45324 20198
rect 45284 17264 45336 17270
rect 45284 17206 45336 17212
rect 45284 16584 45336 16590
rect 45284 16526 45336 16532
rect 45192 13796 45244 13802
rect 45192 13738 45244 13744
rect 45192 13524 45244 13530
rect 45192 13466 45244 13472
rect 45100 10804 45152 10810
rect 45100 10746 45152 10752
rect 45204 10606 45232 13466
rect 45192 10600 45244 10606
rect 45192 10542 45244 10548
rect 45008 8832 45060 8838
rect 45008 8774 45060 8780
rect 44824 6656 44876 6662
rect 44824 6598 44876 6604
rect 44916 5772 44968 5778
rect 44916 5714 44968 5720
rect 44824 3596 44876 3602
rect 44824 3538 44876 3544
rect 44732 2644 44784 2650
rect 44732 2586 44784 2592
rect 44836 800 44864 3538
rect 42248 672 42300 678
rect 42248 614 42300 620
rect 42338 0 42394 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 44928 610 44956 5714
rect 45020 5234 45048 8774
rect 45296 7478 45324 16526
rect 45388 15570 45416 22066
rect 45468 20392 45520 20398
rect 45468 20334 45520 20340
rect 45480 19922 45508 20334
rect 45468 19916 45520 19922
rect 45468 19858 45520 19864
rect 45468 19372 45520 19378
rect 45468 19314 45520 19320
rect 45480 18970 45508 19314
rect 45468 18964 45520 18970
rect 45468 18906 45520 18912
rect 45466 17912 45522 17921
rect 45466 17847 45522 17856
rect 45480 17814 45508 17847
rect 45572 17814 45600 25910
rect 45664 25294 45692 25910
rect 45652 25288 45704 25294
rect 45652 25230 45704 25236
rect 45756 25106 45784 29650
rect 45848 29578 45876 29679
rect 45836 29572 45888 29578
rect 45836 29514 45888 29520
rect 45836 29096 45888 29102
rect 45836 29038 45888 29044
rect 45848 26382 45876 29038
rect 45836 26376 45888 26382
rect 45836 26318 45888 26324
rect 45664 25078 45784 25106
rect 45468 17808 45520 17814
rect 45468 17750 45520 17756
rect 45560 17808 45612 17814
rect 45560 17750 45612 17756
rect 45560 17128 45612 17134
rect 45560 17070 45612 17076
rect 45376 15564 45428 15570
rect 45376 15506 45428 15512
rect 45468 12096 45520 12102
rect 45468 12038 45520 12044
rect 45376 10736 45428 10742
rect 45376 10678 45428 10684
rect 45388 10198 45416 10678
rect 45376 10192 45428 10198
rect 45376 10134 45428 10140
rect 45376 7744 45428 7750
rect 45376 7686 45428 7692
rect 45284 7472 45336 7478
rect 45284 7414 45336 7420
rect 45100 6928 45152 6934
rect 45100 6870 45152 6876
rect 45008 5228 45060 5234
rect 45008 5170 45060 5176
rect 45112 3670 45140 6870
rect 45296 5234 45324 7414
rect 45388 6934 45416 7686
rect 45480 7478 45508 12038
rect 45572 7750 45600 17070
rect 45664 12306 45692 25078
rect 45940 24732 45968 29815
rect 46032 27713 46060 30738
rect 46308 30734 46336 30767
rect 46296 30728 46348 30734
rect 46296 30670 46348 30676
rect 46110 30152 46166 30161
rect 46110 30087 46166 30096
rect 46124 29034 46152 30087
rect 46204 29640 46256 29646
rect 46204 29582 46256 29588
rect 46216 29238 46244 29582
rect 46204 29232 46256 29238
rect 46204 29174 46256 29180
rect 46112 29028 46164 29034
rect 46112 28970 46164 28976
rect 46204 29028 46256 29034
rect 46204 28970 46256 28976
rect 46018 27704 46074 27713
rect 46018 27639 46074 27648
rect 45756 24704 45968 24732
rect 45652 12300 45704 12306
rect 45652 12242 45704 12248
rect 45652 12096 45704 12102
rect 45652 12038 45704 12044
rect 45664 11830 45692 12038
rect 45652 11824 45704 11830
rect 45652 11766 45704 11772
rect 45560 7744 45612 7750
rect 45560 7686 45612 7692
rect 45468 7472 45520 7478
rect 45468 7414 45520 7420
rect 45376 6928 45428 6934
rect 45376 6870 45428 6876
rect 45468 6656 45520 6662
rect 45468 6598 45520 6604
rect 45284 5228 45336 5234
rect 45284 5170 45336 5176
rect 45376 4072 45428 4078
rect 45376 4014 45428 4020
rect 45192 4004 45244 4010
rect 45192 3946 45244 3952
rect 45100 3664 45152 3670
rect 45100 3606 45152 3612
rect 45008 2440 45060 2446
rect 45008 2382 45060 2388
rect 45020 800 45048 2382
rect 45204 800 45232 3946
rect 45388 800 45416 4014
rect 45480 2310 45508 6598
rect 45756 2990 45784 24704
rect 45836 24200 45888 24206
rect 45836 24142 45888 24148
rect 46032 24154 46060 27639
rect 46124 27010 46152 28970
rect 46216 28762 46244 28970
rect 46204 28756 46256 28762
rect 46204 28698 46256 28704
rect 46296 28552 46348 28558
rect 46296 28494 46348 28500
rect 46308 28150 46336 28494
rect 46204 28144 46256 28150
rect 46204 28086 46256 28092
rect 46296 28144 46348 28150
rect 46296 28086 46348 28092
rect 46216 27674 46244 28086
rect 46204 27668 46256 27674
rect 46204 27610 46256 27616
rect 46204 27464 46256 27470
rect 46204 27406 46256 27412
rect 46216 27130 46244 27406
rect 46294 27160 46350 27169
rect 46204 27124 46256 27130
rect 46294 27095 46296 27104
rect 46204 27066 46256 27072
rect 46348 27095 46350 27104
rect 46296 27066 46348 27072
rect 46124 26982 46244 27010
rect 46112 24676 46164 24682
rect 46112 24618 46164 24624
rect 46124 24342 46152 24618
rect 46112 24336 46164 24342
rect 46112 24278 46164 24284
rect 45848 19310 45876 24142
rect 46032 24126 46152 24154
rect 46020 22976 46072 22982
rect 46020 22918 46072 22924
rect 45928 21004 45980 21010
rect 45928 20946 45980 20952
rect 45940 20874 45968 20946
rect 45928 20868 45980 20874
rect 45928 20810 45980 20816
rect 45926 19680 45982 19689
rect 45926 19615 45982 19624
rect 45836 19304 45888 19310
rect 45836 19246 45888 19252
rect 45836 18216 45888 18222
rect 45836 18158 45888 18164
rect 45848 15094 45876 18158
rect 45836 15088 45888 15094
rect 45836 15030 45888 15036
rect 45940 13462 45968 19615
rect 46032 18222 46060 22918
rect 46124 21010 46152 24126
rect 46216 23730 46244 26982
rect 46400 24342 46428 35278
rect 47306 35255 47362 35264
rect 46572 35226 46624 35232
rect 47320 35154 47348 35255
rect 46756 35148 46808 35154
rect 46756 35090 46808 35096
rect 47124 35148 47176 35154
rect 47124 35090 47176 35096
rect 47308 35148 47360 35154
rect 47308 35090 47360 35096
rect 46478 33824 46534 33833
rect 46478 33759 46534 33768
rect 46492 24342 46520 33759
rect 46570 32872 46626 32881
rect 46570 32807 46572 32816
rect 46624 32807 46626 32816
rect 46572 32778 46624 32784
rect 46572 32224 46624 32230
rect 46572 32166 46624 32172
rect 46584 29850 46612 32166
rect 46768 31754 46796 35090
rect 46860 34598 47072 34626
rect 46860 34542 46888 34598
rect 46848 34536 46900 34542
rect 46848 34478 46900 34484
rect 46940 34536 46992 34542
rect 46940 34478 46992 34484
rect 46952 34134 46980 34478
rect 46940 34128 46992 34134
rect 46940 34070 46992 34076
rect 47044 32230 47072 34598
rect 47032 32224 47084 32230
rect 47032 32166 47084 32172
rect 46768 31726 46888 31754
rect 46664 30796 46716 30802
rect 46664 30738 46716 30744
rect 46676 30569 46704 30738
rect 46756 30728 46808 30734
rect 46756 30670 46808 30676
rect 46662 30560 46718 30569
rect 46662 30495 46718 30504
rect 46662 30152 46718 30161
rect 46662 30087 46718 30096
rect 46572 29844 46624 29850
rect 46572 29786 46624 29792
rect 46388 24336 46440 24342
rect 46388 24278 46440 24284
rect 46480 24336 46532 24342
rect 46480 24278 46532 24284
rect 46296 24268 46348 24274
rect 46296 24210 46348 24216
rect 46204 23724 46256 23730
rect 46204 23666 46256 23672
rect 46308 22094 46336 24210
rect 46584 24154 46612 29786
rect 46676 29782 46704 30087
rect 46664 29776 46716 29782
rect 46664 29718 46716 29724
rect 46664 29640 46716 29646
rect 46664 29582 46716 29588
rect 46676 29510 46704 29582
rect 46664 29504 46716 29510
rect 46664 29446 46716 29452
rect 46664 26512 46716 26518
rect 46664 26454 46716 26460
rect 46676 26353 46704 26454
rect 46662 26344 46718 26353
rect 46662 26279 46718 26288
rect 46662 24440 46718 24449
rect 46662 24375 46718 24384
rect 46676 24342 46704 24375
rect 46664 24336 46716 24342
rect 46664 24278 46716 24284
rect 46388 24132 46440 24138
rect 46388 24074 46440 24080
rect 46492 24126 46612 24154
rect 46662 24168 46718 24177
rect 46400 22982 46428 24074
rect 46388 22976 46440 22982
rect 46388 22918 46440 22924
rect 46308 22066 46428 22094
rect 46204 22024 46256 22030
rect 46204 21966 46256 21972
rect 46296 22024 46348 22030
rect 46296 21966 46348 21972
rect 46216 21486 46244 21966
rect 46308 21894 46336 21966
rect 46296 21888 46348 21894
rect 46296 21830 46348 21836
rect 46204 21480 46256 21486
rect 46204 21422 46256 21428
rect 46112 21004 46164 21010
rect 46112 20946 46164 20952
rect 46112 20596 46164 20602
rect 46112 20538 46164 20544
rect 46124 19666 46152 20538
rect 46211 20256 46263 20262
rect 46211 20198 46263 20204
rect 46216 20182 46251 20198
rect 46216 19786 46244 20182
rect 46204 19780 46256 19786
rect 46204 19722 46256 19728
rect 46296 19780 46348 19786
rect 46296 19722 46348 19728
rect 46308 19666 46336 19722
rect 46124 19638 46336 19666
rect 46112 19440 46164 19446
rect 46110 19408 46112 19417
rect 46164 19408 46166 19417
rect 46110 19343 46166 19352
rect 46204 19304 46256 19310
rect 46204 19246 46256 19252
rect 46110 18864 46166 18873
rect 46110 18799 46166 18808
rect 46124 18222 46152 18799
rect 46020 18216 46072 18222
rect 46020 18158 46072 18164
rect 46112 18216 46164 18222
rect 46112 18158 46164 18164
rect 46110 18048 46166 18057
rect 46110 17983 46166 17992
rect 46124 14958 46152 17983
rect 46112 14952 46164 14958
rect 46112 14894 46164 14900
rect 46020 13864 46072 13870
rect 46020 13806 46072 13812
rect 45928 13456 45980 13462
rect 45928 13398 45980 13404
rect 46032 12170 46060 13806
rect 46216 12753 46244 19246
rect 46294 19000 46350 19009
rect 46294 18935 46296 18944
rect 46348 18935 46350 18944
rect 46296 18906 46348 18912
rect 46400 18057 46428 22066
rect 46386 18048 46442 18057
rect 46386 17983 46442 17992
rect 46386 17912 46442 17921
rect 46386 17847 46442 17856
rect 46400 17814 46428 17847
rect 46296 17808 46348 17814
rect 46296 17750 46348 17756
rect 46388 17808 46440 17814
rect 46388 17750 46440 17756
rect 46308 17134 46336 17750
rect 46388 17196 46440 17202
rect 46388 17138 46440 17144
rect 46296 17128 46348 17134
rect 46296 17070 46348 17076
rect 46400 16726 46428 17138
rect 46388 16720 46440 16726
rect 46388 16662 46440 16668
rect 46388 14544 46440 14550
rect 46388 14486 46440 14492
rect 46400 13870 46428 14486
rect 46388 13864 46440 13870
rect 46388 13806 46440 13812
rect 46388 13184 46440 13190
rect 46388 13126 46440 13132
rect 46400 12850 46428 13126
rect 46388 12844 46440 12850
rect 46388 12786 46440 12792
rect 46202 12744 46258 12753
rect 46202 12679 46258 12688
rect 46216 12238 46244 12679
rect 46204 12232 46256 12238
rect 46204 12174 46256 12180
rect 46020 12164 46072 12170
rect 46020 12106 46072 12112
rect 46204 11824 46256 11830
rect 46204 11766 46256 11772
rect 46216 10266 46244 11766
rect 46388 10804 46440 10810
rect 46388 10746 46440 10752
rect 46296 10668 46348 10674
rect 46296 10610 46348 10616
rect 46204 10260 46256 10266
rect 46204 10202 46256 10208
rect 46308 10198 46336 10610
rect 46296 10192 46348 10198
rect 46296 10134 46348 10140
rect 46204 8288 46256 8294
rect 46204 8230 46256 8236
rect 46216 8090 46244 8230
rect 46204 8084 46256 8090
rect 46204 8026 46256 8032
rect 46296 8084 46348 8090
rect 46296 8026 46348 8032
rect 46204 7948 46256 7954
rect 46308 7936 46336 8026
rect 46256 7908 46336 7936
rect 46204 7890 46256 7896
rect 46112 7880 46164 7886
rect 46112 7822 46164 7828
rect 46124 7002 46152 7822
rect 46296 7200 46348 7206
rect 46296 7142 46348 7148
rect 46020 6996 46072 7002
rect 46020 6938 46072 6944
rect 46112 6996 46164 7002
rect 46112 6938 46164 6944
rect 46032 6882 46060 6938
rect 46308 6882 46336 7142
rect 46032 6854 46336 6882
rect 46204 5568 46256 5574
rect 46204 5510 46256 5516
rect 45836 4684 45888 4690
rect 45836 4626 45888 4632
rect 45744 2984 45796 2990
rect 45744 2926 45796 2932
rect 45560 2916 45612 2922
rect 45560 2858 45612 2864
rect 45468 2304 45520 2310
rect 45468 2246 45520 2252
rect 45572 800 45600 2858
rect 45848 800 45876 4626
rect 46020 4072 46072 4078
rect 46020 4014 46072 4020
rect 46032 800 46060 4014
rect 46216 2990 46244 5510
rect 46296 5296 46348 5302
rect 46296 5238 46348 5244
rect 46308 4282 46336 5238
rect 46400 4486 46428 10746
rect 46492 10266 46520 24126
rect 46662 24103 46718 24112
rect 46676 24018 46704 24103
rect 46584 23990 46704 24018
rect 46584 17678 46612 23990
rect 46664 23724 46716 23730
rect 46664 23666 46716 23672
rect 46572 17672 46624 17678
rect 46572 17614 46624 17620
rect 46572 17196 46624 17202
rect 46572 17138 46624 17144
rect 46584 16590 46612 17138
rect 46572 16584 46624 16590
rect 46572 16526 46624 16532
rect 46570 16416 46626 16425
rect 46570 16351 46626 16360
rect 46584 12714 46612 16351
rect 46572 12708 46624 12714
rect 46572 12650 46624 12656
rect 46676 12238 46704 23666
rect 46768 22098 46796 30670
rect 46860 28121 46888 31726
rect 47032 30796 47084 30802
rect 47032 30738 47084 30744
rect 47044 30598 47072 30738
rect 47032 30592 47084 30598
rect 47032 30534 47084 30540
rect 46938 30016 46994 30025
rect 46938 29951 46994 29960
rect 46952 29850 46980 29951
rect 46940 29844 46992 29850
rect 46940 29786 46992 29792
rect 46940 29708 46992 29714
rect 46940 29650 46992 29656
rect 46952 29238 46980 29650
rect 46940 29232 46992 29238
rect 46940 29174 46992 29180
rect 47044 28762 47072 30534
rect 47032 28756 47084 28762
rect 47032 28698 47084 28704
rect 46846 28112 46902 28121
rect 46846 28047 46902 28056
rect 46860 24449 46888 28047
rect 47030 24712 47086 24721
rect 47030 24647 47086 24656
rect 46938 24576 46994 24585
rect 46938 24511 46994 24520
rect 46846 24440 46902 24449
rect 46952 24410 46980 24511
rect 46846 24375 46902 24384
rect 46940 24404 46992 24410
rect 46940 24346 46992 24352
rect 46940 24132 46992 24138
rect 46940 24074 46992 24080
rect 46952 24041 46980 24074
rect 46938 24032 46994 24041
rect 46938 23967 46994 23976
rect 47044 23662 47072 24647
rect 47032 23656 47084 23662
rect 47032 23598 47084 23604
rect 46848 23112 46900 23118
rect 46848 23054 46900 23060
rect 46860 22982 46888 23054
rect 46848 22976 46900 22982
rect 46848 22918 46900 22924
rect 46848 22160 46900 22166
rect 46848 22102 46900 22108
rect 46756 22092 46808 22098
rect 46756 22034 46808 22040
rect 46664 12232 46716 12238
rect 46664 12174 46716 12180
rect 46664 12096 46716 12102
rect 46768 12050 46796 22034
rect 46860 16425 46888 22102
rect 47136 22094 47164 35090
rect 47308 34128 47360 34134
rect 47306 34096 47308 34105
rect 47360 34096 47362 34105
rect 47306 34031 47362 34040
rect 47306 33144 47362 33153
rect 47306 33079 47362 33088
rect 47214 33008 47270 33017
rect 47214 32943 47270 32952
rect 47228 32910 47256 32943
rect 47320 32910 47348 33079
rect 47216 32904 47268 32910
rect 47216 32846 47268 32852
rect 47308 32904 47360 32910
rect 47308 32846 47360 32852
rect 47214 30832 47270 30841
rect 47214 30767 47270 30776
rect 47228 30598 47256 30767
rect 47308 30728 47360 30734
rect 47308 30670 47360 30676
rect 47216 30592 47268 30598
rect 47216 30534 47268 30540
rect 47320 30054 47348 30670
rect 47216 30048 47268 30054
rect 47216 29990 47268 29996
rect 47308 30048 47360 30054
rect 47308 29990 47360 29996
rect 47228 29782 47256 29990
rect 47216 29776 47268 29782
rect 47216 29718 47268 29724
rect 47306 29744 47362 29753
rect 47306 29679 47362 29688
rect 47320 29646 47348 29679
rect 47308 29640 47360 29646
rect 47308 29582 47360 29588
rect 47216 29504 47268 29510
rect 47214 29472 47216 29481
rect 47268 29472 47270 29481
rect 47214 29407 47270 29416
rect 47308 24744 47360 24750
rect 47308 24686 47360 24692
rect 47320 24274 47348 24686
rect 47308 24268 47360 24274
rect 47308 24210 47360 24216
rect 47306 23080 47362 23089
rect 47306 23015 47308 23024
rect 47360 23015 47362 23024
rect 47308 22986 47360 22992
rect 47044 22066 47164 22094
rect 46940 20868 46992 20874
rect 46940 20810 46992 20816
rect 46952 20466 46980 20810
rect 46940 20460 46992 20466
rect 46940 20402 46992 20408
rect 46940 19916 46992 19922
rect 46940 19858 46992 19864
rect 46952 19553 46980 19858
rect 46938 19544 46994 19553
rect 46938 19479 46994 19488
rect 46940 19304 46992 19310
rect 46940 19246 46992 19252
rect 46952 18465 46980 19246
rect 46938 18456 46994 18465
rect 46938 18391 46994 18400
rect 46938 16688 46994 16697
rect 46938 16623 46940 16632
rect 46992 16623 46994 16632
rect 46940 16594 46992 16600
rect 46846 16416 46902 16425
rect 46846 16351 46902 16360
rect 47044 14006 47072 22066
rect 47122 19136 47178 19145
rect 47122 19071 47178 19080
rect 47136 18630 47164 19071
rect 47308 18828 47360 18834
rect 47308 18770 47360 18776
rect 47124 18624 47176 18630
rect 47124 18566 47176 18572
rect 47214 14376 47270 14385
rect 47214 14311 47270 14320
rect 47032 14000 47084 14006
rect 47032 13942 47084 13948
rect 47044 12288 47072 13942
rect 47228 12374 47256 14311
rect 47216 12368 47268 12374
rect 47216 12310 47268 12316
rect 47124 12300 47176 12306
rect 47044 12260 47124 12288
rect 47124 12242 47176 12248
rect 47320 12170 47348 18770
rect 47308 12164 47360 12170
rect 47308 12106 47360 12112
rect 46716 12044 46796 12050
rect 46664 12038 46796 12044
rect 46848 12096 46900 12102
rect 46848 12038 46900 12044
rect 46676 12022 46796 12038
rect 46860 11898 46888 12038
rect 46848 11892 46900 11898
rect 46848 11834 46900 11840
rect 46570 10704 46626 10713
rect 46570 10639 46572 10648
rect 46624 10639 46626 10648
rect 46572 10610 46624 10616
rect 46480 10260 46532 10266
rect 46480 10202 46532 10208
rect 46662 10024 46718 10033
rect 46662 9959 46718 9968
rect 46480 8628 46532 8634
rect 46480 8570 46532 8576
rect 46492 7886 46520 8570
rect 46480 7880 46532 7886
rect 46480 7822 46532 7828
rect 46480 7744 46532 7750
rect 46480 7686 46532 7692
rect 46572 7744 46624 7750
rect 46572 7686 46624 7692
rect 46388 4480 46440 4486
rect 46388 4422 46440 4428
rect 46296 4276 46348 4282
rect 46296 4218 46348 4224
rect 46388 4004 46440 4010
rect 46388 3946 46440 3952
rect 46204 2984 46256 2990
rect 46204 2926 46256 2932
rect 46112 2848 46164 2854
rect 46112 2790 46164 2796
rect 46204 2848 46256 2854
rect 46204 2790 46256 2796
rect 46124 2650 46152 2790
rect 46112 2644 46164 2650
rect 46112 2586 46164 2592
rect 46216 800 46244 2790
rect 46400 800 46428 3946
rect 46492 1329 46520 7686
rect 46584 7342 46612 7686
rect 46572 7336 46624 7342
rect 46572 7278 46624 7284
rect 46572 3596 46624 3602
rect 46572 3538 46624 3544
rect 46478 1320 46534 1329
rect 46478 1255 46534 1264
rect 46584 800 46612 3538
rect 46676 950 46704 9959
rect 47412 7857 47440 35822
rect 47492 35692 47544 35698
rect 47492 35634 47544 35640
rect 47504 35154 47532 35634
rect 47492 35148 47544 35154
rect 47492 35090 47544 35096
rect 47584 30660 47636 30666
rect 47584 30602 47636 30608
rect 47596 29889 47624 30602
rect 47582 29880 47638 29889
rect 47582 29815 47638 29824
rect 47584 26444 47636 26450
rect 47584 26386 47636 26392
rect 47596 25430 47624 26386
rect 47584 25424 47636 25430
rect 47584 25366 47636 25372
rect 47492 25152 47544 25158
rect 47492 25094 47544 25100
rect 47504 23186 47532 25094
rect 47492 23180 47544 23186
rect 47492 23122 47544 23128
rect 47492 15632 47544 15638
rect 47492 15574 47544 15580
rect 47504 8498 47532 15574
rect 47596 8906 47624 25366
rect 47676 23112 47728 23118
rect 47676 23054 47728 23060
rect 47688 22778 47716 23054
rect 47676 22772 47728 22778
rect 47676 22714 47728 22720
rect 47676 21140 47728 21146
rect 47676 21082 47728 21088
rect 47584 8900 47636 8906
rect 47584 8842 47636 8848
rect 47688 8634 47716 21082
rect 47964 20874 47992 37266
rect 48320 37120 48372 37126
rect 48320 37062 48372 37068
rect 48332 36650 48360 37062
rect 48228 36644 48280 36650
rect 48228 36586 48280 36592
rect 48320 36644 48372 36650
rect 48320 36586 48372 36592
rect 48240 35834 48268 36586
rect 48424 36281 48452 37810
rect 48504 37664 48556 37670
rect 48504 37606 48556 37612
rect 48516 37398 48544 37606
rect 48608 37466 48636 39200
rect 48688 38956 48740 38962
rect 48688 38898 48740 38904
rect 48596 37460 48648 37466
rect 48596 37402 48648 37408
rect 48504 37392 48556 37398
rect 48504 37334 48556 37340
rect 48504 37120 48556 37126
rect 48504 37062 48556 37068
rect 48516 36961 48544 37062
rect 48502 36952 48558 36961
rect 48502 36887 48558 36896
rect 48410 36272 48466 36281
rect 48700 36242 48728 38898
rect 49436 37398 49464 39200
rect 50068 38956 50120 38962
rect 50068 38898 50120 38904
rect 49424 37392 49476 37398
rect 49424 37334 49476 37340
rect 49700 37324 49752 37330
rect 49884 37324 49936 37330
rect 49752 37284 49832 37312
rect 49700 37266 49752 37272
rect 49698 36680 49754 36689
rect 49698 36615 49754 36624
rect 48410 36207 48466 36216
rect 48688 36236 48740 36242
rect 48688 36178 48740 36184
rect 49608 36236 49660 36242
rect 49608 36178 49660 36184
rect 48412 36100 48464 36106
rect 48412 36042 48464 36048
rect 48136 35828 48188 35834
rect 48136 35770 48188 35776
rect 48228 35828 48280 35834
rect 48228 35770 48280 35776
rect 48148 35714 48176 35770
rect 48148 35698 48360 35714
rect 48148 35692 48372 35698
rect 48148 35686 48320 35692
rect 48320 35634 48372 35640
rect 48424 31793 48452 36042
rect 48596 36032 48648 36038
rect 48594 36000 48596 36009
rect 48648 36000 48650 36009
rect 48594 35935 48650 35944
rect 49620 33640 49648 36178
rect 49712 34678 49740 36615
rect 49804 34678 49832 37284
rect 49884 37266 49936 37272
rect 49896 35698 49924 37266
rect 49884 35692 49936 35698
rect 49884 35634 49936 35640
rect 49882 35048 49938 35057
rect 49882 34983 49938 34992
rect 49700 34672 49752 34678
rect 49700 34614 49752 34620
rect 49792 34672 49844 34678
rect 49792 34614 49844 34620
rect 49620 33612 49740 33640
rect 49148 33516 49200 33522
rect 49200 33476 49648 33504
rect 49148 33458 49200 33464
rect 49056 33448 49108 33454
rect 49056 33390 49108 33396
rect 49068 33017 49096 33390
rect 49620 33386 49648 33476
rect 49516 33380 49568 33386
rect 49516 33322 49568 33328
rect 49608 33380 49660 33386
rect 49608 33322 49660 33328
rect 49332 33040 49384 33046
rect 49054 33008 49110 33017
rect 49332 32982 49384 32988
rect 49054 32943 49110 32952
rect 48410 31784 48466 31793
rect 48410 31719 48466 31728
rect 48424 31686 48452 31719
rect 48412 31680 48464 31686
rect 48412 31622 48464 31628
rect 49344 31414 49372 32982
rect 49332 31408 49384 31414
rect 49332 31350 49384 31356
rect 49148 30592 49200 30598
rect 49148 30534 49200 30540
rect 48136 30048 48188 30054
rect 48136 29990 48188 29996
rect 48044 28688 48096 28694
rect 48044 28630 48096 28636
rect 48056 28422 48084 28630
rect 48044 28416 48096 28422
rect 48044 28358 48096 28364
rect 48044 26376 48096 26382
rect 48044 26318 48096 26324
rect 48056 26217 48084 26318
rect 48042 26208 48098 26217
rect 48042 26143 48098 26152
rect 48148 24342 48176 29990
rect 48780 29640 48832 29646
rect 48780 29582 48832 29588
rect 48686 27432 48742 27441
rect 48686 27367 48742 27376
rect 48228 26920 48280 26926
rect 48228 26862 48280 26868
rect 48412 26920 48464 26926
rect 48412 26862 48464 26868
rect 48240 26450 48268 26862
rect 48318 26480 48374 26489
rect 48228 26444 48280 26450
rect 48318 26415 48374 26424
rect 48228 26386 48280 26392
rect 48332 26382 48360 26415
rect 48320 26376 48372 26382
rect 48320 26318 48372 26324
rect 48136 24336 48188 24342
rect 48136 24278 48188 24284
rect 48136 23316 48188 23322
rect 48136 23258 48188 23264
rect 48148 23118 48176 23258
rect 48044 23112 48096 23118
rect 48042 23080 48044 23089
rect 48136 23112 48188 23118
rect 48096 23080 48098 23089
rect 48136 23054 48188 23060
rect 48042 23015 48098 23024
rect 48332 22778 48360 26318
rect 48424 25294 48452 26862
rect 48596 26444 48648 26450
rect 48596 26386 48648 26392
rect 48504 25356 48556 25362
rect 48504 25298 48556 25304
rect 48412 25288 48464 25294
rect 48412 25230 48464 25236
rect 48516 23322 48544 25298
rect 48608 25294 48636 26386
rect 48700 26314 48728 27367
rect 48688 26308 48740 26314
rect 48688 26250 48740 26256
rect 48596 25288 48648 25294
rect 48596 25230 48648 25236
rect 48792 24834 48820 29582
rect 48872 26308 48924 26314
rect 48872 26250 48924 26256
rect 48700 24806 48820 24834
rect 48700 23798 48728 24806
rect 48780 24744 48832 24750
rect 48780 24686 48832 24692
rect 48688 23792 48740 23798
rect 48688 23734 48740 23740
rect 48792 23730 48820 24686
rect 48780 23724 48832 23730
rect 48780 23666 48832 23672
rect 48688 23656 48740 23662
rect 48688 23598 48740 23604
rect 48504 23316 48556 23322
rect 48504 23258 48556 23264
rect 48412 23180 48464 23186
rect 48412 23122 48464 23128
rect 48320 22772 48372 22778
rect 48320 22714 48372 22720
rect 47952 20868 48004 20874
rect 47952 20810 48004 20816
rect 47768 19780 47820 19786
rect 47768 19722 47820 19728
rect 47780 11898 47808 19722
rect 47860 19440 47912 19446
rect 47860 19382 47912 19388
rect 47768 11892 47820 11898
rect 47768 11834 47820 11840
rect 47768 10600 47820 10606
rect 47768 10542 47820 10548
rect 47676 8628 47728 8634
rect 47676 8570 47728 8576
rect 47492 8492 47544 8498
rect 47492 8434 47544 8440
rect 47398 7848 47454 7857
rect 47398 7783 47454 7792
rect 46756 5704 46808 5710
rect 46756 5646 46808 5652
rect 46768 2582 46796 5646
rect 47032 4684 47084 4690
rect 47032 4626 47084 4632
rect 47584 4684 47636 4690
rect 47584 4626 47636 4632
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46756 2576 46808 2582
rect 46756 2518 46808 2524
rect 46664 944 46716 950
rect 46664 886 46716 892
rect 46860 800 46888 2926
rect 47044 800 47072 4626
rect 47308 3596 47360 3602
rect 47308 3538 47360 3544
rect 47320 2774 47348 3538
rect 47228 2746 47348 2774
rect 47228 800 47256 2746
rect 47400 2304 47452 2310
rect 47400 2246 47452 2252
rect 47412 800 47440 2246
rect 47596 800 47624 4626
rect 47780 2582 47808 10542
rect 47872 8022 47900 19382
rect 47964 19310 47992 20810
rect 48318 20360 48374 20369
rect 48318 20295 48374 20304
rect 48332 20058 48360 20295
rect 48320 20052 48372 20058
rect 48320 19994 48372 20000
rect 48318 19952 48374 19961
rect 48318 19887 48320 19896
rect 48372 19887 48374 19896
rect 48320 19858 48372 19864
rect 47952 19304 48004 19310
rect 47952 19246 48004 19252
rect 48424 17678 48452 23122
rect 48516 22982 48544 23258
rect 48700 23186 48728 23598
rect 48884 23474 48912 26250
rect 48884 23446 49004 23474
rect 48872 23316 48924 23322
rect 48872 23258 48924 23264
rect 48688 23180 48740 23186
rect 48688 23122 48740 23128
rect 48504 22976 48556 22982
rect 48504 22918 48556 22924
rect 48780 22976 48832 22982
rect 48780 22918 48832 22924
rect 48504 22772 48556 22778
rect 48504 22714 48556 22720
rect 48412 17672 48464 17678
rect 48412 17614 48464 17620
rect 48136 17264 48188 17270
rect 48136 17206 48188 17212
rect 47952 15360 48004 15366
rect 47952 15302 48004 15308
rect 48044 15360 48096 15366
rect 48044 15302 48096 15308
rect 47860 8016 47912 8022
rect 47860 7958 47912 7964
rect 47964 4282 47992 15302
rect 48056 14958 48084 15302
rect 48044 14952 48096 14958
rect 48044 14894 48096 14900
rect 48044 12232 48096 12238
rect 48042 12200 48044 12209
rect 48096 12200 48098 12209
rect 48042 12135 48098 12144
rect 47952 4276 48004 4282
rect 47952 4218 48004 4224
rect 47952 3596 48004 3602
rect 47952 3538 48004 3544
rect 47964 2774 47992 3538
rect 48148 2990 48176 17206
rect 48320 13796 48372 13802
rect 48320 13738 48372 13744
rect 48228 13524 48280 13530
rect 48228 13466 48280 13472
rect 48240 12782 48268 13466
rect 48228 12776 48280 12782
rect 48228 12718 48280 12724
rect 48228 4072 48280 4078
rect 48228 4014 48280 4020
rect 48136 2984 48188 2990
rect 48136 2926 48188 2932
rect 48044 2848 48096 2854
rect 48044 2790 48096 2796
rect 47872 2746 47992 2774
rect 47768 2576 47820 2582
rect 47768 2518 47820 2524
rect 47676 2508 47728 2514
rect 47676 2450 47728 2456
rect 47688 1970 47716 2450
rect 47676 1964 47728 1970
rect 47676 1906 47728 1912
rect 47872 800 47900 2746
rect 48056 800 48084 2790
rect 48240 800 48268 4014
rect 48332 2650 48360 13738
rect 48516 12434 48544 22714
rect 48792 22438 48820 22918
rect 48780 22432 48832 22438
rect 48780 22374 48832 22380
rect 48688 21344 48740 21350
rect 48688 21286 48740 21292
rect 48596 20052 48648 20058
rect 48596 19994 48648 20000
rect 48608 19378 48636 19994
rect 48596 19372 48648 19378
rect 48596 19314 48648 19320
rect 48700 18601 48728 21286
rect 48780 19916 48832 19922
rect 48780 19858 48832 19864
rect 48686 18592 48742 18601
rect 48686 18527 48742 18536
rect 48792 17610 48820 19858
rect 48780 17604 48832 17610
rect 48780 17546 48832 17552
rect 48884 16250 48912 23258
rect 48872 16244 48924 16250
rect 48872 16186 48924 16192
rect 48778 15600 48834 15609
rect 48778 15535 48780 15544
rect 48832 15535 48834 15544
rect 48780 15506 48832 15512
rect 48976 12434 49004 23446
rect 49160 23186 49188 30534
rect 49528 30138 49556 33322
rect 49712 33266 49740 33612
rect 49252 30110 49556 30138
rect 49620 33238 49740 33266
rect 49252 27305 49280 30110
rect 49332 30048 49384 30054
rect 49332 29990 49384 29996
rect 49238 27296 49294 27305
rect 49238 27231 49294 27240
rect 49252 26926 49280 27231
rect 49240 26920 49292 26926
rect 49240 26862 49292 26868
rect 49344 24562 49372 29990
rect 49422 28656 49478 28665
rect 49422 28591 49478 28600
rect 49436 28558 49464 28591
rect 49424 28552 49476 28558
rect 49424 28494 49476 28500
rect 49516 28484 49568 28490
rect 49516 28426 49568 28432
rect 49528 28218 49556 28426
rect 49516 28212 49568 28218
rect 49516 28154 49568 28160
rect 49516 25288 49568 25294
rect 49516 25230 49568 25236
rect 49344 24534 49464 24562
rect 49056 23180 49108 23186
rect 49056 23122 49108 23128
rect 49148 23180 49200 23186
rect 49148 23122 49200 23128
rect 49068 14414 49096 23122
rect 49332 23044 49384 23050
rect 49332 22986 49384 22992
rect 49240 21412 49292 21418
rect 49240 21354 49292 21360
rect 49148 17808 49200 17814
rect 49148 17750 49200 17756
rect 49160 17610 49188 17750
rect 49148 17604 49200 17610
rect 49148 17546 49200 17552
rect 49148 16584 49200 16590
rect 49148 16526 49200 16532
rect 49056 14408 49108 14414
rect 49056 14350 49108 14356
rect 49160 12434 49188 16526
rect 49252 13258 49280 21354
rect 49344 17066 49372 22986
rect 49332 17060 49384 17066
rect 49332 17002 49384 17008
rect 49436 15366 49464 24534
rect 49528 23322 49556 25230
rect 49516 23316 49568 23322
rect 49516 23258 49568 23264
rect 49620 22094 49648 33238
rect 49700 32904 49752 32910
rect 49700 32846 49752 32852
rect 49712 31414 49740 32846
rect 49700 31408 49752 31414
rect 49700 31350 49752 31356
rect 49792 28552 49844 28558
rect 49792 28494 49844 28500
rect 49700 28212 49752 28218
rect 49700 28154 49752 28160
rect 49528 22066 49648 22094
rect 49528 16017 49556 22066
rect 49514 16008 49570 16017
rect 49514 15943 49570 15952
rect 49424 15360 49476 15366
rect 49424 15302 49476 15308
rect 49528 15178 49556 15943
rect 49608 15564 49660 15570
rect 49608 15506 49660 15512
rect 49436 15150 49556 15178
rect 49332 13796 49384 13802
rect 49332 13738 49384 13744
rect 49240 13252 49292 13258
rect 49240 13194 49292 13200
rect 48516 12406 48636 12434
rect 48412 9036 48464 9042
rect 48412 8978 48464 8984
rect 48424 6390 48452 8978
rect 48504 8356 48556 8362
rect 48504 8298 48556 8304
rect 48412 6384 48464 6390
rect 48412 6326 48464 6332
rect 48516 4214 48544 8298
rect 48608 6866 48636 12406
rect 48792 12406 49004 12434
rect 49068 12406 49188 12434
rect 48596 6860 48648 6866
rect 48596 6802 48648 6808
rect 48504 4208 48556 4214
rect 48504 4150 48556 4156
rect 48688 3664 48740 3670
rect 48688 3606 48740 3612
rect 48412 3528 48464 3534
rect 48412 3470 48464 3476
rect 48320 2644 48372 2650
rect 48320 2586 48372 2592
rect 48424 800 48452 3470
rect 48700 2106 48728 3606
rect 48688 2100 48740 2106
rect 48688 2042 48740 2048
rect 48688 1420 48740 1426
rect 48688 1362 48740 1368
rect 48700 800 48728 1362
rect 44916 604 44968 610
rect 44916 546 44968 552
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48792 134 48820 12406
rect 49068 12102 49096 12406
rect 49056 12096 49108 12102
rect 49056 12038 49108 12044
rect 49068 7342 49096 12038
rect 49344 9382 49372 13738
rect 49436 10742 49464 15150
rect 49516 13864 49568 13870
rect 49516 13806 49568 13812
rect 49424 10736 49476 10742
rect 49424 10678 49476 10684
rect 49332 9376 49384 9382
rect 49332 9318 49384 9324
rect 49240 8424 49292 8430
rect 49240 8366 49292 8372
rect 49148 8084 49200 8090
rect 49148 8026 49200 8032
rect 49056 7336 49108 7342
rect 49056 7278 49108 7284
rect 48872 7268 48924 7274
rect 48872 7210 48924 7216
rect 48884 7177 48912 7210
rect 48964 7200 49016 7206
rect 48870 7168 48926 7177
rect 48964 7142 49016 7148
rect 48870 7103 48926 7112
rect 48872 4072 48924 4078
rect 48872 4014 48924 4020
rect 48884 800 48912 4014
rect 48976 1358 49004 7142
rect 49056 3052 49108 3058
rect 49056 2994 49108 3000
rect 48964 1352 49016 1358
rect 48964 1294 49016 1300
rect 49068 800 49096 2994
rect 49160 2990 49188 8026
rect 49252 4690 49280 8366
rect 49332 8356 49384 8362
rect 49332 8298 49384 8304
rect 49344 6934 49372 8298
rect 49424 7336 49476 7342
rect 49424 7278 49476 7284
rect 49332 6928 49384 6934
rect 49332 6870 49384 6876
rect 49240 4684 49292 4690
rect 49240 4626 49292 4632
rect 49148 2984 49200 2990
rect 49148 2926 49200 2932
rect 49240 2916 49292 2922
rect 49240 2858 49292 2864
rect 49252 800 49280 2858
rect 49436 2836 49464 7278
rect 49528 4622 49556 13806
rect 49620 13802 49648 15506
rect 49608 13796 49660 13802
rect 49608 13738 49660 13744
rect 49712 12434 49740 28154
rect 49804 28150 49832 28494
rect 49792 28144 49844 28150
rect 49792 28086 49844 28092
rect 49896 26926 49924 34983
rect 49976 28144 50028 28150
rect 49974 28112 49976 28121
rect 50028 28112 50030 28121
rect 49974 28047 50030 28056
rect 49884 26920 49936 26926
rect 49884 26862 49936 26868
rect 49896 26450 49924 26862
rect 50080 26518 50108 38898
rect 50356 37890 50384 39200
rect 50712 38004 50764 38010
rect 50712 37946 50764 37952
rect 50172 37862 50384 37890
rect 50172 37398 50200 37862
rect 50300 37564 50596 37584
rect 50356 37562 50380 37564
rect 50436 37562 50460 37564
rect 50516 37562 50540 37564
rect 50378 37510 50380 37562
rect 50442 37510 50454 37562
rect 50516 37510 50518 37562
rect 50356 37508 50380 37510
rect 50436 37508 50460 37510
rect 50516 37508 50540 37510
rect 50300 37488 50596 37508
rect 50724 37466 50752 37946
rect 51276 37466 51304 39200
rect 52104 37466 52132 39200
rect 52368 37664 52420 37670
rect 52368 37606 52420 37612
rect 50712 37460 50764 37466
rect 50712 37402 50764 37408
rect 51264 37460 51316 37466
rect 51264 37402 51316 37408
rect 52092 37460 52144 37466
rect 52092 37402 52144 37408
rect 50160 37392 50212 37398
rect 50160 37334 50212 37340
rect 52380 37330 52408 37606
rect 53024 37398 53052 39200
rect 53852 37398 53880 39200
rect 54300 38548 54352 38554
rect 54300 38490 54352 38496
rect 53012 37392 53064 37398
rect 53012 37334 53064 37340
rect 53840 37392 53892 37398
rect 53840 37334 53892 37340
rect 51172 37324 51224 37330
rect 51172 37266 51224 37272
rect 52368 37324 52420 37330
rect 52368 37266 52420 37272
rect 53472 37324 53524 37330
rect 53472 37266 53524 37272
rect 50712 37120 50764 37126
rect 50712 37062 50764 37068
rect 50300 36476 50596 36496
rect 50356 36474 50380 36476
rect 50436 36474 50460 36476
rect 50516 36474 50540 36476
rect 50378 36422 50380 36474
rect 50442 36422 50454 36474
rect 50516 36422 50518 36474
rect 50356 36420 50380 36422
rect 50436 36420 50460 36422
rect 50516 36420 50540 36422
rect 50300 36400 50596 36420
rect 50300 35388 50596 35408
rect 50356 35386 50380 35388
rect 50436 35386 50460 35388
rect 50516 35386 50540 35388
rect 50378 35334 50380 35386
rect 50442 35334 50454 35386
rect 50516 35334 50518 35386
rect 50356 35332 50380 35334
rect 50436 35332 50460 35334
rect 50516 35332 50540 35334
rect 50300 35312 50596 35332
rect 50300 34300 50596 34320
rect 50356 34298 50380 34300
rect 50436 34298 50460 34300
rect 50516 34298 50540 34300
rect 50378 34246 50380 34298
rect 50442 34246 50454 34298
rect 50516 34246 50518 34298
rect 50356 34244 50380 34246
rect 50436 34244 50460 34246
rect 50516 34244 50540 34246
rect 50300 34224 50596 34244
rect 50300 33212 50596 33232
rect 50356 33210 50380 33212
rect 50436 33210 50460 33212
rect 50516 33210 50540 33212
rect 50378 33158 50380 33210
rect 50442 33158 50454 33210
rect 50516 33158 50518 33210
rect 50356 33156 50380 33158
rect 50436 33156 50460 33158
rect 50516 33156 50540 33158
rect 50300 33136 50596 33156
rect 50620 32836 50672 32842
rect 50620 32778 50672 32784
rect 50632 32745 50660 32778
rect 50618 32736 50674 32745
rect 50618 32671 50674 32680
rect 50300 32124 50596 32144
rect 50356 32122 50380 32124
rect 50436 32122 50460 32124
rect 50516 32122 50540 32124
rect 50378 32070 50380 32122
rect 50442 32070 50454 32122
rect 50516 32070 50518 32122
rect 50356 32068 50380 32070
rect 50436 32068 50460 32070
rect 50516 32068 50540 32070
rect 50300 32048 50596 32068
rect 50724 31754 50752 37062
rect 51184 36174 51212 37266
rect 53484 36786 53512 37266
rect 53564 36916 53616 36922
rect 53564 36858 53616 36864
rect 53576 36786 53604 36858
rect 53472 36780 53524 36786
rect 53472 36722 53524 36728
rect 53564 36780 53616 36786
rect 53564 36722 53616 36728
rect 52104 36638 52408 36666
rect 52104 36582 52132 36638
rect 52092 36576 52144 36582
rect 52092 36518 52144 36524
rect 52184 36576 52236 36582
rect 52184 36518 52236 36524
rect 52196 36242 52224 36518
rect 52380 36242 52408 36638
rect 52920 36644 52972 36650
rect 52920 36586 52972 36592
rect 52184 36236 52236 36242
rect 52184 36178 52236 36184
rect 52368 36236 52420 36242
rect 52368 36178 52420 36184
rect 51172 36168 51224 36174
rect 51172 36110 51224 36116
rect 51080 35828 51132 35834
rect 51080 35770 51132 35776
rect 51172 35828 51224 35834
rect 51172 35770 51224 35776
rect 51092 35630 51120 35770
rect 51080 35624 51132 35630
rect 51080 35566 51132 35572
rect 50804 34672 50856 34678
rect 50804 34614 50856 34620
rect 50988 34672 51040 34678
rect 50988 34614 51040 34620
rect 50816 32042 50844 34614
rect 51000 34513 51028 34614
rect 51184 34513 51212 35770
rect 52196 35306 52224 36178
rect 52276 36168 52328 36174
rect 52276 36110 52328 36116
rect 52736 36168 52788 36174
rect 52736 36110 52788 36116
rect 52012 35278 52224 35306
rect 50986 34504 51042 34513
rect 50986 34439 51042 34448
rect 51170 34504 51226 34513
rect 51170 34439 51226 34448
rect 51172 34128 51224 34134
rect 50894 34096 50950 34105
rect 50894 34031 50896 34040
rect 50948 34031 50950 34040
rect 51000 34088 51172 34116
rect 50896 34002 50948 34008
rect 51000 33998 51028 34088
rect 51172 34070 51224 34076
rect 50988 33992 51040 33998
rect 50988 33934 51040 33940
rect 51080 33380 51132 33386
rect 51080 33322 51132 33328
rect 51092 33289 51120 33322
rect 51078 33280 51134 33289
rect 51078 33215 51134 33224
rect 51078 32736 51134 32745
rect 51078 32671 51134 32680
rect 51092 32230 51120 32671
rect 50988 32224 51040 32230
rect 50986 32192 50988 32201
rect 51080 32224 51132 32230
rect 51040 32192 51042 32201
rect 51080 32166 51132 32172
rect 50986 32127 51042 32136
rect 50816 32014 51028 32042
rect 50160 31748 50212 31754
rect 50724 31726 50844 31754
rect 50160 31690 50212 31696
rect 50172 26568 50200 31690
rect 50300 31036 50596 31056
rect 50356 31034 50380 31036
rect 50436 31034 50460 31036
rect 50516 31034 50540 31036
rect 50378 30982 50380 31034
rect 50442 30982 50454 31034
rect 50516 30982 50518 31034
rect 50356 30980 50380 30982
rect 50436 30980 50460 30982
rect 50516 30980 50540 30982
rect 50300 30960 50596 30980
rect 50300 29948 50596 29968
rect 50356 29946 50380 29948
rect 50436 29946 50460 29948
rect 50516 29946 50540 29948
rect 50378 29894 50380 29946
rect 50442 29894 50454 29946
rect 50516 29894 50518 29946
rect 50356 29892 50380 29894
rect 50436 29892 50460 29894
rect 50516 29892 50540 29894
rect 50300 29872 50596 29892
rect 50300 28860 50596 28880
rect 50356 28858 50380 28860
rect 50436 28858 50460 28860
rect 50516 28858 50540 28860
rect 50378 28806 50380 28858
rect 50442 28806 50454 28858
rect 50516 28806 50518 28858
rect 50356 28804 50380 28806
rect 50436 28804 50460 28806
rect 50516 28804 50540 28806
rect 50300 28784 50596 28804
rect 50300 27772 50596 27792
rect 50356 27770 50380 27772
rect 50436 27770 50460 27772
rect 50516 27770 50540 27772
rect 50378 27718 50380 27770
rect 50442 27718 50454 27770
rect 50516 27718 50518 27770
rect 50356 27716 50380 27718
rect 50436 27716 50460 27718
rect 50516 27716 50540 27718
rect 50300 27696 50596 27716
rect 50620 27600 50672 27606
rect 50712 27600 50764 27606
rect 50620 27542 50672 27548
rect 50710 27568 50712 27577
rect 50764 27568 50766 27577
rect 50300 26684 50596 26704
rect 50356 26682 50380 26684
rect 50436 26682 50460 26684
rect 50516 26682 50540 26684
rect 50378 26630 50380 26682
rect 50442 26630 50454 26682
rect 50516 26630 50518 26682
rect 50356 26628 50380 26630
rect 50436 26628 50460 26630
rect 50516 26628 50540 26630
rect 50300 26608 50596 26628
rect 50172 26540 50384 26568
rect 50068 26512 50120 26518
rect 50068 26454 50120 26460
rect 50356 26450 50384 26540
rect 49884 26444 49936 26450
rect 49884 26386 49936 26392
rect 50252 26444 50304 26450
rect 50252 26386 50304 26392
rect 50344 26444 50396 26450
rect 50344 26386 50396 26392
rect 50264 26330 50292 26386
rect 50632 26330 50660 27542
rect 50710 27503 50766 27512
rect 50712 27396 50764 27402
rect 50712 27338 50764 27344
rect 50724 27169 50752 27338
rect 50710 27160 50766 27169
rect 50710 27095 50766 27104
rect 50712 26920 50764 26926
rect 50712 26862 50764 26868
rect 49988 26302 50292 26330
rect 50540 26302 50660 26330
rect 49884 26240 49936 26246
rect 49884 26182 49936 26188
rect 49792 25764 49844 25770
rect 49792 25706 49844 25712
rect 49804 23050 49832 25706
rect 49792 23044 49844 23050
rect 49792 22986 49844 22992
rect 49896 22778 49924 26182
rect 49884 22772 49936 22778
rect 49884 22714 49936 22720
rect 49792 13524 49844 13530
rect 49792 13466 49844 13472
rect 49804 13258 49832 13466
rect 49792 13252 49844 13258
rect 49792 13194 49844 13200
rect 49712 12406 49832 12434
rect 49700 7744 49752 7750
rect 49700 7686 49752 7692
rect 49712 7478 49740 7686
rect 49608 7472 49660 7478
rect 49608 7414 49660 7420
rect 49700 7472 49752 7478
rect 49700 7414 49752 7420
rect 49620 7342 49648 7414
rect 49608 7336 49660 7342
rect 49608 7278 49660 7284
rect 49700 7200 49752 7206
rect 49700 7142 49752 7148
rect 49712 6934 49740 7142
rect 49700 6928 49752 6934
rect 49700 6870 49752 6876
rect 49516 4616 49568 4622
rect 49516 4558 49568 4564
rect 49516 4072 49568 4078
rect 49516 4014 49568 4020
rect 49344 2808 49464 2836
rect 48780 128 48832 134
rect 48780 70 48832 76
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49344 474 49372 2808
rect 49528 2774 49556 4014
rect 49712 3738 49740 6870
rect 49804 3777 49832 12406
rect 49884 9172 49936 9178
rect 49884 9114 49936 9120
rect 49790 3768 49846 3777
rect 49700 3732 49752 3738
rect 49790 3703 49846 3712
rect 49700 3674 49752 3680
rect 49608 3664 49660 3670
rect 49608 3606 49660 3612
rect 49620 2854 49648 3606
rect 49784 3596 49836 3602
rect 49712 3556 49784 3584
rect 49608 2848 49660 2854
rect 49608 2790 49660 2796
rect 49436 2746 49556 2774
rect 49436 800 49464 2746
rect 49712 800 49740 3556
rect 49784 3538 49836 3544
rect 49790 3496 49846 3505
rect 49790 3431 49846 3440
rect 49804 2990 49832 3431
rect 49792 2984 49844 2990
rect 49792 2926 49844 2932
rect 49792 2848 49844 2854
rect 49792 2790 49844 2796
rect 49804 2650 49832 2790
rect 49792 2644 49844 2650
rect 49792 2586 49844 2592
rect 49896 2514 49924 9114
rect 49988 8362 50016 26302
rect 50068 26240 50120 26246
rect 50068 26182 50120 26188
rect 50080 19378 50108 26182
rect 50436 25968 50488 25974
rect 50436 25910 50488 25916
rect 50448 25770 50476 25910
rect 50540 25786 50568 26302
rect 50436 25764 50488 25770
rect 50540 25758 50660 25786
rect 50436 25706 50488 25712
rect 50300 25596 50596 25616
rect 50356 25594 50380 25596
rect 50436 25594 50460 25596
rect 50516 25594 50540 25596
rect 50378 25542 50380 25594
rect 50442 25542 50454 25594
rect 50516 25542 50518 25594
rect 50356 25540 50380 25542
rect 50436 25540 50460 25542
rect 50516 25540 50540 25542
rect 50300 25520 50596 25540
rect 50436 25152 50488 25158
rect 50436 25094 50488 25100
rect 50448 24886 50476 25094
rect 50436 24880 50488 24886
rect 50436 24822 50488 24828
rect 50526 24848 50582 24857
rect 50526 24783 50528 24792
rect 50580 24783 50582 24792
rect 50528 24754 50580 24760
rect 50526 24712 50582 24721
rect 50526 24647 50528 24656
rect 50580 24647 50582 24656
rect 50528 24618 50580 24624
rect 50300 24508 50596 24528
rect 50356 24506 50380 24508
rect 50436 24506 50460 24508
rect 50516 24506 50540 24508
rect 50378 24454 50380 24506
rect 50442 24454 50454 24506
rect 50516 24454 50518 24506
rect 50356 24452 50380 24454
rect 50436 24452 50460 24454
rect 50516 24452 50540 24454
rect 50300 24432 50596 24452
rect 50344 23860 50396 23866
rect 50344 23802 50396 23808
rect 50356 23594 50384 23802
rect 50632 23798 50660 25758
rect 50620 23792 50672 23798
rect 50620 23734 50672 23740
rect 50344 23588 50396 23594
rect 50344 23530 50396 23536
rect 50300 23420 50596 23440
rect 50356 23418 50380 23420
rect 50436 23418 50460 23420
rect 50516 23418 50540 23420
rect 50378 23366 50380 23418
rect 50442 23366 50454 23418
rect 50516 23366 50518 23418
rect 50356 23364 50380 23366
rect 50436 23364 50460 23366
rect 50516 23364 50540 23366
rect 50300 23344 50596 23364
rect 50724 22438 50752 26862
rect 50712 22432 50764 22438
rect 50712 22374 50764 22380
rect 50300 22332 50596 22352
rect 50356 22330 50380 22332
rect 50436 22330 50460 22332
rect 50516 22330 50540 22332
rect 50378 22278 50380 22330
rect 50442 22278 50454 22330
rect 50516 22278 50518 22330
rect 50356 22276 50380 22278
rect 50436 22276 50460 22278
rect 50516 22276 50540 22278
rect 50300 22256 50596 22276
rect 50160 21412 50212 21418
rect 50160 21354 50212 21360
rect 50172 19718 50200 21354
rect 50620 21344 50672 21350
rect 50620 21286 50672 21292
rect 50300 21244 50596 21264
rect 50356 21242 50380 21244
rect 50436 21242 50460 21244
rect 50516 21242 50540 21244
rect 50378 21190 50380 21242
rect 50442 21190 50454 21242
rect 50516 21190 50518 21242
rect 50356 21188 50380 21190
rect 50436 21188 50460 21190
rect 50516 21188 50540 21190
rect 50300 21168 50596 21188
rect 50300 20156 50596 20176
rect 50356 20154 50380 20156
rect 50436 20154 50460 20156
rect 50516 20154 50540 20156
rect 50378 20102 50380 20154
rect 50442 20102 50454 20154
rect 50516 20102 50518 20154
rect 50356 20100 50380 20102
rect 50436 20100 50460 20102
rect 50516 20100 50540 20102
rect 50300 20080 50596 20100
rect 50160 19712 50212 19718
rect 50160 19654 50212 19660
rect 50068 19372 50120 19378
rect 50068 19314 50120 19320
rect 50172 19334 50200 19654
rect 50436 19508 50488 19514
rect 50436 19450 50488 19456
rect 50172 19310 50292 19334
rect 50448 19310 50476 19450
rect 50632 19310 50660 21286
rect 50816 20754 50844 31726
rect 50894 28656 50950 28665
rect 50894 28591 50950 28600
rect 50908 24970 50936 28591
rect 51000 28393 51028 32014
rect 51080 31952 51132 31958
rect 51080 31894 51132 31900
rect 51092 30734 51120 31894
rect 51816 31476 51868 31482
rect 51816 31418 51868 31424
rect 51908 31476 51960 31482
rect 51908 31418 51960 31424
rect 51080 30728 51132 30734
rect 51080 30670 51132 30676
rect 51828 30598 51856 31418
rect 51816 30592 51868 30598
rect 51816 30534 51868 30540
rect 50986 28384 51042 28393
rect 50986 28319 51042 28328
rect 51170 28384 51226 28393
rect 51170 28319 51226 28328
rect 51184 27946 51212 28319
rect 51080 27940 51132 27946
rect 51080 27882 51132 27888
rect 51172 27940 51224 27946
rect 51172 27882 51224 27888
rect 51092 27826 51120 27882
rect 51092 27798 51212 27826
rect 51078 27704 51134 27713
rect 51184 27674 51212 27798
rect 51078 27639 51080 27648
rect 51132 27639 51134 27648
rect 51172 27668 51224 27674
rect 51080 27610 51132 27616
rect 51172 27610 51224 27616
rect 51446 27160 51502 27169
rect 51446 27095 51502 27104
rect 50986 25664 51042 25673
rect 50986 25599 51042 25608
rect 51000 25362 51028 25599
rect 50988 25356 51040 25362
rect 50988 25298 51040 25304
rect 51262 25256 51318 25265
rect 51262 25191 51264 25200
rect 51316 25191 51318 25200
rect 51264 25162 51316 25168
rect 50908 24942 51028 24970
rect 51000 24750 51028 24942
rect 51354 24848 51410 24857
rect 51354 24783 51356 24792
rect 51408 24783 51410 24792
rect 51356 24754 51408 24760
rect 50988 24744 51040 24750
rect 50988 24686 51040 24692
rect 51172 24744 51224 24750
rect 51172 24686 51224 24692
rect 51184 23225 51212 24686
rect 51170 23216 51226 23225
rect 51170 23151 51226 23160
rect 50896 21684 50948 21690
rect 50896 21626 50948 21632
rect 51356 21684 51408 21690
rect 51356 21626 51408 21632
rect 50908 21593 50936 21626
rect 50894 21584 50950 21593
rect 50894 21519 50950 21528
rect 51368 21146 51396 21626
rect 51356 21140 51408 21146
rect 51356 21082 51408 21088
rect 51080 21004 51132 21010
rect 51080 20946 51132 20952
rect 51172 21004 51224 21010
rect 51172 20946 51224 20952
rect 50894 20904 50950 20913
rect 51092 20874 51120 20946
rect 51184 20913 51212 20946
rect 51170 20904 51226 20913
rect 50894 20839 50896 20848
rect 50948 20839 50950 20848
rect 51080 20868 51132 20874
rect 50896 20810 50948 20816
rect 51170 20839 51226 20848
rect 51080 20810 51132 20816
rect 50816 20726 50936 20754
rect 50172 19306 50304 19310
rect 50252 19304 50304 19306
rect 50252 19246 50304 19252
rect 50436 19304 50488 19310
rect 50436 19246 50488 19252
rect 50620 19304 50672 19310
rect 50620 19246 50672 19252
rect 50804 19304 50856 19310
rect 50804 19246 50856 19252
rect 50300 19068 50596 19088
rect 50356 19066 50380 19068
rect 50436 19066 50460 19068
rect 50516 19066 50540 19068
rect 50378 19014 50380 19066
rect 50442 19014 50454 19066
rect 50516 19014 50518 19066
rect 50356 19012 50380 19014
rect 50436 19012 50460 19014
rect 50516 19012 50540 19014
rect 50300 18992 50596 19012
rect 50632 18358 50660 19246
rect 50816 19174 50844 19246
rect 50804 19168 50856 19174
rect 50804 19110 50856 19116
rect 50710 18864 50766 18873
rect 50710 18799 50766 18808
rect 50804 18828 50856 18834
rect 50724 18426 50752 18799
rect 50804 18770 50856 18776
rect 50816 18737 50844 18770
rect 50802 18728 50858 18737
rect 50802 18663 50858 18672
rect 50712 18420 50764 18426
rect 50712 18362 50764 18368
rect 50620 18352 50672 18358
rect 50620 18294 50672 18300
rect 50300 17980 50596 18000
rect 50356 17978 50380 17980
rect 50436 17978 50460 17980
rect 50516 17978 50540 17980
rect 50378 17926 50380 17978
rect 50442 17926 50454 17978
rect 50516 17926 50518 17978
rect 50356 17924 50380 17926
rect 50436 17924 50460 17926
rect 50516 17924 50540 17926
rect 50300 17904 50596 17924
rect 50712 17196 50764 17202
rect 50712 17138 50764 17144
rect 50300 16892 50596 16912
rect 50356 16890 50380 16892
rect 50436 16890 50460 16892
rect 50516 16890 50540 16892
rect 50378 16838 50380 16890
rect 50442 16838 50454 16890
rect 50516 16838 50518 16890
rect 50356 16836 50380 16838
rect 50436 16836 50460 16838
rect 50516 16836 50540 16838
rect 50300 16816 50596 16836
rect 50300 15804 50596 15824
rect 50356 15802 50380 15804
rect 50436 15802 50460 15804
rect 50516 15802 50540 15804
rect 50378 15750 50380 15802
rect 50442 15750 50454 15802
rect 50516 15750 50518 15802
rect 50356 15748 50380 15750
rect 50436 15748 50460 15750
rect 50516 15748 50540 15750
rect 50300 15728 50596 15748
rect 50160 15360 50212 15366
rect 50160 15302 50212 15308
rect 50068 12232 50120 12238
rect 50068 12174 50120 12180
rect 50080 12102 50108 12174
rect 50068 12096 50120 12102
rect 50068 12038 50120 12044
rect 49976 8356 50028 8362
rect 49976 8298 50028 8304
rect 50080 7342 50108 12038
rect 50172 7750 50200 15302
rect 50300 14716 50596 14736
rect 50356 14714 50380 14716
rect 50436 14714 50460 14716
rect 50516 14714 50540 14716
rect 50378 14662 50380 14714
rect 50442 14662 50454 14714
rect 50516 14662 50518 14714
rect 50356 14660 50380 14662
rect 50436 14660 50460 14662
rect 50516 14660 50540 14662
rect 50300 14640 50596 14660
rect 50300 13628 50596 13648
rect 50356 13626 50380 13628
rect 50436 13626 50460 13628
rect 50516 13626 50540 13628
rect 50378 13574 50380 13626
rect 50442 13574 50454 13626
rect 50516 13574 50518 13626
rect 50356 13572 50380 13574
rect 50436 13572 50460 13574
rect 50516 13572 50540 13574
rect 50300 13552 50596 13572
rect 50300 12540 50596 12560
rect 50356 12538 50380 12540
rect 50436 12538 50460 12540
rect 50516 12538 50540 12540
rect 50378 12486 50380 12538
rect 50442 12486 50454 12538
rect 50516 12486 50518 12538
rect 50356 12484 50380 12486
rect 50436 12484 50460 12486
rect 50516 12484 50540 12486
rect 50300 12464 50596 12484
rect 50724 12102 50752 17138
rect 50804 14000 50856 14006
rect 50804 13942 50856 13948
rect 50712 12096 50764 12102
rect 50712 12038 50764 12044
rect 50300 11452 50596 11472
rect 50356 11450 50380 11452
rect 50436 11450 50460 11452
rect 50516 11450 50540 11452
rect 50378 11398 50380 11450
rect 50442 11398 50454 11450
rect 50516 11398 50518 11450
rect 50356 11396 50380 11398
rect 50436 11396 50460 11398
rect 50516 11396 50540 11398
rect 50300 11376 50596 11396
rect 50816 10962 50844 13942
rect 50632 10934 50844 10962
rect 50632 10470 50660 10934
rect 50620 10464 50672 10470
rect 50620 10406 50672 10412
rect 50300 10364 50596 10384
rect 50356 10362 50380 10364
rect 50436 10362 50460 10364
rect 50516 10362 50540 10364
rect 50378 10310 50380 10362
rect 50442 10310 50454 10362
rect 50516 10310 50518 10362
rect 50356 10308 50380 10310
rect 50436 10308 50460 10310
rect 50516 10308 50540 10310
rect 50300 10288 50596 10308
rect 50300 9276 50596 9296
rect 50356 9274 50380 9276
rect 50436 9274 50460 9276
rect 50516 9274 50540 9276
rect 50378 9222 50380 9274
rect 50442 9222 50454 9274
rect 50516 9222 50518 9274
rect 50356 9220 50380 9222
rect 50436 9220 50460 9222
rect 50516 9220 50540 9222
rect 50300 9200 50596 9220
rect 50632 8650 50660 10406
rect 50712 10260 50764 10266
rect 50712 10202 50764 10208
rect 50540 8622 50660 8650
rect 50540 8498 50568 8622
rect 50528 8492 50580 8498
rect 50528 8434 50580 8440
rect 50436 8424 50488 8430
rect 50724 8378 50752 10202
rect 50908 9674 50936 20726
rect 51264 19236 51316 19242
rect 51264 19178 51316 19184
rect 51080 19168 51132 19174
rect 51080 19110 51132 19116
rect 51172 19168 51224 19174
rect 51172 19110 51224 19116
rect 51092 15366 51120 19110
rect 51184 18873 51212 19110
rect 51170 18864 51226 18873
rect 51170 18799 51226 18808
rect 51276 18358 51304 19178
rect 51264 18352 51316 18358
rect 51264 18294 51316 18300
rect 51356 17128 51408 17134
rect 51356 17070 51408 17076
rect 51080 15360 51132 15366
rect 51080 15302 51132 15308
rect 51172 15088 51224 15094
rect 51172 15030 51224 15036
rect 51264 15088 51316 15094
rect 51264 15030 51316 15036
rect 51080 15020 51132 15026
rect 51080 14962 51132 14968
rect 51092 14929 51120 14962
rect 51184 14958 51212 15030
rect 51172 14952 51224 14958
rect 51078 14920 51134 14929
rect 51172 14894 51224 14900
rect 51078 14855 51134 14864
rect 51276 14634 51304 15030
rect 51092 14606 51304 14634
rect 51092 14550 51120 14606
rect 51080 14544 51132 14550
rect 51080 14486 51132 14492
rect 51264 14476 51316 14482
rect 51264 14418 51316 14424
rect 51276 14278 51304 14418
rect 51264 14272 51316 14278
rect 51264 14214 51316 14220
rect 50988 9920 51040 9926
rect 50988 9862 51040 9868
rect 50816 9646 50936 9674
rect 51000 9674 51028 9862
rect 51000 9646 51212 9674
rect 50816 9178 50844 9646
rect 51080 9512 51132 9518
rect 51080 9454 51132 9460
rect 51092 9178 51120 9454
rect 50804 9172 50856 9178
rect 50804 9114 50856 9120
rect 51080 9172 51132 9178
rect 51080 9114 51132 9120
rect 50804 8560 50856 8566
rect 50802 8528 50804 8537
rect 50856 8528 50858 8537
rect 50802 8463 50858 8472
rect 51078 8528 51134 8537
rect 51078 8463 51080 8472
rect 51132 8463 51134 8472
rect 51080 8434 51132 8440
rect 50488 8372 50752 8378
rect 50436 8366 50752 8372
rect 50448 8350 50752 8366
rect 51184 8362 51212 9646
rect 50804 8356 50856 8362
rect 50804 8298 50856 8304
rect 51172 8356 51224 8362
rect 51172 8298 51224 8304
rect 50300 8188 50596 8208
rect 50356 8186 50380 8188
rect 50436 8186 50460 8188
rect 50516 8186 50540 8188
rect 50378 8134 50380 8186
rect 50442 8134 50454 8186
rect 50516 8134 50518 8186
rect 50356 8132 50380 8134
rect 50436 8132 50460 8134
rect 50516 8132 50540 8134
rect 50300 8112 50596 8132
rect 50160 7744 50212 7750
rect 50160 7686 50212 7692
rect 50712 7744 50764 7750
rect 50712 7686 50764 7692
rect 50068 7336 50120 7342
rect 50068 7278 50120 7284
rect 50160 7200 50212 7206
rect 50158 7168 50160 7177
rect 50212 7168 50214 7177
rect 50158 7103 50214 7112
rect 50300 7100 50596 7120
rect 50356 7098 50380 7100
rect 50436 7098 50460 7100
rect 50516 7098 50540 7100
rect 50378 7046 50380 7098
rect 50442 7046 50454 7098
rect 50516 7046 50518 7098
rect 50356 7044 50380 7046
rect 50436 7044 50460 7046
rect 50516 7044 50540 7046
rect 50300 7024 50596 7044
rect 50724 6866 50752 7686
rect 50712 6860 50764 6866
rect 50712 6802 50764 6808
rect 49976 6792 50028 6798
rect 49976 6734 50028 6740
rect 49988 2854 50016 6734
rect 50816 6662 50844 8298
rect 50804 6656 50856 6662
rect 50804 6598 50856 6604
rect 50300 6012 50596 6032
rect 50356 6010 50380 6012
rect 50436 6010 50460 6012
rect 50516 6010 50540 6012
rect 50378 5958 50380 6010
rect 50442 5958 50454 6010
rect 50516 5958 50518 6010
rect 50356 5956 50380 5958
rect 50436 5956 50460 5958
rect 50516 5956 50540 5958
rect 50300 5936 50596 5956
rect 50300 4924 50596 4944
rect 50356 4922 50380 4924
rect 50436 4922 50460 4924
rect 50516 4922 50540 4924
rect 50378 4870 50380 4922
rect 50442 4870 50454 4922
rect 50516 4870 50518 4922
rect 50356 4868 50380 4870
rect 50436 4868 50460 4870
rect 50516 4868 50540 4870
rect 50300 4848 50596 4868
rect 50988 4752 51040 4758
rect 50988 4694 51040 4700
rect 50160 4072 50212 4078
rect 50160 4014 50212 4020
rect 50804 4072 50856 4078
rect 50804 4014 50856 4020
rect 50172 3482 50200 4014
rect 50300 3836 50596 3856
rect 50356 3834 50380 3836
rect 50436 3834 50460 3836
rect 50516 3834 50540 3836
rect 50378 3782 50380 3834
rect 50442 3782 50454 3834
rect 50516 3782 50518 3834
rect 50356 3780 50380 3782
rect 50436 3780 50460 3782
rect 50516 3780 50540 3782
rect 50300 3760 50596 3780
rect 50816 3482 50844 4014
rect 50896 3596 50948 3602
rect 50896 3538 50948 3544
rect 50080 3454 50200 3482
rect 50724 3454 50844 3482
rect 49976 2848 50028 2854
rect 49976 2790 50028 2796
rect 49976 2644 50028 2650
rect 49976 2586 50028 2592
rect 49884 2508 49936 2514
rect 49884 2450 49936 2456
rect 49988 1306 50016 2586
rect 49896 1278 50016 1306
rect 49896 800 49924 1278
rect 50080 800 50108 3454
rect 50160 2916 50212 2922
rect 50160 2858 50212 2864
rect 50172 1442 50200 2858
rect 50300 2748 50596 2768
rect 50356 2746 50380 2748
rect 50436 2746 50460 2748
rect 50516 2746 50540 2748
rect 50378 2694 50380 2746
rect 50442 2694 50454 2746
rect 50516 2694 50518 2746
rect 50356 2692 50380 2694
rect 50436 2692 50460 2694
rect 50516 2692 50540 2694
rect 50300 2672 50596 2692
rect 50528 2440 50580 2446
rect 50528 2382 50580 2388
rect 50436 2372 50488 2378
rect 50436 2314 50488 2320
rect 50172 1414 50292 1442
rect 50264 800 50292 1414
rect 50448 800 50476 2314
rect 50540 1426 50568 2382
rect 50528 1420 50580 1426
rect 50528 1362 50580 1368
rect 50724 800 50752 3454
rect 50804 3052 50856 3058
rect 50804 2994 50856 3000
rect 49332 468 49384 474
rect 49332 410 49384 416
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50816 610 50844 2994
rect 50908 800 50936 3538
rect 51000 3058 51028 4694
rect 51264 4004 51316 4010
rect 51264 3946 51316 3952
rect 50988 3052 51040 3058
rect 50988 2994 51040 3000
rect 51080 2848 51132 2854
rect 51080 2790 51132 2796
rect 51092 800 51120 2790
rect 51276 800 51304 3946
rect 51368 2922 51396 17070
rect 51460 6390 51488 27095
rect 51816 25356 51868 25362
rect 51816 25298 51868 25304
rect 51540 24744 51592 24750
rect 51538 24712 51540 24721
rect 51592 24712 51594 24721
rect 51538 24647 51594 24656
rect 51724 22024 51776 22030
rect 51724 21966 51776 21972
rect 51736 21894 51764 21966
rect 51724 21888 51776 21894
rect 51724 21830 51776 21836
rect 51722 18864 51778 18873
rect 51722 18799 51778 18808
rect 51736 18630 51764 18799
rect 51724 18624 51776 18630
rect 51724 18566 51776 18572
rect 51724 10736 51776 10742
rect 51724 10678 51776 10684
rect 51736 10606 51764 10678
rect 51724 10600 51776 10606
rect 51724 10542 51776 10548
rect 51540 9512 51592 9518
rect 51828 9489 51856 25298
rect 51920 25294 51948 31418
rect 51908 25288 51960 25294
rect 51908 25230 51960 25236
rect 51908 20596 51960 20602
rect 51908 20538 51960 20544
rect 51920 20398 51948 20538
rect 51908 20392 51960 20398
rect 51908 20334 51960 20340
rect 51908 10600 51960 10606
rect 51908 10542 51960 10548
rect 51540 9454 51592 9460
rect 51814 9480 51870 9489
rect 51552 8566 51580 9454
rect 51814 9415 51870 9424
rect 51816 8832 51868 8838
rect 51814 8800 51816 8809
rect 51868 8800 51870 8809
rect 51814 8735 51870 8744
rect 51540 8560 51592 8566
rect 51540 8502 51592 8508
rect 51448 6384 51500 6390
rect 51448 6326 51500 6332
rect 51356 2916 51408 2922
rect 51356 2858 51408 2864
rect 51448 2916 51500 2922
rect 51448 2858 51500 2864
rect 51460 800 51488 2858
rect 51552 2582 51580 8502
rect 51920 6118 51948 10542
rect 52012 6186 52040 35278
rect 52288 35222 52316 36110
rect 52184 35216 52236 35222
rect 52182 35184 52184 35193
rect 52276 35216 52328 35222
rect 52236 35184 52238 35193
rect 52276 35158 52328 35164
rect 52182 35119 52238 35128
rect 52368 35148 52420 35154
rect 52368 35090 52420 35096
rect 52380 34406 52408 35090
rect 52276 34400 52328 34406
rect 52276 34342 52328 34348
rect 52368 34400 52420 34406
rect 52368 34342 52420 34348
rect 52288 33998 52316 34342
rect 52276 33992 52328 33998
rect 52276 33934 52328 33940
rect 52368 32224 52420 32230
rect 52368 32166 52420 32172
rect 52380 31754 52408 32166
rect 52288 31726 52408 31754
rect 52182 31648 52238 31657
rect 52182 31583 52238 31592
rect 52090 25528 52146 25537
rect 52090 25463 52092 25472
rect 52144 25463 52146 25472
rect 52092 25434 52144 25440
rect 52196 25362 52224 31583
rect 52288 30161 52316 31726
rect 52644 31408 52696 31414
rect 52644 31350 52696 31356
rect 52274 30152 52330 30161
rect 52274 30087 52330 30096
rect 52184 25356 52236 25362
rect 52184 25298 52236 25304
rect 52196 22094 52224 25298
rect 52104 22066 52224 22094
rect 52000 6180 52052 6186
rect 52000 6122 52052 6128
rect 51908 6112 51960 6118
rect 51908 6054 51960 6060
rect 52000 5228 52052 5234
rect 52000 5170 52052 5176
rect 52012 5030 52040 5170
rect 52000 5024 52052 5030
rect 52000 4966 52052 4972
rect 52104 4554 52132 22066
rect 52288 21554 52316 30087
rect 52366 29608 52422 29617
rect 52366 29543 52422 29552
rect 52380 28762 52408 29543
rect 52368 28756 52420 28762
rect 52368 28698 52420 28704
rect 52460 28552 52512 28558
rect 52460 28494 52512 28500
rect 52368 27328 52420 27334
rect 52368 27270 52420 27276
rect 52380 25770 52408 27270
rect 52368 25764 52420 25770
rect 52368 25706 52420 25712
rect 52380 22166 52408 25706
rect 52472 24614 52500 28494
rect 52656 26926 52684 31350
rect 52552 26920 52604 26926
rect 52550 26888 52552 26897
rect 52644 26920 52696 26926
rect 52604 26888 52606 26897
rect 52644 26862 52696 26868
rect 52550 26823 52606 26832
rect 52550 26480 52606 26489
rect 52550 26415 52552 26424
rect 52604 26415 52606 26424
rect 52552 26386 52604 26392
rect 52460 24608 52512 24614
rect 52460 24550 52512 24556
rect 52368 22160 52420 22166
rect 52368 22102 52420 22108
rect 52276 21548 52328 21554
rect 52276 21490 52328 21496
rect 52184 21480 52236 21486
rect 52184 21422 52236 21428
rect 52196 5234 52224 21422
rect 52288 21350 52316 21490
rect 52276 21344 52328 21350
rect 52276 21286 52328 21292
rect 52276 20460 52328 20466
rect 52276 20402 52328 20408
rect 52288 20330 52316 20402
rect 52472 20330 52500 24550
rect 52644 22092 52696 22098
rect 52748 22094 52776 36110
rect 52828 31816 52880 31822
rect 52828 31758 52880 31764
rect 52840 31414 52868 31758
rect 52828 31408 52880 31414
rect 52828 31350 52880 31356
rect 52828 27600 52880 27606
rect 52828 27542 52880 27548
rect 52840 26858 52868 27542
rect 52828 26852 52880 26858
rect 52828 26794 52880 26800
rect 52828 26240 52880 26246
rect 52828 26182 52880 26188
rect 52840 25838 52868 26182
rect 52828 25832 52880 25838
rect 52828 25774 52880 25780
rect 52828 25152 52880 25158
rect 52828 25094 52880 25100
rect 52840 24954 52868 25094
rect 52828 24948 52880 24954
rect 52828 24890 52880 24896
rect 52748 22066 52868 22094
rect 52644 22034 52696 22040
rect 52552 21548 52604 21554
rect 52552 21490 52604 21496
rect 52276 20324 52328 20330
rect 52276 20266 52328 20272
rect 52460 20324 52512 20330
rect 52460 20266 52512 20272
rect 52288 19514 52316 20266
rect 52276 19508 52328 19514
rect 52276 19450 52328 19456
rect 52276 18624 52328 18630
rect 52274 18592 52276 18601
rect 52328 18592 52330 18601
rect 52274 18527 52330 18536
rect 52460 15156 52512 15162
rect 52460 15098 52512 15104
rect 52472 14346 52500 15098
rect 52564 14550 52592 21490
rect 52656 19446 52684 22034
rect 52736 21344 52788 21350
rect 52736 21286 52788 21292
rect 52644 19440 52696 19446
rect 52644 19382 52696 19388
rect 52642 19272 52698 19281
rect 52642 19207 52644 19216
rect 52696 19207 52698 19216
rect 52644 19178 52696 19184
rect 52552 14544 52604 14550
rect 52552 14486 52604 14492
rect 52460 14340 52512 14346
rect 52460 14282 52512 14288
rect 52748 10062 52776 21286
rect 52840 16726 52868 22066
rect 52828 16720 52880 16726
rect 52828 16662 52880 16668
rect 52840 12986 52868 16662
rect 52828 12980 52880 12986
rect 52828 12922 52880 12928
rect 52736 10056 52788 10062
rect 52736 9998 52788 10004
rect 52368 8832 52420 8838
rect 52368 8774 52420 8780
rect 52380 6361 52408 8774
rect 52366 6352 52422 6361
rect 52366 6287 52422 6296
rect 52734 6352 52790 6361
rect 52734 6287 52790 6296
rect 52748 6254 52776 6287
rect 52736 6248 52788 6254
rect 52736 6190 52788 6196
rect 52828 5568 52880 5574
rect 52828 5510 52880 5516
rect 52184 5228 52236 5234
rect 52184 5170 52236 5176
rect 52368 4684 52420 4690
rect 52368 4626 52420 4632
rect 52552 4684 52604 4690
rect 52552 4626 52604 4632
rect 52092 4548 52144 4554
rect 52092 4490 52144 4496
rect 52092 3596 52144 3602
rect 52092 3538 52144 3544
rect 51540 2576 51592 2582
rect 51540 2518 51592 2524
rect 51632 2508 51684 2514
rect 51632 2450 51684 2456
rect 51644 2106 51672 2450
rect 51724 2304 51776 2310
rect 51724 2246 51776 2252
rect 51632 2100 51684 2106
rect 51632 2042 51684 2048
rect 51736 800 51764 2246
rect 51908 1896 51960 1902
rect 51908 1838 51960 1844
rect 51920 800 51948 1838
rect 52104 800 52132 3538
rect 52380 2582 52408 4626
rect 52368 2576 52420 2582
rect 52368 2518 52420 2524
rect 52460 2508 52512 2514
rect 52460 2450 52512 2456
rect 52472 1442 52500 2450
rect 52288 1414 52500 1442
rect 52288 800 52316 1414
rect 52564 800 52592 4626
rect 52644 4072 52696 4078
rect 52644 4014 52696 4020
rect 52656 1902 52684 4014
rect 52840 3942 52868 5510
rect 52932 4826 52960 36586
rect 53012 36168 53064 36174
rect 53012 36110 53064 36116
rect 53024 18834 53052 36110
rect 53932 35148 53984 35154
rect 53932 35090 53984 35096
rect 53104 34672 53156 34678
rect 53104 34614 53156 34620
rect 53116 34542 53144 34614
rect 53104 34536 53156 34542
rect 53104 34478 53156 34484
rect 53104 33924 53156 33930
rect 53104 33866 53156 33872
rect 53116 33454 53144 33866
rect 53104 33448 53156 33454
rect 53104 33390 53156 33396
rect 53748 32428 53800 32434
rect 53748 32370 53800 32376
rect 53760 32230 53788 32370
rect 53748 32224 53800 32230
rect 53748 32166 53800 32172
rect 53196 31816 53248 31822
rect 53196 31758 53248 31764
rect 53104 27396 53156 27402
rect 53104 27338 53156 27344
rect 53116 26314 53144 27338
rect 53104 26308 53156 26314
rect 53104 26250 53156 26256
rect 53208 25498 53236 31758
rect 53944 31754 53972 35090
rect 54116 35012 54168 35018
rect 54116 34954 54168 34960
rect 54128 34898 54156 34954
rect 54128 34870 54248 34898
rect 54220 34542 54248 34870
rect 54208 34536 54260 34542
rect 54208 34478 54260 34484
rect 53944 31726 54064 31754
rect 53748 31136 53800 31142
rect 53748 31078 53800 31084
rect 53760 30802 53788 31078
rect 53656 30796 53708 30802
rect 53656 30738 53708 30744
rect 53748 30796 53800 30802
rect 53748 30738 53800 30744
rect 53668 28558 53696 30738
rect 53838 30424 53894 30433
rect 53838 30359 53894 30368
rect 53748 29232 53800 29238
rect 53748 29174 53800 29180
rect 53656 28552 53708 28558
rect 53656 28494 53708 28500
rect 53760 27538 53788 29174
rect 53852 28966 53880 30359
rect 53840 28960 53892 28966
rect 53840 28902 53892 28908
rect 53840 28552 53892 28558
rect 53840 28494 53892 28500
rect 53288 27532 53340 27538
rect 53288 27474 53340 27480
rect 53380 27532 53432 27538
rect 53380 27474 53432 27480
rect 53748 27532 53800 27538
rect 53748 27474 53800 27480
rect 53300 27305 53328 27474
rect 53286 27296 53342 27305
rect 53286 27231 53342 27240
rect 53196 25492 53248 25498
rect 53196 25434 53248 25440
rect 53196 25356 53248 25362
rect 53196 25298 53248 25304
rect 53208 25158 53236 25298
rect 53196 25152 53248 25158
rect 53196 25094 53248 25100
rect 53104 22024 53156 22030
rect 53104 21966 53156 21972
rect 53116 21894 53144 21966
rect 53104 21888 53156 21894
rect 53104 21830 53156 21836
rect 53196 21888 53248 21894
rect 53196 21830 53248 21836
rect 53208 21418 53236 21830
rect 53196 21412 53248 21418
rect 53196 21354 53248 21360
rect 53104 20460 53156 20466
rect 53104 20402 53156 20408
rect 53116 19961 53144 20402
rect 53102 19952 53158 19961
rect 53102 19887 53158 19896
rect 53116 18834 53144 19887
rect 53012 18828 53064 18834
rect 53012 18770 53064 18776
rect 53104 18828 53156 18834
rect 53104 18770 53156 18776
rect 52920 4820 52972 4826
rect 52920 4762 52972 4768
rect 52828 3936 52880 3942
rect 52828 3878 52880 3884
rect 52736 3596 52788 3602
rect 52736 3538 52788 3544
rect 52644 1896 52696 1902
rect 52644 1838 52696 1844
rect 52748 800 52776 3538
rect 52920 1420 52972 1426
rect 52920 1362 52972 1368
rect 52932 800 52960 1362
rect 53024 882 53052 18770
rect 53288 16040 53340 16046
rect 53288 15982 53340 15988
rect 53300 14550 53328 15982
rect 53288 14544 53340 14550
rect 53288 14486 53340 14492
rect 53102 13968 53158 13977
rect 53102 13903 53104 13912
rect 53156 13903 53158 13912
rect 53104 13874 53156 13880
rect 53194 6352 53250 6361
rect 53194 6287 53250 6296
rect 53208 6254 53236 6287
rect 53196 6248 53248 6254
rect 53196 6190 53248 6196
rect 53392 4570 53420 27474
rect 53760 27441 53788 27474
rect 53852 27470 53880 28494
rect 53930 27704 53986 27713
rect 53930 27639 53932 27648
rect 53984 27639 53986 27648
rect 53932 27610 53984 27616
rect 53932 27532 53984 27538
rect 53932 27474 53984 27480
rect 53840 27464 53892 27470
rect 53746 27432 53802 27441
rect 53656 27396 53708 27402
rect 53840 27406 53892 27412
rect 53746 27367 53802 27376
rect 53656 27338 53708 27344
rect 53668 27305 53696 27338
rect 53944 27334 53972 27474
rect 53932 27328 53984 27334
rect 53654 27296 53710 27305
rect 53932 27270 53984 27276
rect 53654 27231 53710 27240
rect 53472 26920 53524 26926
rect 53472 26862 53524 26868
rect 53484 19786 53512 26862
rect 53838 26480 53894 26489
rect 53838 26415 53840 26424
rect 53892 26415 53894 26424
rect 53840 26386 53892 26392
rect 53748 26036 53800 26042
rect 53748 25978 53800 25984
rect 53654 25528 53710 25537
rect 53654 25463 53710 25472
rect 53668 25362 53696 25463
rect 53564 25356 53616 25362
rect 53564 25298 53616 25304
rect 53656 25356 53708 25362
rect 53656 25298 53708 25304
rect 53576 23798 53604 25298
rect 53760 25226 53788 25978
rect 54036 25378 54064 31726
rect 54208 31748 54260 31754
rect 54208 31690 54260 31696
rect 54220 31657 54248 31690
rect 54206 31648 54262 31657
rect 54206 31583 54262 31592
rect 54116 31408 54168 31414
rect 54116 31350 54168 31356
rect 54128 28665 54156 31350
rect 54208 30320 54260 30326
rect 54206 30288 54208 30297
rect 54260 30288 54262 30297
rect 54206 30223 54262 30232
rect 54114 28656 54170 28665
rect 54114 28591 54170 28600
rect 54128 27305 54156 28591
rect 54114 27296 54170 27305
rect 54114 27231 54170 27240
rect 53944 25350 54064 25378
rect 53748 25220 53800 25226
rect 53748 25162 53800 25168
rect 53564 23792 53616 23798
rect 53564 23734 53616 23740
rect 53472 19780 53524 19786
rect 53472 19722 53524 19728
rect 53576 9994 53604 23734
rect 53748 23180 53800 23186
rect 53748 23122 53800 23128
rect 53840 23180 53892 23186
rect 53840 23122 53892 23128
rect 53760 21486 53788 23122
rect 53852 22982 53880 23122
rect 53944 22982 53972 25350
rect 53840 22976 53892 22982
rect 53840 22918 53892 22924
rect 53932 22976 53984 22982
rect 53932 22918 53984 22924
rect 53748 21480 53800 21486
rect 53748 21422 53800 21428
rect 53746 20768 53802 20777
rect 53746 20703 53802 20712
rect 53656 17740 53708 17746
rect 53656 17682 53708 17688
rect 53668 14890 53696 17682
rect 53760 16674 53788 20703
rect 53944 20602 53972 22918
rect 54024 21548 54076 21554
rect 54128 21536 54156 27231
rect 54208 26920 54260 26926
rect 54208 26862 54260 26868
rect 54076 21508 54156 21536
rect 54024 21490 54076 21496
rect 53932 20596 53984 20602
rect 53932 20538 53984 20544
rect 54024 20596 54076 20602
rect 54024 20538 54076 20544
rect 54036 20346 54064 20538
rect 53944 20330 54064 20346
rect 54116 20392 54168 20398
rect 54116 20334 54168 20340
rect 53932 20324 54064 20330
rect 53984 20318 54064 20324
rect 53932 20266 53984 20272
rect 54128 20262 54156 20334
rect 54116 20256 54168 20262
rect 54116 20198 54168 20204
rect 54220 19990 54248 26862
rect 54208 19984 54260 19990
rect 54208 19926 54260 19932
rect 53760 16646 53972 16674
rect 53748 16584 53800 16590
rect 53748 16526 53800 16532
rect 53840 16584 53892 16590
rect 53840 16526 53892 16532
rect 53760 16250 53788 16526
rect 53748 16244 53800 16250
rect 53748 16186 53800 16192
rect 53748 16108 53800 16114
rect 53748 16050 53800 16056
rect 53656 14884 53708 14890
rect 53656 14826 53708 14832
rect 53564 9988 53616 9994
rect 53564 9930 53616 9936
rect 53656 7404 53708 7410
rect 53656 7346 53708 7352
rect 53668 6186 53696 7346
rect 53656 6180 53708 6186
rect 53656 6122 53708 6128
rect 53472 5840 53524 5846
rect 53472 5782 53524 5788
rect 53484 4690 53512 5782
rect 53668 4690 53696 6122
rect 53472 4684 53524 4690
rect 53472 4626 53524 4632
rect 53656 4684 53708 4690
rect 53656 4626 53708 4632
rect 53392 4542 53512 4570
rect 53484 4486 53512 4542
rect 53472 4480 53524 4486
rect 53472 4422 53524 4428
rect 53104 4072 53156 4078
rect 53104 4014 53156 4020
rect 53012 876 53064 882
rect 53012 818 53064 824
rect 53116 800 53144 4014
rect 53656 4004 53708 4010
rect 53656 3946 53708 3952
rect 53288 3596 53340 3602
rect 53288 3538 53340 3544
rect 53300 800 53328 3538
rect 53564 2848 53616 2854
rect 53564 2790 53616 2796
rect 53576 800 53604 2790
rect 53668 1034 53696 3946
rect 53760 2582 53788 16050
rect 53852 15162 53880 16526
rect 53944 16114 53972 16646
rect 53932 16108 53984 16114
rect 53932 16050 53984 16056
rect 54024 16108 54076 16114
rect 54024 16050 54076 16056
rect 54036 15706 54064 16050
rect 54024 15700 54076 15706
rect 54024 15642 54076 15648
rect 54312 15638 54340 38490
rect 54668 37324 54720 37330
rect 54668 37266 54720 37272
rect 54576 36644 54628 36650
rect 54576 36586 54628 36592
rect 54392 34944 54444 34950
rect 54392 34886 54444 34892
rect 54404 31754 54432 34886
rect 54588 34513 54616 36586
rect 54574 34504 54630 34513
rect 54574 34439 54630 34448
rect 54482 33688 54538 33697
rect 54482 33623 54538 33632
rect 54496 33522 54524 33623
rect 54484 33516 54536 33522
rect 54484 33458 54536 33464
rect 54404 31726 54524 31754
rect 54392 21548 54444 21554
rect 54392 21490 54444 21496
rect 53932 15632 53984 15638
rect 53932 15574 53984 15580
rect 54300 15632 54352 15638
rect 54300 15574 54352 15580
rect 53944 15473 53972 15574
rect 53930 15464 53986 15473
rect 54404 15450 54432 21490
rect 54496 20641 54524 31726
rect 54588 25945 54616 34439
rect 54680 30410 54708 37266
rect 54772 36922 54800 39200
rect 54944 37664 54996 37670
rect 54944 37606 54996 37612
rect 54760 36916 54812 36922
rect 54760 36858 54812 36864
rect 54850 36272 54906 36281
rect 54850 36207 54852 36216
rect 54904 36207 54906 36216
rect 54852 36178 54904 36184
rect 54758 35456 54814 35465
rect 54758 35391 54814 35400
rect 54772 31414 54800 35391
rect 54852 34468 54904 34474
rect 54852 34410 54904 34416
rect 54760 31408 54812 31414
rect 54760 31350 54812 31356
rect 54772 31278 54800 31350
rect 54760 31272 54812 31278
rect 54760 31214 54812 31220
rect 54680 30382 54800 30410
rect 54668 30184 54720 30190
rect 54668 30126 54720 30132
rect 54680 30025 54708 30126
rect 54666 30016 54722 30025
rect 54666 29951 54722 29960
rect 54574 25936 54630 25945
rect 54574 25871 54630 25880
rect 54576 25492 54628 25498
rect 54576 25434 54628 25440
rect 54482 20632 54538 20641
rect 54482 20567 54538 20576
rect 54484 20460 54536 20466
rect 54484 20402 54536 20408
rect 54496 19922 54524 20402
rect 54484 19916 54536 19922
rect 54484 19858 54536 19864
rect 54484 15564 54536 15570
rect 54484 15506 54536 15512
rect 53930 15399 53986 15408
rect 54128 15422 54432 15450
rect 54024 15360 54076 15366
rect 54024 15302 54076 15308
rect 53840 15156 53892 15162
rect 53840 15098 53892 15104
rect 53932 9512 53984 9518
rect 53932 9454 53984 9460
rect 53840 8424 53892 8430
rect 53840 8366 53892 8372
rect 53748 2576 53800 2582
rect 53748 2518 53800 2524
rect 53852 1970 53880 8366
rect 53944 3942 53972 9454
rect 54036 7546 54064 15302
rect 54024 7540 54076 7546
rect 54024 7482 54076 7488
rect 53932 3936 53984 3942
rect 53932 3878 53984 3884
rect 53932 3596 53984 3602
rect 53932 3538 53984 3544
rect 53840 1964 53892 1970
rect 53840 1906 53892 1912
rect 53668 1006 53788 1034
rect 53760 800 53788 1006
rect 53944 800 53972 3538
rect 54024 3392 54076 3398
rect 54024 3334 54076 3340
rect 54036 2990 54064 3334
rect 54024 2984 54076 2990
rect 54024 2926 54076 2932
rect 54024 2644 54076 2650
rect 54024 2586 54076 2592
rect 54036 1426 54064 2586
rect 54128 2582 54156 15422
rect 54300 15360 54352 15366
rect 54300 15302 54352 15308
rect 54312 14958 54340 15302
rect 54300 14952 54352 14958
rect 54300 14894 54352 14900
rect 54312 13258 54340 14894
rect 54300 13252 54352 13258
rect 54300 13194 54352 13200
rect 54300 12708 54352 12714
rect 54300 12650 54352 12656
rect 54312 9586 54340 12650
rect 54300 9580 54352 9586
rect 54300 9522 54352 9528
rect 54496 9178 54524 15506
rect 54484 9172 54536 9178
rect 54484 9114 54536 9120
rect 54392 7540 54444 7546
rect 54392 7482 54444 7488
rect 54300 4684 54352 4690
rect 54300 4626 54352 4632
rect 54116 2576 54168 2582
rect 54116 2518 54168 2524
rect 54116 2372 54168 2378
rect 54116 2314 54168 2320
rect 54024 1420 54076 1426
rect 54024 1362 54076 1368
rect 54128 800 54156 2314
rect 54312 800 54340 4626
rect 54404 2038 54432 7482
rect 54588 5166 54616 25434
rect 54772 25158 54800 30382
rect 54760 25152 54812 25158
rect 54760 25094 54812 25100
rect 54668 22432 54720 22438
rect 54668 22374 54720 22380
rect 54680 22166 54708 22374
rect 54668 22160 54720 22166
rect 54668 22102 54720 22108
rect 54680 19922 54708 22102
rect 54864 22094 54892 34410
rect 54956 26926 54984 37606
rect 55404 37392 55456 37398
rect 55404 37334 55456 37340
rect 55220 36916 55272 36922
rect 55220 36858 55272 36864
rect 55128 36168 55180 36174
rect 55128 36110 55180 36116
rect 55140 34474 55168 36110
rect 55128 34468 55180 34474
rect 55128 34410 55180 34416
rect 55034 34096 55090 34105
rect 55034 34031 55090 34040
rect 55048 33862 55076 34031
rect 55036 33856 55088 33862
rect 55036 33798 55088 33804
rect 55036 32564 55088 32570
rect 55036 32506 55088 32512
rect 55048 31754 55076 32506
rect 55036 31748 55088 31754
rect 55036 31690 55088 31696
rect 55036 31272 55088 31278
rect 55036 31214 55088 31220
rect 55048 30433 55076 31214
rect 55232 30666 55260 36858
rect 55312 36236 55364 36242
rect 55312 36178 55364 36184
rect 55324 36038 55352 36178
rect 55312 36032 55364 36038
rect 55312 35974 55364 35980
rect 55324 35737 55352 35974
rect 55310 35728 55366 35737
rect 55310 35663 55366 35672
rect 55310 35592 55366 35601
rect 55310 35527 55312 35536
rect 55364 35527 55366 35536
rect 55312 35498 55364 35504
rect 55310 34504 55366 34513
rect 55310 34439 55312 34448
rect 55364 34439 55366 34448
rect 55312 34410 55364 34416
rect 55310 33688 55366 33697
rect 55310 33623 55366 33632
rect 55324 33386 55352 33623
rect 55312 33380 55364 33386
rect 55312 33322 55364 33328
rect 55312 31272 55364 31278
rect 55312 31214 55364 31220
rect 55324 31142 55352 31214
rect 55312 31136 55364 31142
rect 55312 31078 55364 31084
rect 55220 30660 55272 30666
rect 55220 30602 55272 30608
rect 55034 30424 55090 30433
rect 55034 30359 55090 30368
rect 55128 30320 55180 30326
rect 55128 30262 55180 30268
rect 55140 30190 55168 30262
rect 55128 30184 55180 30190
rect 55128 30126 55180 30132
rect 55220 30184 55272 30190
rect 55220 30126 55272 30132
rect 55036 30116 55088 30122
rect 55036 30058 55088 30064
rect 55048 29850 55076 30058
rect 55036 29844 55088 29850
rect 55036 29786 55088 29792
rect 55034 27160 55090 27169
rect 55034 27095 55090 27104
rect 55048 26926 55076 27095
rect 54944 26920 54996 26926
rect 54944 26862 54996 26868
rect 55036 26920 55088 26926
rect 55036 26862 55088 26868
rect 55034 23216 55090 23225
rect 55034 23151 55090 23160
rect 54864 22066 54984 22094
rect 54758 20632 54814 20641
rect 54758 20567 54814 20576
rect 54668 19916 54720 19922
rect 54668 19858 54720 19864
rect 54772 19174 54800 20567
rect 54760 19168 54812 19174
rect 54760 19110 54812 19116
rect 54852 18624 54904 18630
rect 54852 18566 54904 18572
rect 54760 15564 54812 15570
rect 54760 15506 54812 15512
rect 54772 15026 54800 15506
rect 54760 15020 54812 15026
rect 54760 14962 54812 14968
rect 54772 14482 54800 14962
rect 54760 14476 54812 14482
rect 54760 14418 54812 14424
rect 54864 13802 54892 18566
rect 54956 14482 54984 22066
rect 55048 21690 55076 23151
rect 55128 22976 55180 22982
rect 55128 22918 55180 22924
rect 55140 22438 55168 22918
rect 55128 22432 55180 22438
rect 55128 22374 55180 22380
rect 55036 21684 55088 21690
rect 55036 21626 55088 21632
rect 55034 21584 55090 21593
rect 55034 21519 55090 21528
rect 55048 21418 55076 21519
rect 55036 21412 55088 21418
rect 55036 21354 55088 21360
rect 55128 19916 55180 19922
rect 55128 19858 55180 19864
rect 55036 19712 55088 19718
rect 55036 19654 55088 19660
rect 54944 14476 54996 14482
rect 54944 14418 54996 14424
rect 54852 13796 54904 13802
rect 54852 13738 54904 13744
rect 54852 12980 54904 12986
rect 54852 12922 54904 12928
rect 54668 12368 54720 12374
rect 54668 12310 54720 12316
rect 54680 12102 54708 12310
rect 54668 12096 54720 12102
rect 54668 12038 54720 12044
rect 54680 7750 54708 12038
rect 54760 9580 54812 9586
rect 54760 9522 54812 9528
rect 54668 7744 54720 7750
rect 54668 7686 54720 7692
rect 54772 6934 54800 9522
rect 54760 6928 54812 6934
rect 54760 6870 54812 6876
rect 54576 5160 54628 5166
rect 54576 5102 54628 5108
rect 54576 3596 54628 3602
rect 54576 3538 54628 3544
rect 54392 2032 54444 2038
rect 54392 1974 54444 1980
rect 54588 800 54616 3538
rect 54760 2848 54812 2854
rect 54760 2790 54812 2796
rect 54772 800 54800 2790
rect 50804 604 50856 610
rect 50804 546 50856 552
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54864 542 54892 12922
rect 54944 4072 54996 4078
rect 54944 4014 54996 4020
rect 54956 800 54984 4014
rect 55048 2582 55076 19654
rect 55140 15570 55168 19858
rect 55128 15564 55180 15570
rect 55128 15506 55180 15512
rect 55128 14408 55180 14414
rect 55128 14350 55180 14356
rect 55140 12986 55168 14350
rect 55128 12980 55180 12986
rect 55128 12922 55180 12928
rect 55128 9920 55180 9926
rect 55128 9862 55180 9868
rect 55140 4758 55168 9862
rect 55128 4752 55180 4758
rect 55128 4694 55180 4700
rect 55128 3596 55180 3602
rect 55128 3538 55180 3544
rect 55036 2576 55088 2582
rect 55036 2518 55088 2524
rect 55140 800 55168 3538
rect 55232 3058 55260 30126
rect 55310 29064 55366 29073
rect 55310 28999 55312 29008
rect 55364 28999 55366 29008
rect 55312 28970 55364 28976
rect 55312 22568 55364 22574
rect 55312 22510 55364 22516
rect 55324 12434 55352 22510
rect 55416 15570 55444 37334
rect 55508 36310 55536 39374
rect 55586 39200 55642 40000
rect 56506 39200 56562 40000
rect 57334 39200 57390 40000
rect 58254 39200 58310 40000
rect 59082 39200 59138 40000
rect 60002 39200 60058 40000
rect 60830 39200 60886 40000
rect 61108 39364 61160 39370
rect 61108 39306 61160 39312
rect 55600 36718 55628 39200
rect 56048 37868 56100 37874
rect 56048 37810 56100 37816
rect 55680 37324 55732 37330
rect 55680 37266 55732 37272
rect 55588 36712 55640 36718
rect 55588 36654 55640 36660
rect 55496 36304 55548 36310
rect 55496 36246 55548 36252
rect 55588 36168 55640 36174
rect 55588 36110 55640 36116
rect 55600 36038 55628 36110
rect 55588 36032 55640 36038
rect 55588 35974 55640 35980
rect 55588 35760 55640 35766
rect 55588 35702 55640 35708
rect 55496 35624 55548 35630
rect 55496 35566 55548 35572
rect 55508 30598 55536 35566
rect 55600 35154 55628 35702
rect 55588 35148 55640 35154
rect 55588 35090 55640 35096
rect 55692 31686 55720 37266
rect 55772 36576 55824 36582
rect 55772 36518 55824 36524
rect 55784 36378 55812 36518
rect 55772 36372 55824 36378
rect 55772 36314 55824 36320
rect 55864 36304 55916 36310
rect 55862 36272 55864 36281
rect 55916 36272 55918 36281
rect 55862 36207 55918 36216
rect 55956 36168 56008 36174
rect 55956 36110 56008 36116
rect 55864 36100 55916 36106
rect 55864 36042 55916 36048
rect 55772 35624 55824 35630
rect 55876 35601 55904 36042
rect 55968 36009 55996 36110
rect 55954 36000 56010 36009
rect 55954 35935 56010 35944
rect 56060 35630 56088 37810
rect 56520 37466 56548 39200
rect 56508 37460 56560 37466
rect 56508 37402 56560 37408
rect 57348 36922 57376 39200
rect 57796 38072 57848 38078
rect 57796 38014 57848 38020
rect 57808 37466 57836 38014
rect 57796 37460 57848 37466
rect 57796 37402 57848 37408
rect 58268 37398 58296 39200
rect 59096 37466 59124 39200
rect 59452 39160 59504 39166
rect 59452 39102 59504 39108
rect 59084 37460 59136 37466
rect 59084 37402 59136 37408
rect 58256 37392 58308 37398
rect 58256 37334 58308 37340
rect 58440 37324 58492 37330
rect 58440 37266 58492 37272
rect 58900 37324 58952 37330
rect 58900 37266 58952 37272
rect 57336 36916 57388 36922
rect 57336 36858 57388 36864
rect 57428 36644 57480 36650
rect 57428 36586 57480 36592
rect 56324 36576 56376 36582
rect 56324 36518 56376 36524
rect 56508 36576 56560 36582
rect 56508 36518 56560 36524
rect 55956 35624 56008 35630
rect 55772 35566 55824 35572
rect 55862 35592 55918 35601
rect 55784 35465 55812 35566
rect 55956 35566 56008 35572
rect 56048 35624 56100 35630
rect 56048 35566 56100 35572
rect 55862 35527 55918 35536
rect 55770 35456 55826 35465
rect 55770 35391 55826 35400
rect 55772 32360 55824 32366
rect 55772 32302 55824 32308
rect 55864 32360 55916 32366
rect 55864 32302 55916 32308
rect 55680 31680 55732 31686
rect 55680 31622 55732 31628
rect 55680 31136 55732 31142
rect 55600 31096 55680 31124
rect 55496 30592 55548 30598
rect 55496 30534 55548 30540
rect 55496 29640 55548 29646
rect 55496 29582 55548 29588
rect 55508 29034 55536 29582
rect 55496 29028 55548 29034
rect 55496 28970 55548 28976
rect 55600 28914 55628 31096
rect 55680 31078 55732 31084
rect 55680 30048 55732 30054
rect 55680 29990 55732 29996
rect 55692 29646 55720 29990
rect 55680 29640 55732 29646
rect 55680 29582 55732 29588
rect 55508 28886 55628 28914
rect 55680 28960 55732 28966
rect 55680 28902 55732 28908
rect 55508 23118 55536 28886
rect 55692 28626 55720 28902
rect 55680 28620 55732 28626
rect 55680 28562 55732 28568
rect 55680 27328 55732 27334
rect 55680 27270 55732 27276
rect 55692 27130 55720 27270
rect 55680 27124 55732 27130
rect 55680 27066 55732 27072
rect 55586 26616 55642 26625
rect 55586 26551 55642 26560
rect 55496 23112 55548 23118
rect 55496 23054 55548 23060
rect 55508 22982 55536 23054
rect 55496 22976 55548 22982
rect 55496 22918 55548 22924
rect 55496 22092 55548 22098
rect 55496 22034 55548 22040
rect 55404 15564 55456 15570
rect 55404 15506 55456 15512
rect 55416 14226 55444 15506
rect 55508 14482 55536 22034
rect 55496 14476 55548 14482
rect 55496 14418 55548 14424
rect 55600 14346 55628 26551
rect 55680 24676 55732 24682
rect 55680 24618 55732 24624
rect 55692 24138 55720 24618
rect 55680 24132 55732 24138
rect 55680 24074 55732 24080
rect 55680 23112 55732 23118
rect 55680 23054 55732 23060
rect 55692 22778 55720 23054
rect 55680 22772 55732 22778
rect 55680 22714 55732 22720
rect 55784 22098 55812 32302
rect 55772 22092 55824 22098
rect 55772 22034 55824 22040
rect 55680 21480 55732 21486
rect 55876 21434 55904 32302
rect 55680 21422 55732 21428
rect 55692 20874 55720 21422
rect 55784 21406 55904 21434
rect 55680 20868 55732 20874
rect 55680 20810 55732 20816
rect 55680 19916 55732 19922
rect 55680 19858 55732 19864
rect 55692 15094 55720 19858
rect 55784 18873 55812 21406
rect 55864 21344 55916 21350
rect 55864 21286 55916 21292
rect 55876 21146 55904 21286
rect 55864 21140 55916 21146
rect 55864 21082 55916 21088
rect 55864 20868 55916 20874
rect 55864 20810 55916 20816
rect 55876 20777 55904 20810
rect 55862 20768 55918 20777
rect 55862 20703 55918 20712
rect 55864 19168 55916 19174
rect 55864 19110 55916 19116
rect 55876 18970 55904 19110
rect 55864 18964 55916 18970
rect 55864 18906 55916 18912
rect 55770 18864 55826 18873
rect 55770 18799 55826 18808
rect 55772 16108 55824 16114
rect 55772 16050 55824 16056
rect 55784 15638 55812 16050
rect 55862 16008 55918 16017
rect 55862 15943 55918 15952
rect 55876 15706 55904 15943
rect 55864 15700 55916 15706
rect 55864 15642 55916 15648
rect 55772 15632 55824 15638
rect 55772 15574 55824 15580
rect 55862 15600 55918 15609
rect 55862 15535 55918 15544
rect 55876 15502 55904 15535
rect 55864 15496 55916 15502
rect 55770 15464 55826 15473
rect 55864 15438 55916 15444
rect 55770 15399 55772 15408
rect 55824 15399 55826 15408
rect 55772 15370 55824 15376
rect 55864 15156 55916 15162
rect 55864 15098 55916 15104
rect 55680 15088 55732 15094
rect 55680 15030 55732 15036
rect 55876 14618 55904 15098
rect 55864 14612 55916 14618
rect 55864 14554 55916 14560
rect 55588 14340 55640 14346
rect 55588 14282 55640 14288
rect 55416 14198 55628 14226
rect 55600 12434 55628 14198
rect 55680 13864 55732 13870
rect 55680 13806 55732 13812
rect 55324 12406 55444 12434
rect 55312 8900 55364 8906
rect 55312 8842 55364 8848
rect 55324 4690 55352 8842
rect 55312 4684 55364 4690
rect 55312 4626 55364 4632
rect 55220 3052 55272 3058
rect 55220 2994 55272 3000
rect 55312 2916 55364 2922
rect 55312 2858 55364 2864
rect 55324 800 55352 2858
rect 55416 2582 55444 12406
rect 55508 12406 55628 12434
rect 55508 11150 55536 12406
rect 55496 11144 55548 11150
rect 55496 11086 55548 11092
rect 55588 8900 55640 8906
rect 55588 8842 55640 8848
rect 55600 8566 55628 8842
rect 55588 8560 55640 8566
rect 55588 8502 55640 8508
rect 55692 7562 55720 13806
rect 55772 13796 55824 13802
rect 55772 13738 55824 13744
rect 55784 12782 55812 13738
rect 55772 12776 55824 12782
rect 55772 12718 55824 12724
rect 55508 7534 55720 7562
rect 55404 2576 55456 2582
rect 55404 2518 55456 2524
rect 54852 536 54904 542
rect 54852 478 54904 484
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55508 785 55536 7534
rect 55680 6792 55732 6798
rect 55680 6734 55732 6740
rect 55588 4072 55640 4078
rect 55588 4014 55640 4020
rect 55600 800 55628 4014
rect 55692 3942 55720 6734
rect 55784 5302 55812 12718
rect 55968 12238 55996 35566
rect 56336 35290 56364 36518
rect 56324 35284 56376 35290
rect 56324 35226 56376 35232
rect 56140 33516 56192 33522
rect 56140 33458 56192 33464
rect 56152 33017 56180 33458
rect 56138 33008 56194 33017
rect 56138 32943 56194 32952
rect 56048 32904 56100 32910
rect 56048 32846 56100 32852
rect 56060 32298 56088 32846
rect 56140 32360 56192 32366
rect 56140 32302 56192 32308
rect 56416 32360 56468 32366
rect 56416 32302 56468 32308
rect 56048 32292 56100 32298
rect 56048 32234 56100 32240
rect 56152 31754 56180 32302
rect 56232 31816 56284 31822
rect 56232 31758 56284 31764
rect 56060 31726 56180 31754
rect 56060 31142 56088 31726
rect 56244 31686 56272 31758
rect 56140 31680 56192 31686
rect 56140 31622 56192 31628
rect 56232 31680 56284 31686
rect 56232 31622 56284 31628
rect 56048 31136 56100 31142
rect 56048 31078 56100 31084
rect 56046 27296 56102 27305
rect 56046 27231 56102 27240
rect 56060 27062 56088 27231
rect 56048 27056 56100 27062
rect 56048 26998 56100 27004
rect 56048 25832 56100 25838
rect 56048 25774 56100 25780
rect 56060 25294 56088 25774
rect 56048 25288 56100 25294
rect 56048 25230 56100 25236
rect 56048 23316 56100 23322
rect 56048 23258 56100 23264
rect 56060 22778 56088 23258
rect 56152 23186 56180 31622
rect 56232 31136 56284 31142
rect 56232 31078 56284 31084
rect 56244 26625 56272 31078
rect 56324 28620 56376 28626
rect 56324 28562 56376 28568
rect 56336 28490 56364 28562
rect 56324 28484 56376 28490
rect 56324 28426 56376 28432
rect 56230 26616 56286 26625
rect 56230 26551 56286 26560
rect 56232 25900 56284 25906
rect 56232 25842 56284 25848
rect 56244 25673 56272 25842
rect 56230 25664 56286 25673
rect 56230 25599 56286 25608
rect 56324 25492 56376 25498
rect 56324 25434 56376 25440
rect 56232 25356 56284 25362
rect 56232 25298 56284 25304
rect 56244 24886 56272 25298
rect 56336 24886 56364 25434
rect 56232 24880 56284 24886
rect 56232 24822 56284 24828
rect 56324 24880 56376 24886
rect 56324 24822 56376 24828
rect 56232 23316 56284 23322
rect 56232 23258 56284 23264
rect 56140 23180 56192 23186
rect 56140 23122 56192 23128
rect 56048 22772 56100 22778
rect 56048 22714 56100 22720
rect 56152 22094 56180 23122
rect 56244 22982 56272 23258
rect 56232 22976 56284 22982
rect 56232 22918 56284 22924
rect 56152 22066 56272 22094
rect 56140 21956 56192 21962
rect 56140 21898 56192 21904
rect 56152 20369 56180 21898
rect 56138 20360 56194 20369
rect 56138 20295 56194 20304
rect 56048 18828 56100 18834
rect 56048 18770 56100 18776
rect 56060 18290 56088 18770
rect 56048 18284 56100 18290
rect 56048 18226 56100 18232
rect 56140 18284 56192 18290
rect 56140 18226 56192 18232
rect 56048 16516 56100 16522
rect 56048 16458 56100 16464
rect 56060 16182 56088 16458
rect 56048 16176 56100 16182
rect 56048 16118 56100 16124
rect 56048 16040 56100 16046
rect 56048 15982 56100 15988
rect 56060 13870 56088 15982
rect 56048 13864 56100 13870
rect 56048 13806 56100 13812
rect 56048 12436 56100 12442
rect 56048 12378 56100 12384
rect 55864 12232 55916 12238
rect 55864 12174 55916 12180
rect 55956 12232 56008 12238
rect 55956 12174 56008 12180
rect 55876 12084 55904 12174
rect 56060 12084 56088 12378
rect 55876 12056 56088 12084
rect 55864 11348 55916 11354
rect 55864 11290 55916 11296
rect 55876 11218 55904 11290
rect 55864 11212 55916 11218
rect 55864 11154 55916 11160
rect 55956 5364 56008 5370
rect 55956 5306 56008 5312
rect 55772 5296 55824 5302
rect 55968 5250 55996 5306
rect 55772 5238 55824 5244
rect 55876 5234 55996 5250
rect 55864 5228 55996 5234
rect 55916 5222 55996 5228
rect 55864 5170 55916 5176
rect 55772 4140 55824 4146
rect 55772 4082 55824 4088
rect 55680 3936 55732 3942
rect 55680 3878 55732 3884
rect 55784 3466 55812 4082
rect 55772 3460 55824 3466
rect 55772 3402 55824 3408
rect 55772 2916 55824 2922
rect 55772 2858 55824 2864
rect 55784 800 55812 2858
rect 56152 2582 56180 18226
rect 56244 14618 56272 22066
rect 56428 18970 56456 32302
rect 56520 29238 56548 36518
rect 56600 36236 56652 36242
rect 56600 36178 56652 36184
rect 56612 30297 56640 36178
rect 57152 35828 57204 35834
rect 57152 35770 57204 35776
rect 56692 35692 56744 35698
rect 56692 35634 56744 35640
rect 56704 35222 56732 35634
rect 57164 35630 57192 35770
rect 57242 35728 57298 35737
rect 57242 35663 57298 35672
rect 57152 35624 57204 35630
rect 57152 35566 57204 35572
rect 56782 35456 56838 35465
rect 56782 35391 56838 35400
rect 56796 35222 56824 35391
rect 56692 35216 56744 35222
rect 56692 35158 56744 35164
rect 56784 35216 56836 35222
rect 56784 35158 56836 35164
rect 57152 34944 57204 34950
rect 57152 34886 57204 34892
rect 56784 32496 56836 32502
rect 56784 32438 56836 32444
rect 56796 31657 56824 32438
rect 56782 31648 56838 31657
rect 56782 31583 56838 31592
rect 56598 30288 56654 30297
rect 56598 30223 56654 30232
rect 56508 29232 56560 29238
rect 56508 29174 56560 29180
rect 56508 25492 56560 25498
rect 56508 25434 56560 25440
rect 56520 25158 56548 25434
rect 56508 25152 56560 25158
rect 56508 25094 56560 25100
rect 56612 19990 56640 30223
rect 57164 30025 57192 34886
rect 57150 30016 57206 30025
rect 57150 29951 57206 29960
rect 57164 29238 57192 29951
rect 57152 29232 57204 29238
rect 57152 29174 57204 29180
rect 56690 29064 56746 29073
rect 56690 28999 56746 29008
rect 56600 19984 56652 19990
rect 56600 19926 56652 19932
rect 56612 19446 56640 19926
rect 56508 19440 56560 19446
rect 56508 19382 56560 19388
rect 56600 19440 56652 19446
rect 56600 19382 56652 19388
rect 56416 18964 56468 18970
rect 56416 18906 56468 18912
rect 56428 18222 56456 18906
rect 56520 18426 56548 19382
rect 56508 18420 56560 18426
rect 56508 18362 56560 18368
rect 56416 18216 56468 18222
rect 56416 18158 56468 18164
rect 56416 17536 56468 17542
rect 56416 17478 56468 17484
rect 56428 17134 56456 17478
rect 56416 17128 56468 17134
rect 56416 17070 56468 17076
rect 56520 16658 56548 18362
rect 56600 17536 56652 17542
rect 56600 17478 56652 17484
rect 56508 16652 56560 16658
rect 56508 16594 56560 16600
rect 56324 16040 56376 16046
rect 56324 15982 56376 15988
rect 56508 16040 56560 16046
rect 56508 15982 56560 15988
rect 56232 14612 56284 14618
rect 56232 14554 56284 14560
rect 56336 12434 56364 15982
rect 56520 15570 56548 15982
rect 56508 15564 56560 15570
rect 56508 15506 56560 15512
rect 56508 13796 56560 13802
rect 56508 13738 56560 13744
rect 56336 12406 56456 12434
rect 56232 7744 56284 7750
rect 56232 7686 56284 7692
rect 56244 5234 56272 7686
rect 56232 5228 56284 5234
rect 56232 5170 56284 5176
rect 56232 4072 56284 4078
rect 56232 4014 56284 4020
rect 56140 2576 56192 2582
rect 56140 2518 56192 2524
rect 55956 2440 56008 2446
rect 55956 2382 56008 2388
rect 55968 800 55996 2382
rect 56244 1442 56272 4014
rect 56324 3596 56376 3602
rect 56324 3538 56376 3544
rect 56152 1414 56272 1442
rect 56152 800 56180 1414
rect 56336 800 56364 3538
rect 56428 2106 56456 12406
rect 56520 12102 56548 13738
rect 56508 12096 56560 12102
rect 56508 12038 56560 12044
rect 56612 11830 56640 17478
rect 56600 11824 56652 11830
rect 56600 11766 56652 11772
rect 56506 8800 56562 8809
rect 56506 8735 56562 8744
rect 56520 8566 56548 8735
rect 56600 8628 56652 8634
rect 56600 8570 56652 8576
rect 56508 8560 56560 8566
rect 56508 8502 56560 8508
rect 56612 6730 56640 8570
rect 56600 6724 56652 6730
rect 56600 6666 56652 6672
rect 56704 2990 56732 28999
rect 56968 28484 57020 28490
rect 56968 28426 57020 28432
rect 56874 25256 56930 25265
rect 56784 25220 56836 25226
rect 56874 25191 56930 25200
rect 56784 25162 56836 25168
rect 56796 9110 56824 25162
rect 56888 25158 56916 25191
rect 56876 25152 56928 25158
rect 56876 25094 56928 25100
rect 56980 21894 57008 28426
rect 56968 21888 57020 21894
rect 56968 21830 57020 21836
rect 57152 17196 57204 17202
rect 57152 17138 57204 17144
rect 57164 16726 57192 17138
rect 57152 16720 57204 16726
rect 57152 16662 57204 16668
rect 57256 14550 57284 35663
rect 57440 35193 57468 36586
rect 57426 35184 57482 35193
rect 57426 35119 57482 35128
rect 57336 29232 57388 29238
rect 57336 29174 57388 29180
rect 57244 14544 57296 14550
rect 57244 14486 57296 14492
rect 56874 13968 56930 13977
rect 56874 13903 56876 13912
rect 56928 13903 56930 13912
rect 56876 13874 56928 13880
rect 57348 10538 57376 29174
rect 57440 21078 57468 35119
rect 58164 34128 58216 34134
rect 58164 34070 58216 34076
rect 58072 33856 58124 33862
rect 58072 33798 58124 33804
rect 58084 32434 58112 33798
rect 58176 32570 58204 34070
rect 58164 32564 58216 32570
rect 58164 32506 58216 32512
rect 58072 32428 58124 32434
rect 58072 32370 58124 32376
rect 57978 32192 58034 32201
rect 57978 32127 58034 32136
rect 57886 32056 57942 32065
rect 57886 31991 57942 32000
rect 57518 31920 57574 31929
rect 57900 31890 57928 31991
rect 57992 31890 58020 32127
rect 58084 32026 58296 32042
rect 58072 32020 58308 32026
rect 58124 32014 58256 32020
rect 58072 31962 58124 31968
rect 58256 31962 58308 31968
rect 58162 31920 58218 31929
rect 57518 31855 57574 31864
rect 57888 31884 57940 31890
rect 57532 31754 57560 31855
rect 57888 31826 57940 31832
rect 57980 31884 58032 31890
rect 58162 31855 58164 31864
rect 57980 31826 58032 31832
rect 58216 31855 58218 31864
rect 58164 31826 58216 31832
rect 57886 31784 57942 31793
rect 57520 31748 57572 31754
rect 57942 31754 58112 31770
rect 57942 31748 58400 31754
rect 57942 31742 58348 31748
rect 57886 31719 57942 31728
rect 58084 31726 58348 31742
rect 57520 31690 57572 31696
rect 58348 31690 58400 31696
rect 58072 31680 58124 31686
rect 58072 31622 58124 31628
rect 57520 31204 57572 31210
rect 57520 31146 57572 31152
rect 57532 30938 57560 31146
rect 57520 30932 57572 30938
rect 57520 30874 57572 30880
rect 58084 30122 58112 31622
rect 58072 30116 58124 30122
rect 58072 30058 58124 30064
rect 57520 29232 57572 29238
rect 57520 29174 57572 29180
rect 57532 26897 57560 29174
rect 57518 26888 57574 26897
rect 57518 26823 57574 26832
rect 57532 25226 57560 26823
rect 57888 26444 57940 26450
rect 57888 26386 57940 26392
rect 57520 25220 57572 25226
rect 57520 25162 57572 25168
rect 57428 21072 57480 21078
rect 57428 21014 57480 21020
rect 57520 19712 57572 19718
rect 57520 19654 57572 19660
rect 57532 19446 57560 19654
rect 57428 19440 57480 19446
rect 57428 19382 57480 19388
rect 57520 19440 57572 19446
rect 57520 19382 57572 19388
rect 57440 12374 57468 19382
rect 57520 17128 57572 17134
rect 57520 17070 57572 17076
rect 57532 16726 57560 17070
rect 57520 16720 57572 16726
rect 57520 16662 57572 16668
rect 57796 14952 57848 14958
rect 57794 14920 57796 14929
rect 57848 14920 57850 14929
rect 57794 14855 57850 14864
rect 57796 14544 57848 14550
rect 57796 14486 57848 14492
rect 57428 12368 57480 12374
rect 57428 12310 57480 12316
rect 57704 12096 57756 12102
rect 57704 12038 57756 12044
rect 57336 10532 57388 10538
rect 57336 10474 57388 10480
rect 57348 9518 57376 10474
rect 57336 9512 57388 9518
rect 57336 9454 57388 9460
rect 56784 9104 56836 9110
rect 56784 9046 56836 9052
rect 56796 8906 56824 9046
rect 56784 8900 56836 8906
rect 56784 8842 56836 8848
rect 56876 7744 56928 7750
rect 56876 7686 56928 7692
rect 56784 4072 56836 4078
rect 56784 4014 56836 4020
rect 56692 2984 56744 2990
rect 56692 2926 56744 2932
rect 56600 2848 56652 2854
rect 56600 2790 56652 2796
rect 56416 2100 56468 2106
rect 56416 2042 56468 2048
rect 56612 800 56640 2790
rect 56796 800 56824 4014
rect 56888 3398 56916 7686
rect 57716 7478 57744 12038
rect 57808 10062 57836 14486
rect 57796 10056 57848 10062
rect 57796 9998 57848 10004
rect 57704 7472 57756 7478
rect 57704 7414 57756 7420
rect 57900 5302 57928 26386
rect 58452 19310 58480 37266
rect 58624 34468 58676 34474
rect 58624 34410 58676 34416
rect 58636 34134 58664 34410
rect 58624 34128 58676 34134
rect 58624 34070 58676 34076
rect 58716 33380 58768 33386
rect 58716 33322 58768 33328
rect 58532 32836 58584 32842
rect 58532 32778 58584 32784
rect 58544 31890 58572 32778
rect 58532 31884 58584 31890
rect 58532 31826 58584 31832
rect 58530 29608 58586 29617
rect 58530 29543 58586 29552
rect 58440 19304 58492 19310
rect 58440 19246 58492 19252
rect 57980 16788 58032 16794
rect 57980 16730 58032 16736
rect 57992 13802 58020 16730
rect 58072 16584 58124 16590
rect 58072 16526 58124 16532
rect 58084 15638 58112 16526
rect 58072 15632 58124 15638
rect 58072 15574 58124 15580
rect 58452 14958 58480 19246
rect 58544 18442 58572 29543
rect 58624 21888 58676 21894
rect 58624 21830 58676 21836
rect 58636 21554 58664 21830
rect 58624 21548 58676 21554
rect 58624 21490 58676 21496
rect 58622 20632 58678 20641
rect 58622 20567 58678 20576
rect 58636 19310 58664 20567
rect 58624 19304 58676 19310
rect 58624 19246 58676 19252
rect 58544 18414 58664 18442
rect 58532 16788 58584 16794
rect 58532 16730 58584 16736
rect 58544 15570 58572 16730
rect 58532 15564 58584 15570
rect 58532 15506 58584 15512
rect 58348 14952 58400 14958
rect 58346 14920 58348 14929
rect 58440 14952 58492 14958
rect 58400 14920 58402 14929
rect 58440 14894 58492 14900
rect 58346 14855 58402 14864
rect 57980 13796 58032 13802
rect 57980 13738 58032 13744
rect 58636 12714 58664 18414
rect 58728 17134 58756 33322
rect 58806 32056 58862 32065
rect 58806 31991 58862 32000
rect 58820 31958 58848 31991
rect 58808 31952 58860 31958
rect 58808 31894 58860 31900
rect 58912 31754 58940 37266
rect 59360 36168 59412 36174
rect 59360 36110 59412 36116
rect 59372 35290 59400 36110
rect 59360 35284 59412 35290
rect 59360 35226 59412 35232
rect 59360 34944 59412 34950
rect 59360 34886 59412 34892
rect 59372 34542 59400 34886
rect 59360 34536 59412 34542
rect 59360 34478 59412 34484
rect 59464 34354 59492 39102
rect 60016 36922 60044 39200
rect 60844 37398 60872 39200
rect 61120 37398 61148 39306
rect 61750 39200 61806 40000
rect 62578 39200 62634 40000
rect 63498 39200 63554 40000
rect 64418 39200 64474 40000
rect 65246 39200 65302 40000
rect 66166 39200 66222 40000
rect 66994 39200 67050 40000
rect 67914 39200 67970 40000
rect 68742 39200 68798 40000
rect 69662 39200 69718 40000
rect 70490 39200 70546 40000
rect 71410 39200 71466 40000
rect 72238 39200 72294 40000
rect 73158 39200 73214 40000
rect 73986 39200 74042 40000
rect 74906 39200 74962 40000
rect 75826 39200 75882 40000
rect 76654 39200 76710 40000
rect 77574 39200 77630 40000
rect 78402 39200 78458 40000
rect 79322 39200 79378 40000
rect 80150 39200 80206 40000
rect 81070 39200 81126 40000
rect 81898 39200 81954 40000
rect 82818 39200 82874 40000
rect 83646 39200 83702 40000
rect 84566 39200 84622 40000
rect 85394 39200 85450 40000
rect 86314 39200 86370 40000
rect 87142 39200 87198 40000
rect 88062 39200 88118 40000
rect 88982 39200 89038 40000
rect 89444 39296 89496 39302
rect 89444 39238 89496 39244
rect 61764 37482 61792 39200
rect 61764 37466 61884 37482
rect 61764 37460 61896 37466
rect 61764 37454 61844 37460
rect 61844 37402 61896 37408
rect 60832 37392 60884 37398
rect 60832 37334 60884 37340
rect 61108 37392 61160 37398
rect 61108 37334 61160 37340
rect 61660 37324 61712 37330
rect 61660 37266 61712 37272
rect 60004 36916 60056 36922
rect 60004 36858 60056 36864
rect 60096 36644 60148 36650
rect 60096 36586 60148 36592
rect 59818 36544 59874 36553
rect 59818 36479 59874 36488
rect 59832 36310 59860 36479
rect 59820 36304 59872 36310
rect 59820 36246 59872 36252
rect 59636 34536 59688 34542
rect 59636 34478 59688 34484
rect 59372 34326 59492 34354
rect 59372 33862 59400 34326
rect 59360 33856 59412 33862
rect 59360 33798 59412 33804
rect 59372 33454 59400 33798
rect 59360 33448 59412 33454
rect 59360 33390 59412 33396
rect 59452 33380 59504 33386
rect 59452 33322 59504 33328
rect 59268 32836 59320 32842
rect 59268 32778 59320 32784
rect 58912 31726 59124 31754
rect 58808 31680 58860 31686
rect 58808 31622 58860 31628
rect 58820 30734 58848 31622
rect 58808 30728 58860 30734
rect 58808 30670 58860 30676
rect 58820 22574 58848 30670
rect 59096 30666 59124 31726
rect 59084 30660 59136 30666
rect 59084 30602 59136 30608
rect 58808 22568 58860 22574
rect 58808 22510 58860 22516
rect 58900 21956 58952 21962
rect 58900 21898 58952 21904
rect 58912 21146 58940 21898
rect 58992 21548 59044 21554
rect 58992 21490 59044 21496
rect 59004 21146 59032 21490
rect 58900 21140 58952 21146
rect 58900 21082 58952 21088
rect 58992 21140 59044 21146
rect 58992 21082 59044 21088
rect 58900 20460 58952 20466
rect 58900 20402 58952 20408
rect 58716 17128 58768 17134
rect 58716 17070 58768 17076
rect 58728 16794 58756 17070
rect 58716 16788 58768 16794
rect 58716 16730 58768 16736
rect 58808 15700 58860 15706
rect 58808 15642 58860 15648
rect 58820 15502 58848 15642
rect 58808 15496 58860 15502
rect 58808 15438 58860 15444
rect 58716 14476 58768 14482
rect 58716 14418 58768 14424
rect 58728 14006 58756 14418
rect 58716 14000 58768 14006
rect 58716 13942 58768 13948
rect 58624 12708 58676 12714
rect 58624 12650 58676 12656
rect 58912 12434 58940 20402
rect 59096 16590 59124 30602
rect 59174 27024 59230 27033
rect 59174 26959 59176 26968
rect 59228 26959 59230 26968
rect 59176 26930 59228 26936
rect 59280 26858 59308 32778
rect 59360 30932 59412 30938
rect 59360 30874 59412 30880
rect 59372 30734 59400 30874
rect 59360 30728 59412 30734
rect 59360 30670 59412 30676
rect 59360 27668 59412 27674
rect 59360 27610 59412 27616
rect 59268 26852 59320 26858
rect 59268 26794 59320 26800
rect 59266 26616 59322 26625
rect 59266 26551 59322 26560
rect 59280 26450 59308 26551
rect 59268 26444 59320 26450
rect 59268 26386 59320 26392
rect 59372 22094 59400 27610
rect 59464 26450 59492 33322
rect 59648 30734 59676 34478
rect 59728 33380 59780 33386
rect 59728 33322 59780 33328
rect 59740 32978 59768 33322
rect 59728 32972 59780 32978
rect 59728 32914 59780 32920
rect 59740 32298 59768 32914
rect 59728 32292 59780 32298
rect 59728 32234 59780 32240
rect 59726 31376 59782 31385
rect 59726 31311 59728 31320
rect 59780 31311 59782 31320
rect 59728 31282 59780 31288
rect 59636 30728 59688 30734
rect 59636 30670 59688 30676
rect 59544 30320 59596 30326
rect 59544 30262 59596 30268
rect 59452 26444 59504 26450
rect 59452 26386 59504 26392
rect 59372 22066 59492 22094
rect 59360 21480 59412 21486
rect 59360 21422 59412 21428
rect 59372 19718 59400 21422
rect 59360 19712 59412 19718
rect 59360 19654 59412 19660
rect 59358 19136 59414 19145
rect 59358 19071 59414 19080
rect 59372 18970 59400 19071
rect 59464 18970 59492 22066
rect 59360 18964 59412 18970
rect 59360 18906 59412 18912
rect 59452 18964 59504 18970
rect 59452 18906 59504 18912
rect 59360 18828 59412 18834
rect 59360 18770 59412 18776
rect 59372 18222 59400 18770
rect 59360 18216 59412 18222
rect 59360 18158 59412 18164
rect 59084 16584 59136 16590
rect 59084 16526 59136 16532
rect 59176 16584 59228 16590
rect 59176 16526 59228 16532
rect 58992 16244 59044 16250
rect 58992 16186 59044 16192
rect 59004 15706 59032 16186
rect 59188 16046 59216 16526
rect 59176 16040 59228 16046
rect 59176 15982 59228 15988
rect 59360 16040 59412 16046
rect 59360 15982 59412 15988
rect 58992 15700 59044 15706
rect 58992 15642 59044 15648
rect 59004 15502 59032 15642
rect 58992 15496 59044 15502
rect 58992 15438 59044 15444
rect 59176 15496 59228 15502
rect 59176 15438 59228 15444
rect 58820 12406 58940 12434
rect 58820 12306 58848 12406
rect 58808 12300 58860 12306
rect 58808 12242 58860 12248
rect 58072 12232 58124 12238
rect 58072 12174 58124 12180
rect 58532 12232 58584 12238
rect 58532 12174 58584 12180
rect 58992 12232 59044 12238
rect 58992 12174 59044 12180
rect 58084 11898 58112 12174
rect 57980 11892 58032 11898
rect 57980 11834 58032 11840
rect 58072 11892 58124 11898
rect 58072 11834 58124 11840
rect 57992 10810 58020 11834
rect 58072 11144 58124 11150
rect 58072 11086 58124 11092
rect 57980 10804 58032 10810
rect 57980 10746 58032 10752
rect 58084 8906 58112 11086
rect 58164 10600 58216 10606
rect 58164 10542 58216 10548
rect 58176 10062 58204 10542
rect 58164 10056 58216 10062
rect 58164 9998 58216 10004
rect 58072 8900 58124 8906
rect 58072 8842 58124 8848
rect 58544 5846 58572 12174
rect 59004 11830 59032 12174
rect 58992 11824 59044 11830
rect 58992 11766 59044 11772
rect 58900 7472 58952 7478
rect 58900 7414 58952 7420
rect 58532 5840 58584 5846
rect 58532 5782 58584 5788
rect 57888 5296 57940 5302
rect 57888 5238 57940 5244
rect 57336 4684 57388 4690
rect 57336 4626 57388 4632
rect 57152 3596 57204 3602
rect 57152 3538 57204 3544
rect 56876 3392 56928 3398
rect 56876 3334 56928 3340
rect 57164 2496 57192 3538
rect 57348 2650 57376 4626
rect 58256 4548 58308 4554
rect 58256 4490 58308 4496
rect 57428 4072 57480 4078
rect 57428 4014 57480 4020
rect 57336 2644 57388 2650
rect 57336 2586 57388 2592
rect 56980 2468 57192 2496
rect 56980 800 57008 2468
rect 57152 2372 57204 2378
rect 57152 2314 57204 2320
rect 57164 800 57192 2314
rect 57440 800 57468 4014
rect 58164 3596 58216 3602
rect 58164 3538 58216 3544
rect 57980 3528 58032 3534
rect 57980 3470 58032 3476
rect 57612 2984 57664 2990
rect 57612 2926 57664 2932
rect 57624 800 57652 2926
rect 57796 2916 57848 2922
rect 57796 2858 57848 2864
rect 57808 800 57836 2858
rect 57992 800 58020 3470
rect 58072 2508 58124 2514
rect 58072 2450 58124 2456
rect 58084 2310 58112 2450
rect 58072 2304 58124 2310
rect 58072 2246 58124 2252
rect 58084 1358 58112 2246
rect 58072 1352 58124 1358
rect 58072 1294 58124 1300
rect 58176 800 58204 3538
rect 58268 1086 58296 4490
rect 58348 3052 58400 3058
rect 58348 2994 58400 3000
rect 58360 2582 58388 2994
rect 58544 2774 58572 5782
rect 58912 5166 58940 7414
rect 59004 5778 59032 11766
rect 58992 5772 59044 5778
rect 58992 5714 59044 5720
rect 59084 5228 59136 5234
rect 59084 5170 59136 5176
rect 58900 5160 58952 5166
rect 59096 5137 59124 5170
rect 58900 5102 58952 5108
rect 59082 5128 59138 5137
rect 59082 5063 59138 5072
rect 58624 4072 58676 4078
rect 58624 4014 58676 4020
rect 58452 2746 58572 2774
rect 58348 2576 58400 2582
rect 58348 2518 58400 2524
rect 58452 1986 58480 2746
rect 58360 1958 58480 1986
rect 58360 1154 58388 1958
rect 58440 1488 58492 1494
rect 58440 1430 58492 1436
rect 58348 1148 58400 1154
rect 58348 1090 58400 1096
rect 58256 1080 58308 1086
rect 58256 1022 58308 1028
rect 58452 800 58480 1430
rect 58636 800 58664 4014
rect 59084 4004 59136 4010
rect 59084 3946 59136 3952
rect 58808 3596 58860 3602
rect 58808 3538 58860 3544
rect 58820 800 58848 3538
rect 58992 2848 59044 2854
rect 58992 2790 59044 2796
rect 59004 800 59032 2790
rect 59096 1442 59124 3946
rect 59188 2582 59216 15438
rect 59268 14952 59320 14958
rect 59268 14894 59320 14900
rect 59280 12306 59308 14894
rect 59268 12300 59320 12306
rect 59268 12242 59320 12248
rect 59268 12164 59320 12170
rect 59268 12106 59320 12112
rect 59280 11898 59308 12106
rect 59268 11892 59320 11898
rect 59268 11834 59320 11840
rect 59268 9104 59320 9110
rect 59268 9046 59320 9052
rect 59280 8673 59308 9046
rect 59266 8664 59322 8673
rect 59266 8599 59322 8608
rect 59268 5092 59320 5098
rect 59268 5034 59320 5040
rect 59176 2576 59228 2582
rect 59176 2518 59228 2524
rect 59096 1414 59216 1442
rect 59188 800 59216 1414
rect 59280 882 59308 5034
rect 59372 2990 59400 15982
rect 59464 14958 59492 18906
rect 59452 14952 59504 14958
rect 59452 14894 59504 14900
rect 59556 12442 59584 30262
rect 59648 28966 59676 30670
rect 59636 28960 59688 28966
rect 59636 28902 59688 28908
rect 59728 28960 59780 28966
rect 59728 28902 59780 28908
rect 59740 28490 59768 28902
rect 59728 28484 59780 28490
rect 59728 28426 59780 28432
rect 59832 27146 59860 36246
rect 60004 31680 60056 31686
rect 60004 31622 60056 31628
rect 60016 31278 60044 31622
rect 60004 31272 60056 31278
rect 60004 31214 60056 31220
rect 60016 31142 60044 31214
rect 60004 31136 60056 31142
rect 60004 31078 60056 31084
rect 59912 30932 59964 30938
rect 59912 30874 59964 30880
rect 59924 29866 59952 30874
rect 60016 30802 60044 31078
rect 60004 30796 60056 30802
rect 60004 30738 60056 30744
rect 60016 30054 60044 30738
rect 60004 30048 60056 30054
rect 60004 29990 60056 29996
rect 59924 29838 60044 29866
rect 59740 27118 59860 27146
rect 59740 22094 59768 27118
rect 59912 26920 59964 26926
rect 59912 26862 59964 26868
rect 59648 22066 59768 22094
rect 59648 14482 59676 22066
rect 59728 20460 59780 20466
rect 59728 20402 59780 20408
rect 59740 19990 59768 20402
rect 59728 19984 59780 19990
rect 59728 19926 59780 19932
rect 59728 18828 59780 18834
rect 59728 18770 59780 18776
rect 59820 18828 59872 18834
rect 59820 18770 59872 18776
rect 59740 17746 59768 18770
rect 59832 18630 59860 18770
rect 59820 18624 59872 18630
rect 59820 18566 59872 18572
rect 59728 17740 59780 17746
rect 59728 17682 59780 17688
rect 59636 14476 59688 14482
rect 59636 14418 59688 14424
rect 59728 14476 59780 14482
rect 59728 14418 59780 14424
rect 59544 12436 59596 12442
rect 59544 12378 59596 12384
rect 59740 11150 59768 14418
rect 59728 11144 59780 11150
rect 59728 11086 59780 11092
rect 59452 9104 59504 9110
rect 59452 9046 59504 9052
rect 59464 5710 59492 9046
rect 59452 5704 59504 5710
rect 59452 5646 59504 5652
rect 59360 2984 59412 2990
rect 59360 2926 59412 2932
rect 59452 2984 59504 2990
rect 59452 2926 59504 2932
rect 59268 876 59320 882
rect 59268 818 59320 824
rect 59464 800 59492 2926
rect 59636 2304 59688 2310
rect 59636 2246 59688 2252
rect 59648 800 59676 2246
rect 59740 1358 59768 11086
rect 59924 7206 59952 26862
rect 60016 25226 60044 29838
rect 60004 25220 60056 25226
rect 60004 25162 60056 25168
rect 60108 16726 60136 36586
rect 61198 35048 61254 35057
rect 61198 34983 61254 34992
rect 60370 33688 60426 33697
rect 60370 33623 60426 33632
rect 60384 33522 60412 33623
rect 60372 33516 60424 33522
rect 60372 33458 60424 33464
rect 60280 33448 60332 33454
rect 60280 33390 60332 33396
rect 60740 33448 60792 33454
rect 60924 33448 60976 33454
rect 60792 33408 60872 33436
rect 60740 33390 60792 33396
rect 60292 31686 60320 33390
rect 60372 33380 60424 33386
rect 60372 33322 60424 33328
rect 60384 33289 60412 33322
rect 60740 33312 60792 33318
rect 60370 33280 60426 33289
rect 60370 33215 60426 33224
rect 60738 33280 60740 33289
rect 60792 33280 60794 33289
rect 60738 33215 60794 33224
rect 60280 31680 60332 31686
rect 60280 31622 60332 31628
rect 60280 31340 60332 31346
rect 60280 31282 60332 31288
rect 60188 31136 60240 31142
rect 60188 31078 60240 31084
rect 60200 26246 60228 31078
rect 60292 30938 60320 31282
rect 60280 30932 60332 30938
rect 60280 30874 60332 30880
rect 60384 28694 60412 33215
rect 60556 31680 60608 31686
rect 60556 31622 60608 31628
rect 60568 30734 60596 31622
rect 60646 31376 60702 31385
rect 60646 31311 60648 31320
rect 60700 31311 60702 31320
rect 60648 31282 60700 31288
rect 60740 31272 60792 31278
rect 60740 31214 60792 31220
rect 60556 30728 60608 30734
rect 60556 30670 60608 30676
rect 60372 28688 60424 28694
rect 60372 28630 60424 28636
rect 60464 27464 60516 27470
rect 60464 27406 60516 27412
rect 60280 26444 60332 26450
rect 60280 26386 60332 26392
rect 60372 26444 60424 26450
rect 60372 26386 60424 26392
rect 60188 26240 60240 26246
rect 60188 26182 60240 26188
rect 60188 25220 60240 25226
rect 60188 25162 60240 25168
rect 60096 16720 60148 16726
rect 60096 16662 60148 16668
rect 60200 14482 60228 25162
rect 60292 14618 60320 26386
rect 60384 26314 60412 26386
rect 60476 26314 60504 27406
rect 60648 27328 60700 27334
rect 60648 27270 60700 27276
rect 60660 27130 60688 27270
rect 60648 27124 60700 27130
rect 60648 27066 60700 27072
rect 60646 26616 60702 26625
rect 60646 26551 60702 26560
rect 60660 26518 60688 26551
rect 60556 26512 60608 26518
rect 60554 26480 60556 26489
rect 60648 26512 60700 26518
rect 60608 26480 60610 26489
rect 60648 26454 60700 26460
rect 60554 26415 60610 26424
rect 60372 26308 60424 26314
rect 60372 26250 60424 26256
rect 60464 26308 60516 26314
rect 60464 26250 60516 26256
rect 60752 25498 60780 31214
rect 60844 26330 60872 33408
rect 60924 33390 60976 33396
rect 60936 32910 60964 33390
rect 61108 33312 61160 33318
rect 61108 33254 61160 33260
rect 60924 32904 60976 32910
rect 60924 32846 60976 32852
rect 61016 32020 61068 32026
rect 61016 31962 61068 31968
rect 61028 29578 61056 31962
rect 61120 30870 61148 33254
rect 61108 30864 61160 30870
rect 61108 30806 61160 30812
rect 61016 29572 61068 29578
rect 61016 29514 61068 29520
rect 60924 27328 60976 27334
rect 60924 27270 60976 27276
rect 60936 27033 60964 27270
rect 60922 27024 60978 27033
rect 61212 26994 61240 34983
rect 61672 33998 61700 37266
rect 62592 36922 62620 39200
rect 63512 37398 63540 39200
rect 64432 37754 64460 39200
rect 64432 37726 64552 37754
rect 63776 37664 63828 37670
rect 63776 37606 63828 37612
rect 63788 37398 63816 37606
rect 64524 37466 64552 37726
rect 64880 37664 64932 37670
rect 64880 37606 64932 37612
rect 64512 37460 64564 37466
rect 64512 37402 64564 37408
rect 63500 37392 63552 37398
rect 63500 37334 63552 37340
rect 63776 37392 63828 37398
rect 63776 37334 63828 37340
rect 64328 37324 64380 37330
rect 64328 37266 64380 37272
rect 62580 36916 62632 36922
rect 62580 36858 62632 36864
rect 62672 36644 62724 36650
rect 62672 36586 62724 36592
rect 61844 35624 61896 35630
rect 61844 35566 61896 35572
rect 61856 35154 61884 35566
rect 62026 35184 62082 35193
rect 61844 35148 61896 35154
rect 62026 35119 62028 35128
rect 61844 35090 61896 35096
rect 62080 35119 62082 35128
rect 62580 35148 62632 35154
rect 62028 35090 62080 35096
rect 62580 35090 62632 35096
rect 62212 35080 62264 35086
rect 61856 35028 62212 35034
rect 62592 35057 62620 35090
rect 61856 35022 62264 35028
rect 62578 35048 62634 35057
rect 61856 35006 62252 35022
rect 61856 34950 61884 35006
rect 62578 34983 62634 34992
rect 61844 34944 61896 34950
rect 61844 34886 61896 34892
rect 61660 33992 61712 33998
rect 61660 33934 61712 33940
rect 61290 33688 61346 33697
rect 61290 33623 61346 33632
rect 61304 33454 61332 33623
rect 61384 33516 61436 33522
rect 61384 33458 61436 33464
rect 61292 33448 61344 33454
rect 61292 33390 61344 33396
rect 61396 29782 61424 33458
rect 61476 33380 61528 33386
rect 61476 33322 61528 33328
rect 61488 33289 61516 33322
rect 61474 33280 61530 33289
rect 61474 33215 61530 33224
rect 61856 32774 61884 34886
rect 62028 33992 62080 33998
rect 62028 33934 62080 33940
rect 62040 33522 62068 33934
rect 62684 33833 62712 36586
rect 63040 36576 63092 36582
rect 63040 36518 63092 36524
rect 63052 36106 63080 36518
rect 63132 36168 63184 36174
rect 63132 36110 63184 36116
rect 63408 36168 63460 36174
rect 63408 36110 63460 36116
rect 63040 36100 63092 36106
rect 63040 36042 63092 36048
rect 63144 35193 63172 36110
rect 63130 35184 63186 35193
rect 63130 35119 63186 35128
rect 62670 33824 62726 33833
rect 62670 33759 62726 33768
rect 62028 33516 62080 33522
rect 62028 33458 62080 33464
rect 61844 32768 61896 32774
rect 61844 32710 61896 32716
rect 62028 31272 62080 31278
rect 62028 31214 62080 31220
rect 62040 30054 62068 31214
rect 62488 30592 62540 30598
rect 62488 30534 62540 30540
rect 62028 30048 62080 30054
rect 62028 29990 62080 29996
rect 61384 29776 61436 29782
rect 61384 29718 61436 29724
rect 62028 29776 62080 29782
rect 62028 29718 62080 29724
rect 61936 28620 61988 28626
rect 61936 28562 61988 28568
rect 61844 28552 61896 28558
rect 61844 28494 61896 28500
rect 61856 27674 61884 28494
rect 61844 27668 61896 27674
rect 61844 27610 61896 27616
rect 60922 26959 60978 26968
rect 61200 26988 61252 26994
rect 61200 26930 61252 26936
rect 61212 26489 61240 26930
rect 61198 26480 61254 26489
rect 61198 26415 61254 26424
rect 60844 26302 61792 26330
rect 60740 25492 60792 25498
rect 60740 25434 60792 25440
rect 60844 21962 60872 26302
rect 61292 26240 61344 26246
rect 61292 26182 61344 26188
rect 61200 25832 61252 25838
rect 61200 25774 61252 25780
rect 61212 24070 61240 25774
rect 61304 25362 61332 26182
rect 61764 25838 61792 26302
rect 61660 25832 61712 25838
rect 61660 25774 61712 25780
rect 61752 25832 61804 25838
rect 61752 25774 61804 25780
rect 61384 25492 61436 25498
rect 61384 25434 61436 25440
rect 61396 25362 61424 25434
rect 61292 25356 61344 25362
rect 61292 25298 61344 25304
rect 61384 25356 61436 25362
rect 61384 25298 61436 25304
rect 61200 24064 61252 24070
rect 61200 24006 61252 24012
rect 61384 23588 61436 23594
rect 61384 23530 61436 23536
rect 61016 23112 61068 23118
rect 61016 23054 61068 23060
rect 61028 22545 61056 23054
rect 61014 22536 61070 22545
rect 61014 22471 61070 22480
rect 60832 21956 60884 21962
rect 60832 21898 60884 21904
rect 60830 21720 60886 21729
rect 60830 21655 60886 21664
rect 60844 21622 60872 21655
rect 61028 21622 61056 22471
rect 61106 21720 61162 21729
rect 61106 21655 61162 21664
rect 61120 21622 61148 21655
rect 60832 21616 60884 21622
rect 60832 21558 60884 21564
rect 61016 21616 61068 21622
rect 61016 21558 61068 21564
rect 61108 21616 61160 21622
rect 61108 21558 61160 21564
rect 60464 21480 60516 21486
rect 60464 21422 60516 21428
rect 60832 21480 60884 21486
rect 60884 21440 61056 21468
rect 60832 21422 60884 21428
rect 60372 19304 60424 19310
rect 60372 19246 60424 19252
rect 60280 14612 60332 14618
rect 60280 14554 60332 14560
rect 60188 14476 60240 14482
rect 60188 14418 60240 14424
rect 60200 7546 60228 14418
rect 60278 14376 60334 14385
rect 60278 14311 60280 14320
rect 60332 14311 60334 14320
rect 60280 14282 60332 14288
rect 60384 11354 60412 19246
rect 60476 18714 60504 21422
rect 60554 20904 60610 20913
rect 60554 20839 60556 20848
rect 60608 20839 60610 20848
rect 60556 20810 60608 20816
rect 60924 19712 60976 19718
rect 60924 19654 60976 19660
rect 60738 19544 60794 19553
rect 60738 19479 60794 19488
rect 60752 19378 60780 19479
rect 60740 19372 60792 19378
rect 60740 19314 60792 19320
rect 60832 19372 60884 19378
rect 60832 19314 60884 19320
rect 60738 19272 60794 19281
rect 60648 19236 60700 19242
rect 60738 19207 60794 19216
rect 60648 19178 60700 19184
rect 60476 18686 60596 18714
rect 60462 18320 60518 18329
rect 60462 18255 60518 18264
rect 60476 18086 60504 18255
rect 60568 18222 60596 18686
rect 60660 18601 60688 19178
rect 60752 19174 60780 19207
rect 60740 19168 60792 19174
rect 60844 19145 60872 19314
rect 60740 19110 60792 19116
rect 60830 19136 60886 19145
rect 60830 19071 60886 19080
rect 60832 18896 60884 18902
rect 60832 18838 60884 18844
rect 60844 18698 60872 18838
rect 60936 18698 60964 19654
rect 60832 18692 60884 18698
rect 60832 18634 60884 18640
rect 60924 18692 60976 18698
rect 60924 18634 60976 18640
rect 60646 18592 60702 18601
rect 60646 18527 60702 18536
rect 60556 18216 60608 18222
rect 60556 18158 60608 18164
rect 60464 18080 60516 18086
rect 60464 18022 60516 18028
rect 60464 14952 60516 14958
rect 60464 14894 60516 14900
rect 60476 14346 60504 14894
rect 60464 14340 60516 14346
rect 60464 14282 60516 14288
rect 60464 12912 60516 12918
rect 60464 12854 60516 12860
rect 60372 11348 60424 11354
rect 60372 11290 60424 11296
rect 60188 7540 60240 7546
rect 60188 7482 60240 7488
rect 59912 7200 59964 7206
rect 59912 7142 59964 7148
rect 59820 4004 59872 4010
rect 59820 3946 59872 3952
rect 59728 1352 59780 1358
rect 59728 1294 59780 1300
rect 59832 800 59860 3946
rect 60096 2984 60148 2990
rect 60096 2926 60148 2932
rect 60108 2774 60136 2926
rect 60280 2916 60332 2922
rect 60280 2858 60332 2864
rect 60016 2746 60136 2774
rect 60016 800 60044 2746
rect 60292 2650 60320 2858
rect 60280 2644 60332 2650
rect 60280 2586 60332 2592
rect 60476 2582 60504 12854
rect 60568 12714 60596 18158
rect 61028 14521 61056 21440
rect 61290 21448 61346 21457
rect 61290 21383 61346 21392
rect 61304 21350 61332 21383
rect 61292 21344 61344 21350
rect 61292 21286 61344 21292
rect 61108 19712 61160 19718
rect 61108 19654 61160 19660
rect 61120 19553 61148 19654
rect 61106 19544 61162 19553
rect 61106 19479 61162 19488
rect 61108 19304 61160 19310
rect 61106 19272 61108 19281
rect 61160 19272 61162 19281
rect 61106 19207 61162 19216
rect 61292 17536 61344 17542
rect 61292 17478 61344 17484
rect 61304 16726 61332 17478
rect 61292 16720 61344 16726
rect 61292 16662 61344 16668
rect 61292 14952 61344 14958
rect 61292 14894 61344 14900
rect 61014 14512 61070 14521
rect 60740 14476 60792 14482
rect 61014 14447 61070 14456
rect 60740 14418 60792 14424
rect 60752 14278 60780 14418
rect 60740 14272 60792 14278
rect 60740 14214 60792 14220
rect 60832 14272 60884 14278
rect 60832 14214 60884 14220
rect 60844 14006 60872 14214
rect 60832 14000 60884 14006
rect 60832 13942 60884 13948
rect 60556 12708 60608 12714
rect 60556 12650 60608 12656
rect 60830 8664 60886 8673
rect 60740 8628 60792 8634
rect 60830 8599 60832 8608
rect 60740 8570 60792 8576
rect 60884 8599 60886 8608
rect 60832 8570 60884 8576
rect 60752 8537 60780 8570
rect 60738 8528 60794 8537
rect 60738 8463 60794 8472
rect 60832 8424 60884 8430
rect 60832 8366 60884 8372
rect 60740 4072 60792 4078
rect 60568 4032 60740 4060
rect 60464 2576 60516 2582
rect 60464 2518 60516 2524
rect 60372 2372 60424 2378
rect 60372 2314 60424 2320
rect 60384 1494 60412 2314
rect 60568 2088 60596 4032
rect 60740 4014 60792 4020
rect 60648 3596 60700 3602
rect 60648 3538 60700 3544
rect 60476 2060 60596 2088
rect 60372 1488 60424 1494
rect 60372 1430 60424 1436
rect 60188 1420 60240 1426
rect 60188 1362 60240 1368
rect 60200 800 60228 1362
rect 60476 800 60504 2060
rect 60660 800 60688 3538
rect 60844 3058 60872 8366
rect 61028 4622 61056 14447
rect 61106 14376 61162 14385
rect 61106 14311 61108 14320
rect 61160 14311 61162 14320
rect 61108 14282 61160 14288
rect 61304 7562 61332 14894
rect 61396 7698 61424 23530
rect 61474 23080 61530 23089
rect 61474 23015 61530 23024
rect 61488 11014 61516 23015
rect 61568 21480 61620 21486
rect 61566 21448 61568 21457
rect 61620 21448 61622 21457
rect 61566 21383 61622 21392
rect 61566 21312 61622 21321
rect 61566 21247 61622 21256
rect 61580 12102 61608 21247
rect 61568 12096 61620 12102
rect 61568 12038 61620 12044
rect 61476 11008 61528 11014
rect 61476 10950 61528 10956
rect 61568 11008 61620 11014
rect 61568 10950 61620 10956
rect 61580 10690 61608 10950
rect 61672 10742 61700 25774
rect 61752 23588 61804 23594
rect 61752 23530 61804 23536
rect 61764 19922 61792 23530
rect 61948 22094 61976 28562
rect 62040 25265 62068 29718
rect 62026 25256 62082 25265
rect 62026 25191 62082 25200
rect 62500 23186 62528 30534
rect 62684 28626 62712 33759
rect 62856 32428 62908 32434
rect 62856 32370 62908 32376
rect 62764 30184 62816 30190
rect 62762 30152 62764 30161
rect 62816 30152 62818 30161
rect 62762 30087 62818 30096
rect 62672 28620 62724 28626
rect 62672 28562 62724 28568
rect 62120 23180 62172 23186
rect 62120 23122 62172 23128
rect 62488 23180 62540 23186
rect 62488 23122 62540 23128
rect 61948 22066 62068 22094
rect 61844 21548 61896 21554
rect 61844 21490 61896 21496
rect 61856 21078 61884 21490
rect 61844 21072 61896 21078
rect 61844 21014 61896 21020
rect 61752 19916 61804 19922
rect 61752 19858 61804 19864
rect 61936 19440 61988 19446
rect 61936 19382 61988 19388
rect 61948 18630 61976 19382
rect 61936 18624 61988 18630
rect 61936 18566 61988 18572
rect 61844 16720 61896 16726
rect 61844 16662 61896 16668
rect 61856 12714 61884 16662
rect 61752 12708 61804 12714
rect 61752 12650 61804 12656
rect 61844 12708 61896 12714
rect 61844 12650 61896 12656
rect 61488 10674 61608 10690
rect 61660 10736 61712 10742
rect 61660 10678 61712 10684
rect 61476 10668 61608 10674
rect 61528 10662 61608 10668
rect 61476 10610 61528 10616
rect 61660 10600 61712 10606
rect 61660 10542 61712 10548
rect 61672 9602 61700 10542
rect 61764 9738 61792 12650
rect 61856 10606 61884 12650
rect 62040 12434 62068 22066
rect 62132 18970 62160 23122
rect 62212 23112 62264 23118
rect 62212 23054 62264 23060
rect 62224 22545 62252 23054
rect 62210 22536 62266 22545
rect 62210 22471 62266 22480
rect 62120 18964 62172 18970
rect 62120 18906 62172 18912
rect 62396 18964 62448 18970
rect 62396 18906 62448 18912
rect 62210 18728 62266 18737
rect 62210 18663 62266 18672
rect 62120 15088 62172 15094
rect 62120 15030 62172 15036
rect 62132 14890 62160 15030
rect 62120 14884 62172 14890
rect 62120 14826 62172 14832
rect 62120 13728 62172 13734
rect 62120 13670 62172 13676
rect 61948 12406 62068 12434
rect 61844 10600 61896 10606
rect 61844 10542 61896 10548
rect 61764 9710 61884 9738
rect 61672 9574 61792 9602
rect 61658 8936 61714 8945
rect 61764 8906 61792 9574
rect 61658 8871 61660 8880
rect 61712 8871 61714 8880
rect 61752 8900 61804 8906
rect 61660 8842 61712 8848
rect 61752 8842 61804 8848
rect 61658 8664 61714 8673
rect 61658 8599 61714 8608
rect 61672 8430 61700 8599
rect 61660 8424 61712 8430
rect 61660 8366 61712 8372
rect 61396 7670 61516 7698
rect 61304 7534 61424 7562
rect 61016 4616 61068 4622
rect 61016 4558 61068 4564
rect 60924 4140 60976 4146
rect 60924 4082 60976 4088
rect 61016 4140 61068 4146
rect 61016 4082 61068 4088
rect 60936 4010 60964 4082
rect 60924 4004 60976 4010
rect 60924 3946 60976 3952
rect 60832 3052 60884 3058
rect 60832 2994 60884 3000
rect 60924 2984 60976 2990
rect 60924 2926 60976 2932
rect 60740 2576 60792 2582
rect 60936 2564 60964 2926
rect 60740 2518 60792 2524
rect 60844 2536 60964 2564
rect 60752 2310 60780 2518
rect 60740 2304 60792 2310
rect 60740 2246 60792 2252
rect 60844 800 60872 2536
rect 61028 800 61056 4082
rect 61292 3596 61344 3602
rect 61292 3538 61344 3544
rect 61200 2508 61252 2514
rect 61200 2450 61252 2456
rect 61212 2106 61240 2450
rect 61200 2100 61252 2106
rect 61200 2042 61252 2048
rect 61304 800 61332 3538
rect 61396 2650 61424 7534
rect 61488 5574 61516 7670
rect 61568 7404 61620 7410
rect 61568 7346 61620 7352
rect 61476 5568 61528 5574
rect 61476 5510 61528 5516
rect 61580 2922 61608 7346
rect 61764 6798 61792 8842
rect 61856 8362 61884 9710
rect 61844 8356 61896 8362
rect 61844 8298 61896 8304
rect 61844 7336 61896 7342
rect 61844 7278 61896 7284
rect 61752 6792 61804 6798
rect 61752 6734 61804 6740
rect 61764 6118 61792 6734
rect 61752 6112 61804 6118
rect 61752 6054 61804 6060
rect 61764 4593 61792 6054
rect 61856 4690 61884 7278
rect 61844 4684 61896 4690
rect 61844 4626 61896 4632
rect 61750 4584 61806 4593
rect 61750 4519 61806 4528
rect 61948 3890 61976 12406
rect 62132 10470 62160 13670
rect 62120 10464 62172 10470
rect 62120 10406 62172 10412
rect 62224 9674 62252 18663
rect 62408 18290 62436 18906
rect 62396 18284 62448 18290
rect 62396 18226 62448 18232
rect 62396 16244 62448 16250
rect 62396 16186 62448 16192
rect 62408 15502 62436 16186
rect 62396 15496 62448 15502
rect 62396 15438 62448 15444
rect 62304 15156 62356 15162
rect 62304 15098 62356 15104
rect 62132 9646 62252 9674
rect 62028 8968 62080 8974
rect 62028 8910 62080 8916
rect 62040 6390 62068 8910
rect 62028 6384 62080 6390
rect 62028 6326 62080 6332
rect 62028 4752 62080 4758
rect 62026 4720 62028 4729
rect 62080 4720 62082 4729
rect 62026 4655 62082 4664
rect 62132 4554 62160 9646
rect 62210 8528 62266 8537
rect 62210 8463 62266 8472
rect 62224 8430 62252 8463
rect 62212 8424 62264 8430
rect 62212 8366 62264 8372
rect 62316 4690 62344 15098
rect 62396 15020 62448 15026
rect 62396 14962 62448 14968
rect 62408 14929 62436 14962
rect 62394 14920 62450 14929
rect 62394 14855 62450 14864
rect 62500 9518 62528 23122
rect 62580 23112 62632 23118
rect 62580 23054 62632 23060
rect 62592 21418 62620 23054
rect 62868 23050 62896 32370
rect 63144 28966 63172 35119
rect 63224 33856 63276 33862
rect 63224 33798 63276 33804
rect 63316 33856 63368 33862
rect 63316 33798 63368 33804
rect 63236 33318 63264 33798
rect 63224 33312 63276 33318
rect 63224 33254 63276 33260
rect 63224 30728 63276 30734
rect 63224 30670 63276 30676
rect 63236 30598 63264 30670
rect 63224 30592 63276 30598
rect 63224 30534 63276 30540
rect 63040 28960 63092 28966
rect 63040 28902 63092 28908
rect 63132 28960 63184 28966
rect 63132 28902 63184 28908
rect 63052 28150 63080 28902
rect 63144 28422 63172 28902
rect 63132 28416 63184 28422
rect 63132 28358 63184 28364
rect 63224 28416 63276 28422
rect 63224 28358 63276 28364
rect 62948 28144 63000 28150
rect 62948 28086 63000 28092
rect 63040 28144 63092 28150
rect 63040 28086 63092 28092
rect 62960 27962 62988 28086
rect 63236 27962 63264 28358
rect 62960 27934 63264 27962
rect 63040 26852 63092 26858
rect 63040 26794 63092 26800
rect 62856 23044 62908 23050
rect 62856 22986 62908 22992
rect 62764 22976 62816 22982
rect 62764 22918 62816 22924
rect 62672 22568 62724 22574
rect 62672 22510 62724 22516
rect 62684 21962 62712 22510
rect 62672 21956 62724 21962
rect 62672 21898 62724 21904
rect 62672 21684 62724 21690
rect 62672 21626 62724 21632
rect 62684 21418 62712 21626
rect 62776 21434 62804 22918
rect 63052 22420 63080 26794
rect 63132 25424 63184 25430
rect 63132 25366 63184 25372
rect 63144 22574 63172 25366
rect 63224 24064 63276 24070
rect 63224 24006 63276 24012
rect 63132 22568 63184 22574
rect 63132 22510 63184 22516
rect 63052 22392 63172 22420
rect 62580 21412 62632 21418
rect 62580 21354 62632 21360
rect 62672 21412 62724 21418
rect 62776 21406 63080 21434
rect 62672 21354 62724 21360
rect 62592 18290 62620 21354
rect 62948 21344 63000 21350
rect 62948 21286 63000 21292
rect 62856 20800 62908 20806
rect 62856 20742 62908 20748
rect 62764 20460 62816 20466
rect 62764 20402 62816 20408
rect 62580 18284 62632 18290
rect 62580 18226 62632 18232
rect 62672 18216 62724 18222
rect 62672 18158 62724 18164
rect 62684 16182 62712 18158
rect 62672 16176 62724 16182
rect 62672 16118 62724 16124
rect 62670 15600 62726 15609
rect 62670 15535 62726 15544
rect 62684 15434 62712 15535
rect 62672 15428 62724 15434
rect 62672 15370 62724 15376
rect 62776 15094 62804 20402
rect 62764 15088 62816 15094
rect 62764 15030 62816 15036
rect 62580 13456 62632 13462
rect 62580 13398 62632 13404
rect 62396 9512 62448 9518
rect 62394 9480 62396 9489
rect 62488 9512 62540 9518
rect 62448 9480 62450 9489
rect 62488 9454 62540 9460
rect 62394 9415 62450 9424
rect 62396 4752 62448 4758
rect 62396 4694 62448 4700
rect 62304 4684 62356 4690
rect 62304 4626 62356 4632
rect 62120 4548 62172 4554
rect 62120 4490 62172 4496
rect 62028 4480 62080 4486
rect 62026 4448 62028 4457
rect 62304 4480 62356 4486
rect 62080 4448 62082 4457
rect 62304 4422 62356 4428
rect 62026 4383 62082 4392
rect 62316 4298 62344 4422
rect 62224 4270 62344 4298
rect 62028 4072 62080 4078
rect 62028 4014 62080 4020
rect 61764 3862 61976 3890
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 61568 2916 61620 2922
rect 61568 2858 61620 2864
rect 61476 2848 61528 2854
rect 61476 2790 61528 2796
rect 61384 2644 61436 2650
rect 61384 2586 61436 2592
rect 61396 2514 61424 2586
rect 61384 2508 61436 2514
rect 61384 2450 61436 2456
rect 61488 800 61516 2790
rect 61672 800 61700 3334
rect 61764 2106 61792 3862
rect 61844 3528 61896 3534
rect 61844 3470 61896 3476
rect 61752 2100 61804 2106
rect 61752 2042 61804 2048
rect 61856 800 61884 3470
rect 62040 3398 62068 4014
rect 62028 3392 62080 3398
rect 62028 3334 62080 3340
rect 62120 2984 62172 2990
rect 62120 2926 62172 2932
rect 62132 2650 62160 2926
rect 62120 2644 62172 2650
rect 62120 2586 62172 2592
rect 62028 2304 62080 2310
rect 62028 2246 62080 2252
rect 62040 1426 62068 2246
rect 62120 2100 62172 2106
rect 62120 2042 62172 2048
rect 62028 1420 62080 1426
rect 62028 1362 62080 1368
rect 62132 1306 62160 2042
rect 62040 1278 62160 1306
rect 62040 800 62068 1278
rect 55494 776 55550 785
rect 55494 711 55550 720
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62026 0 62082 800
rect 62224 746 62252 4270
rect 62304 4140 62356 4146
rect 62304 4082 62356 4088
rect 62316 800 62344 4082
rect 62408 1358 62436 4694
rect 62592 4690 62620 13398
rect 62672 12232 62724 12238
rect 62672 12174 62724 12180
rect 62684 11898 62712 12174
rect 62672 11892 62724 11898
rect 62672 11834 62724 11840
rect 62684 11694 62712 11834
rect 62672 11688 62724 11694
rect 62672 11630 62724 11636
rect 62868 11014 62896 20742
rect 62960 20641 62988 21286
rect 62946 20632 63002 20641
rect 62946 20567 63002 20576
rect 62948 19848 63000 19854
rect 62948 19790 63000 19796
rect 62960 15570 62988 19790
rect 62948 15564 63000 15570
rect 62948 15506 63000 15512
rect 62948 11212 63000 11218
rect 62948 11154 63000 11160
rect 62960 11121 62988 11154
rect 62946 11112 63002 11121
rect 62946 11047 63002 11056
rect 62856 11008 62908 11014
rect 62856 10950 62908 10956
rect 62948 10464 63000 10470
rect 62948 10406 63000 10412
rect 62672 10124 62724 10130
rect 62672 10066 62724 10072
rect 62684 9722 62712 10066
rect 62672 9716 62724 9722
rect 62672 9658 62724 9664
rect 62856 9444 62908 9450
rect 62856 9386 62908 9392
rect 62868 9110 62896 9386
rect 62856 9104 62908 9110
rect 62856 9046 62908 9052
rect 62960 7478 62988 10406
rect 63052 9042 63080 21406
rect 63040 9036 63092 9042
rect 63040 8978 63092 8984
rect 62948 7472 63000 7478
rect 62948 7414 63000 7420
rect 62764 5568 62816 5574
rect 62764 5510 62816 5516
rect 62580 4684 62632 4690
rect 62580 4626 62632 4632
rect 62488 3664 62540 3670
rect 62488 3606 62540 3612
rect 62396 1352 62448 1358
rect 62396 1294 62448 1300
rect 62212 740 62264 746
rect 62212 682 62264 688
rect 62302 0 62358 800
rect 62408 270 62436 1294
rect 62500 800 62528 3606
rect 62776 2990 62804 5510
rect 62854 4584 62910 4593
rect 62854 4519 62856 4528
rect 62908 4519 62910 4528
rect 62856 4490 62908 4496
rect 63040 3528 63092 3534
rect 63040 3470 63092 3476
rect 62856 3392 62908 3398
rect 62856 3334 62908 3340
rect 62764 2984 62816 2990
rect 62764 2926 62816 2932
rect 62672 2848 62724 2854
rect 62672 2790 62724 2796
rect 62684 800 62712 2790
rect 62868 800 62896 3334
rect 63052 800 63080 3470
rect 63144 2582 63172 22392
rect 63236 21010 63264 24006
rect 63224 21004 63276 21010
rect 63224 20946 63276 20952
rect 63236 19854 63264 20946
rect 63224 19848 63276 19854
rect 63224 19790 63276 19796
rect 63224 19236 63276 19242
rect 63224 19178 63276 19184
rect 63236 18154 63264 19178
rect 63224 18148 63276 18154
rect 63224 18090 63276 18096
rect 63236 16114 63264 18090
rect 63224 16108 63276 16114
rect 63224 16050 63276 16056
rect 63328 12434 63356 33798
rect 63420 24682 63448 36110
rect 63500 34944 63552 34950
rect 63500 34886 63552 34892
rect 64236 34944 64288 34950
rect 64236 34886 64288 34892
rect 63512 26246 63540 34886
rect 63500 26240 63552 26246
rect 63500 26182 63552 26188
rect 63408 24676 63460 24682
rect 63408 24618 63460 24624
rect 63512 24426 63540 26182
rect 63512 24398 63632 24426
rect 63500 24336 63552 24342
rect 63500 24278 63552 24284
rect 63408 24064 63460 24070
rect 63408 24006 63460 24012
rect 63420 23798 63448 24006
rect 63512 23798 63540 24278
rect 63408 23792 63460 23798
rect 63408 23734 63460 23740
rect 63500 23792 63552 23798
rect 63500 23734 63552 23740
rect 63604 22094 63632 24398
rect 63684 23044 63736 23050
rect 63684 22986 63736 22992
rect 63512 22066 63632 22094
rect 63512 18902 63540 22066
rect 63592 21344 63644 21350
rect 63590 21312 63592 21321
rect 63644 21312 63646 21321
rect 63590 21247 63646 21256
rect 63696 21010 63724 22986
rect 63684 21004 63736 21010
rect 63684 20946 63736 20952
rect 63696 20466 63724 20946
rect 64144 20800 64196 20806
rect 64144 20742 64196 20748
rect 63684 20460 63736 20466
rect 63684 20402 63736 20408
rect 63960 20392 64012 20398
rect 63960 20334 64012 20340
rect 64050 20360 64106 20369
rect 63972 19786 64000 20334
rect 64050 20295 64106 20304
rect 64064 20262 64092 20295
rect 64052 20256 64104 20262
rect 64052 20198 64104 20204
rect 63960 19780 64012 19786
rect 63960 19722 64012 19728
rect 63776 19712 63828 19718
rect 63776 19654 63828 19660
rect 63408 18896 63460 18902
rect 63408 18838 63460 18844
rect 63500 18896 63552 18902
rect 63500 18838 63552 18844
rect 63420 18442 63448 18838
rect 63420 18414 63724 18442
rect 63696 18358 63724 18414
rect 63592 18352 63644 18358
rect 63592 18294 63644 18300
rect 63684 18352 63736 18358
rect 63684 18294 63736 18300
rect 63408 15156 63460 15162
rect 63408 15098 63460 15104
rect 63420 14618 63448 15098
rect 63408 14612 63460 14618
rect 63408 14554 63460 14560
rect 63500 14476 63552 14482
rect 63500 14418 63552 14424
rect 63236 12406 63356 12434
rect 63236 10470 63264 12406
rect 63224 10464 63276 10470
rect 63224 10406 63276 10412
rect 63512 10130 63540 14418
rect 63408 10124 63460 10130
rect 63408 10066 63460 10072
rect 63500 10124 63552 10130
rect 63500 10066 63552 10072
rect 63420 9722 63448 10066
rect 63408 9716 63460 9722
rect 63408 9658 63460 9664
rect 63224 9512 63276 9518
rect 63224 9454 63276 9460
rect 63316 9512 63368 9518
rect 63316 9454 63368 9460
rect 63236 8974 63264 9454
rect 63224 8968 63276 8974
rect 63224 8910 63276 8916
rect 63328 8673 63356 9454
rect 63314 8664 63370 8673
rect 63314 8599 63370 8608
rect 63604 6866 63632 18294
rect 63682 14512 63738 14521
rect 63682 14447 63684 14456
rect 63736 14447 63738 14456
rect 63684 14418 63736 14424
rect 63684 13728 63736 13734
rect 63684 13670 63736 13676
rect 63696 12850 63724 13670
rect 63684 12844 63736 12850
rect 63684 12786 63736 12792
rect 63592 6860 63644 6866
rect 63592 6802 63644 6808
rect 63500 4140 63552 4146
rect 63500 4082 63552 4088
rect 63224 4072 63276 4078
rect 63224 4014 63276 4020
rect 63236 3398 63264 4014
rect 63224 3392 63276 3398
rect 63224 3334 63276 3340
rect 63132 2576 63184 2582
rect 63132 2518 63184 2524
rect 63408 2440 63460 2446
rect 63408 2382 63460 2388
rect 63316 2372 63368 2378
rect 63316 2314 63368 2320
rect 63328 800 63356 2314
rect 63420 2038 63448 2382
rect 63408 2032 63460 2038
rect 63408 1974 63460 1980
rect 63512 800 63540 4082
rect 63684 3528 63736 3534
rect 63684 3470 63736 3476
rect 63592 2984 63644 2990
rect 63592 2926 63644 2932
rect 63604 1154 63632 2926
rect 63592 1148 63644 1154
rect 63592 1090 63644 1096
rect 63696 800 63724 3470
rect 63788 2582 63816 19654
rect 64156 16250 64184 20742
rect 64144 16244 64196 16250
rect 64144 16186 64196 16192
rect 63960 12232 64012 12238
rect 63960 12174 64012 12180
rect 63868 9104 63920 9110
rect 63868 9046 63920 9052
rect 63880 8362 63908 9046
rect 63868 8356 63920 8362
rect 63868 8298 63920 8304
rect 63972 7750 64000 12174
rect 63960 7744 64012 7750
rect 63960 7686 64012 7692
rect 64248 4690 64276 34886
rect 64340 32910 64368 37266
rect 64604 36032 64656 36038
rect 64604 35974 64656 35980
rect 64616 35154 64644 35974
rect 64604 35148 64656 35154
rect 64604 35090 64656 35096
rect 64788 34196 64840 34202
rect 64788 34138 64840 34144
rect 64800 33998 64828 34138
rect 64788 33992 64840 33998
rect 64788 33934 64840 33940
rect 64328 32904 64380 32910
rect 64328 32846 64380 32852
rect 64328 28076 64380 28082
rect 64328 28018 64380 28024
rect 64340 11014 64368 28018
rect 64604 26444 64656 26450
rect 64604 26386 64656 26392
rect 64696 26444 64748 26450
rect 64696 26386 64748 26392
rect 64420 23044 64472 23050
rect 64420 22986 64472 22992
rect 64432 22642 64460 22986
rect 64420 22636 64472 22642
rect 64420 22578 64472 22584
rect 64616 22250 64644 26386
rect 64708 26314 64736 26386
rect 64696 26308 64748 26314
rect 64696 26250 64748 26256
rect 64696 23180 64748 23186
rect 64696 23122 64748 23128
rect 64708 22438 64736 23122
rect 64788 22704 64840 22710
rect 64788 22646 64840 22652
rect 64696 22432 64748 22438
rect 64696 22374 64748 22380
rect 64616 22222 64736 22250
rect 64604 22160 64656 22166
rect 64604 22102 64656 22108
rect 64420 21548 64472 21554
rect 64420 21490 64472 21496
rect 64432 20806 64460 21490
rect 64420 20800 64472 20806
rect 64420 20742 64472 20748
rect 64512 20528 64564 20534
rect 64510 20496 64512 20505
rect 64564 20496 64566 20505
rect 64510 20431 64566 20440
rect 64616 19446 64644 22102
rect 64604 19440 64656 19446
rect 64604 19382 64656 19388
rect 64512 18692 64564 18698
rect 64512 18634 64564 18640
rect 64328 11008 64380 11014
rect 64328 10950 64380 10956
rect 64524 8838 64552 18634
rect 64512 8832 64564 8838
rect 64512 8774 64564 8780
rect 64616 5166 64644 19382
rect 64604 5160 64656 5166
rect 64604 5102 64656 5108
rect 64418 4720 64474 4729
rect 64236 4684 64288 4690
rect 64236 4626 64288 4632
rect 64328 4684 64380 4690
rect 64418 4655 64474 4664
rect 64328 4626 64380 4632
rect 63868 4616 63920 4622
rect 64340 4570 64368 4626
rect 64432 4622 64460 4655
rect 63920 4564 64368 4570
rect 63868 4558 64368 4564
rect 64420 4616 64472 4622
rect 64420 4558 64472 4564
rect 63880 4542 64368 4558
rect 64052 3664 64104 3670
rect 64052 3606 64104 3612
rect 63776 2576 63828 2582
rect 63776 2518 63828 2524
rect 63868 2576 63920 2582
rect 63868 2518 63920 2524
rect 63880 800 63908 2518
rect 63960 2304 64012 2310
rect 63960 2246 64012 2252
rect 63972 2106 64000 2246
rect 63960 2100 64012 2106
rect 63960 2042 64012 2048
rect 64064 800 64092 3606
rect 64420 3052 64472 3058
rect 64420 2994 64472 3000
rect 64328 2984 64380 2990
rect 64328 2926 64380 2932
rect 64340 800 64368 2926
rect 64432 2514 64460 2994
rect 64708 2922 64736 22222
rect 64800 22166 64828 22646
rect 64788 22160 64840 22166
rect 64788 22102 64840 22108
rect 64786 20632 64842 20641
rect 64786 20567 64842 20576
rect 64800 20330 64828 20567
rect 64788 20324 64840 20330
rect 64788 20266 64840 20272
rect 64788 17740 64840 17746
rect 64788 17682 64840 17688
rect 64800 17202 64828 17682
rect 64788 17196 64840 17202
rect 64788 17138 64840 17144
rect 64788 7472 64840 7478
rect 64788 7414 64840 7420
rect 64800 5098 64828 7414
rect 64892 5166 64920 37606
rect 64972 37256 65024 37262
rect 64972 37198 65024 37204
rect 65064 37256 65116 37262
rect 65064 37198 65116 37204
rect 64984 36174 65012 37198
rect 65076 37126 65104 37198
rect 65064 37120 65116 37126
rect 65064 37062 65116 37068
rect 65156 37120 65208 37126
rect 65156 37062 65208 37068
rect 65064 36916 65116 36922
rect 65064 36858 65116 36864
rect 64972 36168 65024 36174
rect 64972 36110 65024 36116
rect 64972 34536 65024 34542
rect 64972 34478 65024 34484
rect 64984 34202 65012 34478
rect 64972 34196 65024 34202
rect 64972 34138 65024 34144
rect 64972 25356 65024 25362
rect 64972 25298 65024 25304
rect 64984 22817 65012 25298
rect 64970 22808 65026 22817
rect 64970 22743 65026 22752
rect 65076 22642 65104 36858
rect 65168 36786 65196 37062
rect 65156 36780 65208 36786
rect 65156 36722 65208 36728
rect 65260 36530 65288 39200
rect 66180 37398 66208 39200
rect 66444 37868 66496 37874
rect 66444 37810 66496 37816
rect 66456 37398 66484 37810
rect 66536 37800 66588 37806
rect 66536 37742 66588 37748
rect 66168 37392 66220 37398
rect 66168 37334 66220 37340
rect 66444 37392 66496 37398
rect 66444 37334 66496 37340
rect 65660 37020 65956 37040
rect 65716 37018 65740 37020
rect 65796 37018 65820 37020
rect 65876 37018 65900 37020
rect 65738 36966 65740 37018
rect 65802 36966 65814 37018
rect 65876 36966 65878 37018
rect 65716 36964 65740 36966
rect 65796 36964 65820 36966
rect 65876 36964 65900 36966
rect 65660 36944 65956 36964
rect 65432 36712 65484 36718
rect 65432 36654 65484 36660
rect 65168 36502 65288 36530
rect 65168 36106 65196 36502
rect 65444 36378 65472 36654
rect 65616 36644 65668 36650
rect 65616 36586 65668 36592
rect 65800 36644 65852 36650
rect 65800 36586 65852 36592
rect 65524 36576 65576 36582
rect 65524 36518 65576 36524
rect 65536 36378 65564 36518
rect 65432 36372 65484 36378
rect 65432 36314 65484 36320
rect 65524 36372 65576 36378
rect 65524 36314 65576 36320
rect 65340 36236 65392 36242
rect 65340 36178 65392 36184
rect 65156 36100 65208 36106
rect 65156 36042 65208 36048
rect 65156 35556 65208 35562
rect 65156 35498 65208 35504
rect 64972 22636 65024 22642
rect 64972 22578 65024 22584
rect 65064 22636 65116 22642
rect 65064 22578 65116 22584
rect 64984 22094 65012 22578
rect 65062 22536 65118 22545
rect 65062 22471 65064 22480
rect 65116 22471 65118 22480
rect 65064 22442 65116 22448
rect 64984 22066 65104 22094
rect 65076 20890 65104 22066
rect 65168 21554 65196 35498
rect 65352 31754 65380 36178
rect 65628 36174 65656 36586
rect 65812 36553 65840 36586
rect 65798 36544 65854 36553
rect 65854 36502 66024 36530
rect 65798 36479 65854 36488
rect 65616 36168 65668 36174
rect 65616 36110 65668 36116
rect 65660 35932 65956 35952
rect 65716 35930 65740 35932
rect 65796 35930 65820 35932
rect 65876 35930 65900 35932
rect 65738 35878 65740 35930
rect 65802 35878 65814 35930
rect 65876 35878 65878 35930
rect 65716 35876 65740 35878
rect 65796 35876 65820 35878
rect 65876 35876 65900 35878
rect 65660 35856 65956 35876
rect 65996 35222 66024 36502
rect 66168 36032 66220 36038
rect 66168 35974 66220 35980
rect 65984 35216 66036 35222
rect 65984 35158 66036 35164
rect 65660 34844 65956 34864
rect 65716 34842 65740 34844
rect 65796 34842 65820 34844
rect 65876 34842 65900 34844
rect 65738 34790 65740 34842
rect 65802 34790 65814 34842
rect 65876 34790 65878 34842
rect 65716 34788 65740 34790
rect 65796 34788 65820 34790
rect 65876 34788 65900 34790
rect 65660 34768 65956 34788
rect 65984 34536 66036 34542
rect 65984 34478 66036 34484
rect 65660 33756 65956 33776
rect 65716 33754 65740 33756
rect 65796 33754 65820 33756
rect 65876 33754 65900 33756
rect 65738 33702 65740 33754
rect 65802 33702 65814 33754
rect 65876 33702 65878 33754
rect 65716 33700 65740 33702
rect 65796 33700 65820 33702
rect 65876 33700 65900 33702
rect 65660 33680 65956 33700
rect 65996 33318 66024 34478
rect 65984 33312 66036 33318
rect 65984 33254 66036 33260
rect 65660 32668 65956 32688
rect 65716 32666 65740 32668
rect 65796 32666 65820 32668
rect 65876 32666 65900 32668
rect 65738 32614 65740 32666
rect 65802 32614 65814 32666
rect 65876 32614 65878 32666
rect 65716 32612 65740 32614
rect 65796 32612 65820 32614
rect 65876 32612 65900 32614
rect 65660 32592 65956 32612
rect 65352 31726 65564 31754
rect 65432 29844 65484 29850
rect 65432 29786 65484 29792
rect 65444 29238 65472 29786
rect 65432 29232 65484 29238
rect 65432 29174 65484 29180
rect 65536 26874 65564 31726
rect 65660 31580 65956 31600
rect 65716 31578 65740 31580
rect 65796 31578 65820 31580
rect 65876 31578 65900 31580
rect 65738 31526 65740 31578
rect 65802 31526 65814 31578
rect 65876 31526 65878 31578
rect 65716 31524 65740 31526
rect 65796 31524 65820 31526
rect 65876 31524 65900 31526
rect 65660 31504 65956 31524
rect 65660 30492 65956 30512
rect 65716 30490 65740 30492
rect 65796 30490 65820 30492
rect 65876 30490 65900 30492
rect 65738 30438 65740 30490
rect 65802 30438 65814 30490
rect 65876 30438 65878 30490
rect 65716 30436 65740 30438
rect 65796 30436 65820 30438
rect 65876 30436 65900 30438
rect 65660 30416 65956 30436
rect 65616 30320 65668 30326
rect 65616 30262 65668 30268
rect 65628 29617 65656 30262
rect 65614 29608 65670 29617
rect 65614 29543 65670 29552
rect 65660 29404 65956 29424
rect 65716 29402 65740 29404
rect 65796 29402 65820 29404
rect 65876 29402 65900 29404
rect 65738 29350 65740 29402
rect 65802 29350 65814 29402
rect 65876 29350 65878 29402
rect 65716 29348 65740 29350
rect 65796 29348 65820 29350
rect 65876 29348 65900 29350
rect 65660 29328 65956 29348
rect 65660 28316 65956 28336
rect 65716 28314 65740 28316
rect 65796 28314 65820 28316
rect 65876 28314 65900 28316
rect 65738 28262 65740 28314
rect 65802 28262 65814 28314
rect 65876 28262 65878 28314
rect 65716 28260 65740 28262
rect 65796 28260 65820 28262
rect 65876 28260 65900 28262
rect 65660 28240 65956 28260
rect 65660 27228 65956 27248
rect 65716 27226 65740 27228
rect 65796 27226 65820 27228
rect 65876 27226 65900 27228
rect 65738 27174 65740 27226
rect 65802 27174 65814 27226
rect 65876 27174 65878 27226
rect 65716 27172 65740 27174
rect 65796 27172 65820 27174
rect 65876 27172 65900 27174
rect 65660 27152 65956 27172
rect 65352 26846 65564 26874
rect 65248 25832 65300 25838
rect 65248 25774 65300 25780
rect 65260 25498 65288 25774
rect 65248 25492 65300 25498
rect 65248 25434 65300 25440
rect 65248 22976 65300 22982
rect 65248 22918 65300 22924
rect 65260 22574 65288 22918
rect 65248 22568 65300 22574
rect 65248 22510 65300 22516
rect 65246 22400 65302 22409
rect 65246 22335 65302 22344
rect 65260 21554 65288 22335
rect 65156 21548 65208 21554
rect 65156 21490 65208 21496
rect 65248 21548 65300 21554
rect 65248 21490 65300 21496
rect 64984 20862 65104 20890
rect 64984 17678 65012 20862
rect 65064 20800 65116 20806
rect 65064 20742 65116 20748
rect 65156 20800 65208 20806
rect 65156 20742 65208 20748
rect 65076 20262 65104 20742
rect 65168 20398 65196 20742
rect 65156 20392 65208 20398
rect 65248 20392 65300 20398
rect 65156 20334 65208 20340
rect 65246 20360 65248 20369
rect 65300 20360 65302 20369
rect 65246 20295 65302 20304
rect 65064 20256 65116 20262
rect 65064 20198 65116 20204
rect 64972 17672 65024 17678
rect 64972 17614 65024 17620
rect 65352 17354 65380 26846
rect 65432 26240 65484 26246
rect 65432 26182 65484 26188
rect 65444 26042 65472 26182
rect 65660 26140 65956 26160
rect 65716 26138 65740 26140
rect 65796 26138 65820 26140
rect 65876 26138 65900 26140
rect 65738 26086 65740 26138
rect 65802 26086 65814 26138
rect 65876 26086 65878 26138
rect 65716 26084 65740 26086
rect 65796 26084 65820 26086
rect 65876 26084 65900 26086
rect 65660 26064 65956 26084
rect 65432 26036 65484 26042
rect 65432 25978 65484 25984
rect 65432 25900 65484 25906
rect 65432 25842 65484 25848
rect 65444 25430 65472 25842
rect 65432 25424 65484 25430
rect 65432 25366 65484 25372
rect 65614 25256 65670 25265
rect 65614 25191 65616 25200
rect 65668 25191 65670 25200
rect 65616 25162 65668 25168
rect 65660 25052 65956 25072
rect 65716 25050 65740 25052
rect 65796 25050 65820 25052
rect 65876 25050 65900 25052
rect 65738 24998 65740 25050
rect 65802 24998 65814 25050
rect 65876 24998 65878 25050
rect 65716 24996 65740 24998
rect 65796 24996 65820 24998
rect 65876 24996 65900 24998
rect 65660 24976 65956 24996
rect 65524 24744 65576 24750
rect 65524 24686 65576 24692
rect 65536 24410 65564 24686
rect 65524 24404 65576 24410
rect 65524 24346 65576 24352
rect 65432 24064 65484 24070
rect 65432 24006 65484 24012
rect 65444 23594 65472 24006
rect 65660 23964 65956 23984
rect 65716 23962 65740 23964
rect 65796 23962 65820 23964
rect 65876 23962 65900 23964
rect 65738 23910 65740 23962
rect 65802 23910 65814 23962
rect 65876 23910 65878 23962
rect 65716 23908 65740 23910
rect 65796 23908 65820 23910
rect 65876 23908 65900 23910
rect 65660 23888 65956 23908
rect 65616 23656 65668 23662
rect 65892 23656 65944 23662
rect 65668 23604 65892 23610
rect 65616 23598 65944 23604
rect 65432 23588 65484 23594
rect 65628 23582 65932 23598
rect 65432 23530 65484 23536
rect 65892 23520 65944 23526
rect 65892 23462 65944 23468
rect 65904 23089 65932 23462
rect 65890 23080 65946 23089
rect 65890 23015 65946 23024
rect 65660 22876 65956 22896
rect 65716 22874 65740 22876
rect 65796 22874 65820 22876
rect 65876 22874 65900 22876
rect 65738 22822 65740 22874
rect 65802 22822 65814 22874
rect 65876 22822 65878 22874
rect 65716 22820 65740 22822
rect 65796 22820 65820 22822
rect 65876 22820 65900 22822
rect 65660 22800 65956 22820
rect 65432 22704 65484 22710
rect 65484 22652 65748 22658
rect 65432 22646 65748 22652
rect 65444 22630 65748 22646
rect 65720 22574 65748 22630
rect 65432 22568 65484 22574
rect 65432 22510 65484 22516
rect 65708 22568 65760 22574
rect 65708 22510 65760 22516
rect 64984 17326 65380 17354
rect 64984 13326 65012 17326
rect 65444 17218 65472 22510
rect 65660 21788 65956 21808
rect 65716 21786 65740 21788
rect 65796 21786 65820 21788
rect 65876 21786 65900 21788
rect 65738 21734 65740 21786
rect 65802 21734 65814 21786
rect 65876 21734 65878 21786
rect 65716 21732 65740 21734
rect 65796 21732 65820 21734
rect 65876 21732 65900 21734
rect 65660 21712 65956 21732
rect 65522 21584 65578 21593
rect 65522 21519 65578 21528
rect 65536 18816 65564 21519
rect 65996 21298 66024 33254
rect 66180 31754 66208 35974
rect 66088 31726 66208 31754
rect 66548 31754 66576 37742
rect 67008 37482 67036 39200
rect 67928 37890 67956 39200
rect 67928 37862 68324 37890
rect 67008 37466 67220 37482
rect 67008 37460 67232 37466
rect 67008 37454 67180 37460
rect 67180 37402 67232 37408
rect 66996 37324 67048 37330
rect 66996 37266 67048 37272
rect 67008 35766 67036 37266
rect 67836 36786 68232 36802
rect 67732 36780 67784 36786
rect 67732 36722 67784 36728
rect 67836 36780 68244 36786
rect 67836 36774 68192 36780
rect 67744 35766 67772 36722
rect 67836 36718 67864 36774
rect 68192 36722 68244 36728
rect 67824 36712 67876 36718
rect 67824 36654 67876 36660
rect 68296 36650 68324 37862
rect 68756 37330 68784 39200
rect 68836 38616 68888 38622
rect 68836 38558 68888 38564
rect 68744 37324 68796 37330
rect 68744 37266 68796 37272
rect 68560 37256 68612 37262
rect 68560 37198 68612 37204
rect 68468 36712 68520 36718
rect 68468 36654 68520 36660
rect 68008 36644 68060 36650
rect 68008 36586 68060 36592
rect 68284 36644 68336 36650
rect 68284 36586 68336 36592
rect 66996 35760 67048 35766
rect 66996 35702 67048 35708
rect 67732 35760 67784 35766
rect 67732 35702 67784 35708
rect 67008 35630 67036 35702
rect 66720 35624 66772 35630
rect 66720 35566 66772 35572
rect 66996 35624 67048 35630
rect 66996 35566 67048 35572
rect 66548 31726 66668 31754
rect 66088 21434 66116 31726
rect 66536 29640 66588 29646
rect 66534 29608 66536 29617
rect 66588 29608 66590 29617
rect 66534 29543 66590 29552
rect 66352 25832 66404 25838
rect 66352 25774 66404 25780
rect 66260 24948 66312 24954
rect 66260 24890 66312 24896
rect 66272 24342 66300 24890
rect 66260 24336 66312 24342
rect 66260 24278 66312 24284
rect 66168 23248 66220 23254
rect 66168 23190 66220 23196
rect 66180 21593 66208 23190
rect 66260 21684 66312 21690
rect 66260 21626 66312 21632
rect 66166 21584 66222 21593
rect 66166 21519 66222 21528
rect 66088 21406 66208 21434
rect 65996 21270 66116 21298
rect 65660 20700 65956 20720
rect 65716 20698 65740 20700
rect 65796 20698 65820 20700
rect 65876 20698 65900 20700
rect 65738 20646 65740 20698
rect 65802 20646 65814 20698
rect 65876 20646 65878 20698
rect 65716 20644 65740 20646
rect 65796 20644 65820 20646
rect 65876 20644 65900 20646
rect 65660 20624 65956 20644
rect 65982 20496 66038 20505
rect 65982 20431 66038 20440
rect 65996 20262 66024 20431
rect 65984 20256 66036 20262
rect 65984 20198 66036 20204
rect 65660 19612 65956 19632
rect 65716 19610 65740 19612
rect 65796 19610 65820 19612
rect 65876 19610 65900 19612
rect 65738 19558 65740 19610
rect 65802 19558 65814 19610
rect 65876 19558 65878 19610
rect 65716 19556 65740 19558
rect 65796 19556 65820 19558
rect 65876 19556 65900 19558
rect 65660 19536 65956 19556
rect 65536 18788 66024 18816
rect 65524 18692 65576 18698
rect 65524 18634 65576 18640
rect 65536 18426 65564 18634
rect 65660 18524 65956 18544
rect 65716 18522 65740 18524
rect 65796 18522 65820 18524
rect 65876 18522 65900 18524
rect 65738 18470 65740 18522
rect 65802 18470 65814 18522
rect 65876 18470 65878 18522
rect 65716 18468 65740 18470
rect 65796 18468 65820 18470
rect 65876 18468 65900 18470
rect 65660 18448 65956 18468
rect 65524 18420 65576 18426
rect 65524 18362 65576 18368
rect 65616 18352 65668 18358
rect 65800 18352 65852 18358
rect 65668 18300 65800 18306
rect 65616 18294 65852 18300
rect 65524 18284 65576 18290
rect 65628 18278 65840 18294
rect 65524 18226 65576 18232
rect 65168 17190 65472 17218
rect 65064 16584 65116 16590
rect 65064 16526 65116 16532
rect 65076 15366 65104 16526
rect 65064 15360 65116 15366
rect 65064 15302 65116 15308
rect 64972 13320 65024 13326
rect 64972 13262 65024 13268
rect 65064 12912 65116 12918
rect 65064 12854 65116 12860
rect 64972 12300 65024 12306
rect 64972 12242 65024 12248
rect 64984 10606 65012 12242
rect 65076 11121 65104 12854
rect 65062 11112 65118 11121
rect 65062 11047 65118 11056
rect 64972 10600 65024 10606
rect 64972 10542 65024 10548
rect 65076 9674 65104 11047
rect 64984 9646 65104 9674
rect 64984 7478 65012 9646
rect 65062 8936 65118 8945
rect 65062 8871 65118 8880
rect 65076 7834 65104 8871
rect 65168 7993 65196 17190
rect 65536 17082 65564 18226
rect 65660 17436 65956 17456
rect 65716 17434 65740 17436
rect 65796 17434 65820 17436
rect 65876 17434 65900 17436
rect 65738 17382 65740 17434
rect 65802 17382 65814 17434
rect 65876 17382 65878 17434
rect 65716 17380 65740 17382
rect 65796 17380 65820 17382
rect 65876 17380 65900 17382
rect 65660 17360 65956 17380
rect 65444 17054 65564 17082
rect 65248 16584 65300 16590
rect 65248 16526 65300 16532
rect 65260 12918 65288 16526
rect 65444 16250 65472 17054
rect 65524 16448 65576 16454
rect 65524 16390 65576 16396
rect 65432 16244 65484 16250
rect 65432 16186 65484 16192
rect 65536 16182 65564 16390
rect 65660 16348 65956 16368
rect 65716 16346 65740 16348
rect 65796 16346 65820 16348
rect 65876 16346 65900 16348
rect 65738 16294 65740 16346
rect 65802 16294 65814 16346
rect 65876 16294 65878 16346
rect 65716 16292 65740 16294
rect 65796 16292 65820 16294
rect 65876 16292 65900 16294
rect 65660 16272 65956 16292
rect 65524 16176 65576 16182
rect 65524 16118 65576 16124
rect 65340 16108 65392 16114
rect 65340 16050 65392 16056
rect 65352 15910 65380 16050
rect 65340 15904 65392 15910
rect 65340 15846 65392 15852
rect 65432 15904 65484 15910
rect 65432 15846 65484 15852
rect 65444 15706 65472 15846
rect 65432 15700 65484 15706
rect 65432 15642 65484 15648
rect 65616 15632 65668 15638
rect 65614 15600 65616 15609
rect 65668 15600 65670 15609
rect 65432 15564 65484 15570
rect 65614 15535 65670 15544
rect 65432 15506 65484 15512
rect 65248 12912 65300 12918
rect 65248 12854 65300 12860
rect 65444 12866 65472 15506
rect 65660 15260 65956 15280
rect 65716 15258 65740 15260
rect 65796 15258 65820 15260
rect 65876 15258 65900 15260
rect 65738 15206 65740 15258
rect 65802 15206 65814 15258
rect 65876 15206 65878 15258
rect 65716 15204 65740 15206
rect 65796 15204 65820 15206
rect 65876 15204 65900 15206
rect 65660 15184 65956 15204
rect 65660 14172 65956 14192
rect 65716 14170 65740 14172
rect 65796 14170 65820 14172
rect 65876 14170 65900 14172
rect 65738 14118 65740 14170
rect 65802 14118 65814 14170
rect 65876 14118 65878 14170
rect 65716 14116 65740 14118
rect 65796 14116 65820 14118
rect 65876 14116 65900 14118
rect 65660 14096 65956 14116
rect 65996 14056 66024 18788
rect 65904 14028 66024 14056
rect 65524 13796 65576 13802
rect 65524 13738 65576 13744
rect 65536 13394 65564 13738
rect 65524 13388 65576 13394
rect 65524 13330 65576 13336
rect 65904 13274 65932 14028
rect 65984 13932 66036 13938
rect 65984 13874 66036 13880
rect 65996 13734 66024 13874
rect 65984 13728 66036 13734
rect 65984 13670 66036 13676
rect 65996 13462 66024 13670
rect 65984 13456 66036 13462
rect 65984 13398 66036 13404
rect 65904 13246 66024 13274
rect 65660 13084 65956 13104
rect 65716 13082 65740 13084
rect 65796 13082 65820 13084
rect 65876 13082 65900 13084
rect 65738 13030 65740 13082
rect 65802 13030 65814 13082
rect 65876 13030 65878 13082
rect 65716 13028 65740 13030
rect 65796 13028 65820 13030
rect 65876 13028 65900 13030
rect 65660 13008 65956 13028
rect 65444 12838 65840 12866
rect 65432 12708 65484 12714
rect 65432 12650 65484 12656
rect 65444 12442 65472 12650
rect 65432 12436 65484 12442
rect 65432 12378 65484 12384
rect 65524 12232 65576 12238
rect 65524 12174 65576 12180
rect 65812 12186 65840 12838
rect 65996 12714 66024 13246
rect 65984 12708 66036 12714
rect 65984 12650 66036 12656
rect 65892 12436 65944 12442
rect 66088 12434 66116 21270
rect 66180 16590 66208 21406
rect 66272 21350 66300 21626
rect 66260 21344 66312 21350
rect 66260 21286 66312 21292
rect 66260 18420 66312 18426
rect 66260 18362 66312 18368
rect 66272 18329 66300 18362
rect 66258 18320 66314 18329
rect 66258 18255 66314 18264
rect 66260 17672 66312 17678
rect 66260 17614 66312 17620
rect 66168 16584 66220 16590
rect 66168 16526 66220 16532
rect 66272 16250 66300 17614
rect 66168 16244 66220 16250
rect 66168 16186 66220 16192
rect 66260 16244 66312 16250
rect 66260 16186 66312 16192
rect 66180 13462 66208 16186
rect 66260 13932 66312 13938
rect 66260 13874 66312 13880
rect 66168 13456 66220 13462
rect 66168 13398 66220 13404
rect 66272 13274 66300 13874
rect 66180 13246 66300 13274
rect 66180 12782 66208 13246
rect 66168 12776 66220 12782
rect 66168 12718 66220 12724
rect 66088 12406 66208 12434
rect 65892 12378 65944 12384
rect 65904 12306 65932 12378
rect 65892 12300 65944 12306
rect 65892 12242 65944 12248
rect 65340 12096 65392 12102
rect 65340 12038 65392 12044
rect 65248 10532 65300 10538
rect 65248 10474 65300 10480
rect 65260 10266 65288 10474
rect 65248 10260 65300 10266
rect 65248 10202 65300 10208
rect 65352 9450 65380 12038
rect 65536 11830 65564 12174
rect 65812 12158 66116 12186
rect 65660 11996 65956 12016
rect 65716 11994 65740 11996
rect 65796 11994 65820 11996
rect 65876 11994 65900 11996
rect 65738 11942 65740 11994
rect 65802 11942 65814 11994
rect 65876 11942 65878 11994
rect 65716 11940 65740 11942
rect 65796 11940 65820 11942
rect 65876 11940 65900 11942
rect 65660 11920 65956 11940
rect 65524 11824 65576 11830
rect 65524 11766 65576 11772
rect 65660 10908 65956 10928
rect 65716 10906 65740 10908
rect 65796 10906 65820 10908
rect 65876 10906 65900 10908
rect 65738 10854 65740 10906
rect 65802 10854 65814 10906
rect 65876 10854 65878 10906
rect 65716 10852 65740 10854
rect 65796 10852 65820 10854
rect 65876 10852 65900 10854
rect 65660 10832 65956 10852
rect 65660 9820 65956 9840
rect 65716 9818 65740 9820
rect 65796 9818 65820 9820
rect 65876 9818 65900 9820
rect 65738 9766 65740 9818
rect 65802 9766 65814 9818
rect 65876 9766 65878 9818
rect 65716 9764 65740 9766
rect 65796 9764 65820 9766
rect 65876 9764 65900 9766
rect 65660 9744 65956 9764
rect 65522 9480 65578 9489
rect 65340 9444 65392 9450
rect 65522 9415 65524 9424
rect 65340 9386 65392 9392
rect 65576 9415 65578 9424
rect 65524 9386 65576 9392
rect 65524 8968 65576 8974
rect 65524 8910 65576 8916
rect 65536 8430 65564 8910
rect 65660 8732 65956 8752
rect 65716 8730 65740 8732
rect 65796 8730 65820 8732
rect 65876 8730 65900 8732
rect 65738 8678 65740 8730
rect 65802 8678 65814 8730
rect 65876 8678 65878 8730
rect 65716 8676 65740 8678
rect 65796 8676 65820 8678
rect 65876 8676 65900 8678
rect 65660 8656 65956 8676
rect 65524 8424 65576 8430
rect 65524 8366 65576 8372
rect 65984 8424 66036 8430
rect 65984 8366 66036 8372
rect 65248 8356 65300 8362
rect 65248 8298 65300 8304
rect 65154 7984 65210 7993
rect 65154 7919 65210 7928
rect 65076 7806 65196 7834
rect 64972 7472 65024 7478
rect 64972 7414 65024 7420
rect 65168 5302 65196 7806
rect 64972 5296 65024 5302
rect 64972 5238 65024 5244
rect 65156 5296 65208 5302
rect 65156 5238 65208 5244
rect 64880 5160 64932 5166
rect 64984 5148 65012 5238
rect 65064 5160 65116 5166
rect 64984 5120 65064 5148
rect 64880 5102 64932 5108
rect 65156 5160 65208 5166
rect 65064 5102 65116 5108
rect 65154 5128 65156 5137
rect 65208 5128 65210 5137
rect 64788 5092 64840 5098
rect 65154 5063 65210 5072
rect 64788 5034 64840 5040
rect 64972 4548 65024 4554
rect 64972 4490 65024 4496
rect 64984 4457 65012 4490
rect 64970 4448 65026 4457
rect 64970 4383 65026 4392
rect 64788 4140 64840 4146
rect 64788 4082 64840 4088
rect 64512 2916 64564 2922
rect 64512 2858 64564 2864
rect 64696 2916 64748 2922
rect 64696 2858 64748 2864
rect 64420 2508 64472 2514
rect 64420 2450 64472 2456
rect 64524 800 64552 2858
rect 64800 2774 64828 4082
rect 64880 3596 64932 3602
rect 64880 3538 64932 3544
rect 64708 2746 64828 2774
rect 64708 800 64736 2746
rect 64892 800 64920 3538
rect 65064 1420 65116 1426
rect 65064 1362 65116 1368
rect 65076 800 65104 1362
rect 65260 1290 65288 8298
rect 65660 7644 65956 7664
rect 65716 7642 65740 7644
rect 65796 7642 65820 7644
rect 65876 7642 65900 7644
rect 65738 7590 65740 7642
rect 65802 7590 65814 7642
rect 65876 7590 65878 7642
rect 65716 7588 65740 7590
rect 65796 7588 65820 7590
rect 65876 7588 65900 7590
rect 65660 7568 65956 7588
rect 65340 7540 65392 7546
rect 65340 7482 65392 7488
rect 65352 5234 65380 7482
rect 65996 6662 66024 8366
rect 66088 8362 66116 12158
rect 66180 8430 66208 12406
rect 66168 8424 66220 8430
rect 66168 8366 66220 8372
rect 66076 8356 66128 8362
rect 66076 8298 66128 8304
rect 65984 6656 66036 6662
rect 65984 6598 66036 6604
rect 65660 6556 65956 6576
rect 65716 6554 65740 6556
rect 65796 6554 65820 6556
rect 65876 6554 65900 6556
rect 65738 6502 65740 6554
rect 65802 6502 65814 6554
rect 65876 6502 65878 6554
rect 65716 6500 65740 6502
rect 65796 6500 65820 6502
rect 65876 6500 65900 6502
rect 65660 6480 65956 6500
rect 65660 5468 65956 5488
rect 65716 5466 65740 5468
rect 65796 5466 65820 5468
rect 65876 5466 65900 5468
rect 65738 5414 65740 5466
rect 65802 5414 65814 5466
rect 65876 5414 65878 5466
rect 65716 5412 65740 5414
rect 65796 5412 65820 5414
rect 65876 5412 65900 5414
rect 65660 5392 65956 5412
rect 66168 5364 66220 5370
rect 66168 5306 66220 5312
rect 65524 5296 65576 5302
rect 65524 5238 65576 5244
rect 65340 5228 65392 5234
rect 65340 5170 65392 5176
rect 65536 5030 65564 5238
rect 65524 5024 65576 5030
rect 65524 4966 65576 4972
rect 66180 4758 66208 5306
rect 66168 4752 66220 4758
rect 66168 4694 66220 4700
rect 65432 4684 65484 4690
rect 65432 4626 65484 4632
rect 65984 4684 66036 4690
rect 65984 4626 66036 4632
rect 65340 4140 65392 4146
rect 65340 4082 65392 4088
rect 65248 1284 65300 1290
rect 65248 1226 65300 1232
rect 65352 800 65380 4082
rect 65444 2582 65472 4626
rect 65660 4380 65956 4400
rect 65716 4378 65740 4380
rect 65796 4378 65820 4380
rect 65876 4378 65900 4380
rect 65738 4326 65740 4378
rect 65802 4326 65814 4378
rect 65876 4326 65878 4378
rect 65716 4324 65740 4326
rect 65796 4324 65820 4326
rect 65876 4324 65900 4326
rect 65660 4304 65956 4324
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 65536 3126 65564 3470
rect 65660 3292 65956 3312
rect 65716 3290 65740 3292
rect 65796 3290 65820 3292
rect 65876 3290 65900 3292
rect 65738 3238 65740 3290
rect 65802 3238 65814 3290
rect 65876 3238 65878 3290
rect 65716 3236 65740 3238
rect 65796 3236 65820 3238
rect 65876 3236 65900 3238
rect 65660 3216 65956 3236
rect 65524 3120 65576 3126
rect 65524 3062 65576 3068
rect 65524 2984 65576 2990
rect 65524 2926 65576 2932
rect 65432 2576 65484 2582
rect 65432 2518 65484 2524
rect 65536 800 65564 2926
rect 65660 2204 65956 2224
rect 65716 2202 65740 2204
rect 65796 2202 65820 2204
rect 65876 2202 65900 2204
rect 65738 2150 65740 2202
rect 65802 2150 65814 2202
rect 65876 2150 65878 2202
rect 65716 2148 65740 2150
rect 65796 2148 65820 2150
rect 65876 2148 65900 2150
rect 65660 2128 65956 2148
rect 65708 1488 65760 1494
rect 65996 1442 66024 4626
rect 66168 2848 66220 2854
rect 66168 2790 66220 2796
rect 65708 1430 65760 1436
rect 65720 800 65748 1430
rect 65904 1414 66024 1442
rect 65904 800 65932 1414
rect 66180 800 66208 2790
rect 66260 2304 66312 2310
rect 66260 2246 66312 2252
rect 66272 1494 66300 2246
rect 66364 1902 66392 25774
rect 66444 25356 66496 25362
rect 66444 25298 66496 25304
rect 66456 12918 66484 25298
rect 66536 23044 66588 23050
rect 66536 22986 66588 22992
rect 66548 22642 66576 22986
rect 66536 22636 66588 22642
rect 66536 22578 66588 22584
rect 66536 13864 66588 13870
rect 66536 13806 66588 13812
rect 66444 12912 66496 12918
rect 66444 12854 66496 12860
rect 66456 12782 66484 12854
rect 66444 12776 66496 12782
rect 66444 12718 66496 12724
rect 66548 9994 66576 13806
rect 66536 9988 66588 9994
rect 66536 9930 66588 9936
rect 66536 4072 66588 4078
rect 66536 4014 66588 4020
rect 66352 1896 66404 1902
rect 66352 1838 66404 1844
rect 66260 1488 66312 1494
rect 66260 1430 66312 1436
rect 66352 1488 66404 1494
rect 66352 1430 66404 1436
rect 66364 800 66392 1430
rect 66548 800 66576 4014
rect 66640 2650 66668 31726
rect 66732 5658 66760 35566
rect 67100 34598 67588 34626
rect 67100 34542 67128 34598
rect 67560 34542 67588 34598
rect 67088 34536 67140 34542
rect 67088 34478 67140 34484
rect 67456 34536 67508 34542
rect 67456 34478 67508 34484
rect 67548 34536 67600 34542
rect 67548 34478 67600 34484
rect 67468 34406 67496 34478
rect 67456 34400 67508 34406
rect 67456 34342 67508 34348
rect 67086 33960 67142 33969
rect 66904 33924 66956 33930
rect 67086 33895 67142 33904
rect 66904 33866 66956 33872
rect 66812 31884 66864 31890
rect 66812 31826 66864 31832
rect 66824 7562 66852 31826
rect 66916 31754 66944 33866
rect 66916 31726 67036 31754
rect 66904 30592 66956 30598
rect 66904 30534 66956 30540
rect 66916 24682 66944 30534
rect 66904 24676 66956 24682
rect 66904 24618 66956 24624
rect 66904 14068 66956 14074
rect 66904 14010 66956 14016
rect 66916 13938 66944 14010
rect 66904 13932 66956 13938
rect 66904 13874 66956 13880
rect 67008 7750 67036 31726
rect 66996 7744 67048 7750
rect 66996 7686 67048 7692
rect 66824 7534 67036 7562
rect 66732 5630 66852 5658
rect 66720 3596 66772 3602
rect 66720 3538 66772 3544
rect 66628 2644 66680 2650
rect 66628 2586 66680 2592
rect 66732 800 66760 3538
rect 66824 3126 66852 5630
rect 66812 3120 66864 3126
rect 66812 3062 66864 3068
rect 66904 2916 66956 2922
rect 66904 2858 66956 2864
rect 66812 2372 66864 2378
rect 66812 2314 66864 2320
rect 66824 1426 66852 2314
rect 66812 1420 66864 1426
rect 66812 1362 66864 1368
rect 66916 800 66944 2858
rect 67008 2650 67036 7534
rect 67100 5302 67128 33895
rect 67824 33652 67876 33658
rect 67824 33594 67876 33600
rect 67548 30864 67600 30870
rect 67548 30806 67600 30812
rect 67560 29646 67588 30806
rect 67180 29640 67232 29646
rect 67456 29640 67508 29646
rect 67180 29582 67232 29588
rect 67454 29608 67456 29617
rect 67548 29640 67600 29646
rect 67508 29608 67510 29617
rect 67192 28966 67220 29582
rect 67548 29582 67600 29588
rect 67454 29543 67510 29552
rect 67836 29238 67864 33594
rect 67824 29232 67876 29238
rect 67824 29174 67876 29180
rect 67914 29064 67970 29073
rect 67914 28999 67916 29008
rect 67968 28999 67970 29008
rect 67916 28970 67968 28976
rect 67180 28960 67232 28966
rect 67180 28902 67232 28908
rect 67192 25838 67220 28902
rect 67180 25832 67232 25838
rect 67180 25774 67232 25780
rect 67548 25832 67600 25838
rect 67548 25774 67600 25780
rect 67192 23118 67220 25774
rect 67272 24676 67324 24682
rect 67272 24618 67324 24624
rect 67180 23112 67232 23118
rect 67180 23054 67232 23060
rect 67284 19446 67312 24618
rect 67456 23112 67508 23118
rect 67456 23054 67508 23060
rect 67364 21004 67416 21010
rect 67364 20946 67416 20952
rect 67376 20913 67404 20946
rect 67362 20904 67418 20913
rect 67362 20839 67418 20848
rect 67468 20806 67496 23054
rect 67456 20800 67508 20806
rect 67456 20742 67508 20748
rect 67272 19440 67324 19446
rect 67272 19382 67324 19388
rect 67456 14408 67508 14414
rect 67456 14350 67508 14356
rect 67180 12912 67232 12918
rect 67180 12854 67232 12860
rect 67192 9518 67220 12854
rect 67364 12096 67416 12102
rect 67364 12038 67416 12044
rect 67272 11620 67324 11626
rect 67272 11562 67324 11568
rect 67284 10742 67312 11562
rect 67272 10736 67324 10742
rect 67272 10678 67324 10684
rect 67376 10266 67404 12038
rect 67468 11354 67496 14350
rect 67456 11348 67508 11354
rect 67456 11290 67508 11296
rect 67364 10260 67416 10266
rect 67364 10202 67416 10208
rect 67180 9512 67232 9518
rect 67180 9454 67232 9460
rect 67364 9104 67416 9110
rect 67364 9046 67416 9052
rect 67376 8634 67404 9046
rect 67364 8628 67416 8634
rect 67364 8570 67416 8576
rect 67468 8430 67496 11290
rect 67456 8424 67508 8430
rect 67456 8366 67508 8372
rect 67272 7744 67324 7750
rect 67272 7686 67324 7692
rect 67088 5296 67140 5302
rect 67088 5238 67140 5244
rect 67180 4072 67232 4078
rect 67180 4014 67232 4020
rect 66996 2644 67048 2650
rect 66996 2586 67048 2592
rect 67192 800 67220 4014
rect 67284 3058 67312 7686
rect 67272 3052 67324 3058
rect 67272 2994 67324 3000
rect 67364 2916 67416 2922
rect 67364 2858 67416 2864
rect 67376 800 67404 2858
rect 67560 2774 67588 25774
rect 67640 23112 67692 23118
rect 67640 23054 67692 23060
rect 67652 11558 67680 23054
rect 67824 18352 67876 18358
rect 67824 18294 67876 18300
rect 67732 16652 67784 16658
rect 67732 16594 67784 16600
rect 67640 11552 67692 11558
rect 67640 11494 67692 11500
rect 67744 7886 67772 16594
rect 67836 11286 67864 18294
rect 68020 15162 68048 36586
rect 68480 36582 68508 36654
rect 68572 36582 68600 37198
rect 68468 36576 68520 36582
rect 68468 36518 68520 36524
rect 68560 36576 68612 36582
rect 68560 36518 68612 36524
rect 68100 35148 68152 35154
rect 68100 35090 68152 35096
rect 68192 35148 68244 35154
rect 68192 35090 68244 35096
rect 68112 32298 68140 35090
rect 68100 32292 68152 32298
rect 68100 32234 68152 32240
rect 68112 27334 68140 32234
rect 68100 27328 68152 27334
rect 68100 27270 68152 27276
rect 68008 15156 68060 15162
rect 68008 15098 68060 15104
rect 68020 14958 68048 15098
rect 68008 14952 68060 14958
rect 68008 14894 68060 14900
rect 67824 11280 67876 11286
rect 67824 11222 67876 11228
rect 68100 8560 68152 8566
rect 68100 8502 68152 8508
rect 68112 8362 68140 8502
rect 68100 8356 68152 8362
rect 68100 8298 68152 8304
rect 67732 7880 67784 7886
rect 67732 7822 67784 7828
rect 68204 7002 68232 35090
rect 68480 34066 68508 36518
rect 68848 35154 68876 38558
rect 69676 37482 69704 39200
rect 70400 38004 70452 38010
rect 70400 37946 70452 37952
rect 70124 37732 70176 37738
rect 70124 37674 70176 37680
rect 69676 37466 69796 37482
rect 69676 37460 69808 37466
rect 69676 37454 69756 37460
rect 69756 37402 69808 37408
rect 68926 37360 68982 37369
rect 68926 37295 68982 37304
rect 69480 37324 69532 37330
rect 68940 37194 68968 37295
rect 69480 37266 69532 37272
rect 68928 37188 68980 37194
rect 68928 37130 68980 37136
rect 68836 35148 68888 35154
rect 68836 35090 68888 35096
rect 68744 35080 68796 35086
rect 68744 35022 68796 35028
rect 68468 34060 68520 34066
rect 68468 34002 68520 34008
rect 68468 30184 68520 30190
rect 68468 30126 68520 30132
rect 68560 30184 68612 30190
rect 68560 30126 68612 30132
rect 68284 30048 68336 30054
rect 68284 29990 68336 29996
rect 68296 29850 68324 29990
rect 68284 29844 68336 29850
rect 68284 29786 68336 29792
rect 68282 29200 68338 29209
rect 68282 29135 68338 29144
rect 68296 28966 68324 29135
rect 68480 29102 68508 30126
rect 68572 29646 68600 30126
rect 68560 29640 68612 29646
rect 68560 29582 68612 29588
rect 68652 29640 68704 29646
rect 68652 29582 68704 29588
rect 68560 29504 68612 29510
rect 68664 29458 68692 29582
rect 68612 29452 68692 29458
rect 68560 29446 68692 29452
rect 68572 29430 68692 29446
rect 68468 29096 68520 29102
rect 68468 29038 68520 29044
rect 68284 28960 68336 28966
rect 68284 28902 68336 28908
rect 68376 28144 68428 28150
rect 68376 28086 68428 28092
rect 68282 10568 68338 10577
rect 68282 10503 68338 10512
rect 68296 10470 68324 10503
rect 68284 10464 68336 10470
rect 68284 10406 68336 10412
rect 68282 9752 68338 9761
rect 68388 9722 68416 28086
rect 68572 22094 68600 29430
rect 68652 29232 68704 29238
rect 68652 29174 68704 29180
rect 68664 29102 68692 29174
rect 68652 29096 68704 29102
rect 68652 29038 68704 29044
rect 68480 22066 68600 22094
rect 68480 15638 68508 22066
rect 68468 15632 68520 15638
rect 68468 15574 68520 15580
rect 68282 9687 68284 9696
rect 68336 9687 68338 9696
rect 68376 9716 68428 9722
rect 68284 9658 68336 9664
rect 68376 9658 68428 9664
rect 68284 9444 68336 9450
rect 68284 9386 68336 9392
rect 68296 8566 68324 9386
rect 68284 8560 68336 8566
rect 68284 8502 68336 8508
rect 68192 6996 68244 7002
rect 68192 6938 68244 6944
rect 68480 6798 68508 15574
rect 68560 15156 68612 15162
rect 68560 15098 68612 15104
rect 68468 6792 68520 6798
rect 68468 6734 68520 6740
rect 67640 5636 67692 5642
rect 67640 5578 67692 5584
rect 67652 4486 67680 5578
rect 68572 5302 68600 15098
rect 68652 10600 68704 10606
rect 68652 10542 68704 10548
rect 68664 10169 68692 10542
rect 68650 10160 68706 10169
rect 68650 10095 68706 10104
rect 68756 9450 68784 35022
rect 68848 32774 68876 35090
rect 68928 35080 68980 35086
rect 68928 35022 68980 35028
rect 68940 34542 68968 35022
rect 68928 34536 68980 34542
rect 68928 34478 68980 34484
rect 69204 34400 69256 34406
rect 69204 34342 69256 34348
rect 69296 34400 69348 34406
rect 69296 34342 69348 34348
rect 68928 32904 68980 32910
rect 68928 32846 68980 32852
rect 68836 32768 68888 32774
rect 68836 32710 68888 32716
rect 68940 29646 68968 32846
rect 69112 30388 69164 30394
rect 69112 30330 69164 30336
rect 68928 29640 68980 29646
rect 68928 29582 68980 29588
rect 68836 29232 68888 29238
rect 68836 29174 68888 29180
rect 68848 26858 68876 29174
rect 68928 29096 68980 29102
rect 68928 29038 68980 29044
rect 68940 28150 68968 29038
rect 68928 28144 68980 28150
rect 68928 28086 68980 28092
rect 68836 26852 68888 26858
rect 68836 26794 68888 26800
rect 69020 26852 69072 26858
rect 69020 26794 69072 26800
rect 69032 23662 69060 26794
rect 69124 25974 69152 30330
rect 69112 25968 69164 25974
rect 69112 25910 69164 25916
rect 69020 23656 69072 23662
rect 69020 23598 69072 23604
rect 69112 22976 69164 22982
rect 69112 22918 69164 22924
rect 69020 19168 69072 19174
rect 69020 19110 69072 19116
rect 69032 13870 69060 19110
rect 69020 13864 69072 13870
rect 69020 13806 69072 13812
rect 69124 13326 69152 22918
rect 69112 13320 69164 13326
rect 69112 13262 69164 13268
rect 69112 10736 69164 10742
rect 69112 10678 69164 10684
rect 69124 10577 69152 10678
rect 69110 10568 69166 10577
rect 69110 10503 69166 10512
rect 68744 9444 68796 9450
rect 68744 9386 68796 9392
rect 68100 5296 68152 5302
rect 68100 5238 68152 5244
rect 68560 5296 68612 5302
rect 68560 5238 68612 5244
rect 67640 4480 67692 4486
rect 67640 4422 67692 4428
rect 67824 4072 67876 4078
rect 67824 4014 67876 4020
rect 67836 2774 67864 4014
rect 67916 3596 67968 3602
rect 67916 3538 67968 3544
rect 67468 2746 67588 2774
rect 67744 2746 67864 2774
rect 62396 264 62448 270
rect 62396 206 62448 212
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63498 0 63554 800
rect 63682 0 63738 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65338 0 65394 800
rect 65522 0 65578 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67468 513 67496 2746
rect 67548 2100 67600 2106
rect 67548 2042 67600 2048
rect 67560 800 67588 2042
rect 67744 800 67772 2746
rect 67928 800 67956 3538
rect 68112 2650 68140 5238
rect 68836 5024 68888 5030
rect 68836 4966 68888 4972
rect 68376 4684 68428 4690
rect 68376 4626 68428 4632
rect 68192 2848 68244 2854
rect 68192 2790 68244 2796
rect 68100 2644 68152 2650
rect 68100 2586 68152 2592
rect 68204 800 68232 2790
rect 68388 800 68416 4626
rect 68560 3596 68612 3602
rect 68560 3538 68612 3544
rect 68468 2372 68520 2378
rect 68468 2314 68520 2320
rect 68480 1494 68508 2314
rect 68468 1488 68520 1494
rect 68468 1430 68520 1436
rect 68572 800 68600 3538
rect 68848 2650 68876 4966
rect 68928 4072 68980 4078
rect 68928 4014 68980 4020
rect 68836 2644 68888 2650
rect 68836 2586 68888 2592
rect 68744 2032 68796 2038
rect 68744 1974 68796 1980
rect 68756 800 68784 1974
rect 68940 800 68968 4014
rect 69216 3754 69244 34342
rect 69308 33522 69336 34342
rect 69296 33516 69348 33522
rect 69296 33458 69348 33464
rect 69492 31754 69520 37266
rect 70032 37120 70084 37126
rect 69570 37088 69626 37097
rect 70032 37062 70084 37068
rect 69570 37023 69626 37032
rect 69308 31726 69520 31754
rect 69308 25809 69336 31726
rect 69480 30592 69532 30598
rect 69480 30534 69532 30540
rect 69386 29064 69442 29073
rect 69386 28999 69388 29008
rect 69440 28999 69442 29008
rect 69388 28970 69440 28976
rect 69492 28422 69520 30534
rect 69480 28416 69532 28422
rect 69480 28358 69532 28364
rect 69294 25800 69350 25809
rect 69294 25735 69350 25744
rect 69308 24954 69336 25735
rect 69296 24948 69348 24954
rect 69296 24890 69348 24896
rect 69492 22094 69520 28358
rect 69400 22066 69520 22094
rect 69296 18896 69348 18902
rect 69294 18864 69296 18873
rect 69348 18864 69350 18873
rect 69294 18799 69350 18808
rect 69296 17196 69348 17202
rect 69296 17138 69348 17144
rect 69308 11354 69336 17138
rect 69400 16794 69428 22066
rect 69480 19440 69532 19446
rect 69480 19382 69532 19388
rect 69492 18834 69520 19382
rect 69480 18828 69532 18834
rect 69480 18770 69532 18776
rect 69388 16788 69440 16794
rect 69388 16730 69440 16736
rect 69400 15570 69520 15586
rect 69388 15564 69520 15570
rect 69440 15558 69520 15564
rect 69388 15506 69440 15512
rect 69492 11762 69520 15558
rect 69480 11756 69532 11762
rect 69480 11698 69532 11704
rect 69480 11620 69532 11626
rect 69480 11562 69532 11568
rect 69296 11348 69348 11354
rect 69296 11290 69348 11296
rect 69492 7410 69520 11562
rect 69584 7546 69612 37023
rect 70044 35154 70072 37062
rect 70032 35148 70084 35154
rect 70032 35090 70084 35096
rect 70136 33658 70164 37674
rect 70214 36272 70270 36281
rect 70214 36207 70216 36216
rect 70268 36207 70270 36216
rect 70308 36236 70360 36242
rect 70216 36178 70268 36184
rect 70308 36178 70360 36184
rect 70320 33980 70348 36178
rect 70228 33952 70348 33980
rect 70124 33652 70176 33658
rect 70124 33594 70176 33600
rect 69664 32768 69716 32774
rect 69664 32710 69716 32716
rect 69676 31890 69704 32710
rect 69664 31884 69716 31890
rect 69664 31826 69716 31832
rect 69676 15638 69704 31826
rect 70228 30394 70256 33952
rect 70308 33652 70360 33658
rect 70308 33594 70360 33600
rect 70216 30388 70268 30394
rect 70216 30330 70268 30336
rect 69848 27940 69900 27946
rect 69848 27882 69900 27888
rect 69756 27668 69808 27674
rect 69756 27610 69808 27616
rect 69768 20398 69796 27610
rect 69756 20392 69808 20398
rect 69756 20334 69808 20340
rect 69756 18828 69808 18834
rect 69756 18770 69808 18776
rect 69768 18358 69796 18770
rect 69756 18352 69808 18358
rect 69756 18294 69808 18300
rect 69756 18216 69808 18222
rect 69756 18158 69808 18164
rect 69768 16658 69796 18158
rect 69860 17202 69888 27882
rect 70124 25764 70176 25770
rect 70124 25706 70176 25712
rect 70136 25498 70164 25706
rect 70124 25492 70176 25498
rect 70124 25434 70176 25440
rect 70216 25492 70268 25498
rect 70216 25434 70268 25440
rect 69940 24880 69992 24886
rect 69940 24822 69992 24828
rect 69952 23798 69980 24822
rect 69940 23792 69992 23798
rect 69940 23734 69992 23740
rect 70136 20398 70164 25434
rect 70228 25226 70256 25434
rect 70216 25220 70268 25226
rect 70216 25162 70268 25168
rect 70228 20466 70256 25162
rect 70216 20460 70268 20466
rect 70216 20402 70268 20408
rect 69940 20392 69992 20398
rect 69940 20334 69992 20340
rect 70124 20392 70176 20398
rect 70124 20334 70176 20340
rect 69848 17196 69900 17202
rect 69848 17138 69900 17144
rect 69848 16788 69900 16794
rect 69848 16730 69900 16736
rect 69756 16652 69808 16658
rect 69756 16594 69808 16600
rect 69768 16046 69796 16594
rect 69756 16040 69808 16046
rect 69756 15982 69808 15988
rect 69664 15632 69716 15638
rect 69664 15574 69716 15580
rect 69768 14958 69796 15982
rect 69756 14952 69808 14958
rect 69756 14894 69808 14900
rect 69664 14816 69716 14822
rect 69662 14784 69664 14793
rect 69716 14784 69718 14793
rect 69662 14719 69718 14728
rect 69768 13802 69796 14894
rect 69860 14482 69888 16730
rect 69848 14476 69900 14482
rect 69848 14418 69900 14424
rect 69756 13796 69808 13802
rect 69756 13738 69808 13744
rect 69768 12918 69796 13738
rect 69756 12912 69808 12918
rect 69756 12854 69808 12860
rect 69848 12708 69900 12714
rect 69848 12650 69900 12656
rect 69860 11354 69888 12650
rect 69848 11348 69900 11354
rect 69848 11290 69900 11296
rect 69952 9761 69980 20334
rect 70214 18864 70270 18873
rect 70214 18799 70270 18808
rect 70228 18290 70256 18799
rect 70216 18284 70268 18290
rect 70216 18226 70268 18232
rect 70032 18216 70084 18222
rect 70084 18176 70164 18204
rect 70032 18158 70084 18164
rect 70030 15192 70086 15201
rect 70030 15127 70086 15136
rect 70044 15094 70072 15127
rect 70032 15088 70084 15094
rect 70032 15030 70084 15036
rect 70032 13864 70084 13870
rect 70032 13806 70084 13812
rect 69938 9752 69994 9761
rect 69938 9687 69994 9696
rect 69572 7540 69624 7546
rect 69572 7482 69624 7488
rect 69480 7404 69532 7410
rect 69480 7346 69532 7352
rect 69480 6248 69532 6254
rect 69480 6190 69532 6196
rect 69492 6118 69520 6190
rect 69480 6112 69532 6118
rect 69480 6054 69532 6060
rect 69952 5642 69980 9687
rect 69940 5636 69992 5642
rect 69940 5578 69992 5584
rect 69572 4140 69624 4146
rect 69572 4082 69624 4088
rect 69216 3726 69336 3754
rect 69204 3596 69256 3602
rect 69204 3538 69256 3544
rect 69216 800 69244 3538
rect 69308 3126 69336 3726
rect 69296 3120 69348 3126
rect 69296 3062 69348 3068
rect 69388 2916 69440 2922
rect 69388 2858 69440 2864
rect 69296 2848 69348 2854
rect 69296 2790 69348 2796
rect 69308 2514 69336 2790
rect 69296 2508 69348 2514
rect 69296 2450 69348 2456
rect 69296 2304 69348 2310
rect 69296 2246 69348 2252
rect 69308 2106 69336 2246
rect 69296 2100 69348 2106
rect 69296 2042 69348 2048
rect 69400 800 69428 2858
rect 69584 800 69612 4082
rect 69756 3596 69808 3602
rect 69756 3538 69808 3544
rect 69768 800 69796 3538
rect 70044 3126 70072 13806
rect 70136 13326 70164 18176
rect 70320 15201 70348 33594
rect 70306 15192 70362 15201
rect 70306 15127 70362 15136
rect 70320 14958 70348 15127
rect 70308 14952 70360 14958
rect 70308 14894 70360 14900
rect 70412 14550 70440 37946
rect 70504 37346 70532 39200
rect 71424 37398 71452 39200
rect 71504 38072 71556 38078
rect 71504 38014 71556 38020
rect 71412 37392 71464 37398
rect 70504 37318 70624 37346
rect 71412 37334 71464 37340
rect 70596 36922 70624 37318
rect 70676 37256 70728 37262
rect 70676 37198 70728 37204
rect 70688 37097 70716 37198
rect 71516 37126 71544 38014
rect 71688 37324 71740 37330
rect 72252 37312 72280 39200
rect 72332 37324 72384 37330
rect 72252 37284 72332 37312
rect 71688 37266 71740 37272
rect 72332 37266 72384 37272
rect 71504 37120 71556 37126
rect 70674 37088 70730 37097
rect 71504 37062 71556 37068
rect 70674 37023 70730 37032
rect 70492 36916 70544 36922
rect 70492 36858 70544 36864
rect 70584 36916 70636 36922
rect 70584 36858 70636 36864
rect 70504 36825 70532 36858
rect 70490 36816 70546 36825
rect 70490 36751 70546 36760
rect 70584 36712 70636 36718
rect 70584 36654 70636 36660
rect 70490 36408 70546 36417
rect 70596 36378 70624 36654
rect 70490 36343 70492 36352
rect 70544 36343 70546 36352
rect 70584 36372 70636 36378
rect 70492 36314 70544 36320
rect 70584 36314 70636 36320
rect 70676 34060 70728 34066
rect 70676 34002 70728 34008
rect 70584 33992 70636 33998
rect 70584 33934 70636 33940
rect 70596 32842 70624 33934
rect 70584 32836 70636 32842
rect 70584 32778 70636 32784
rect 70688 31754 70716 34002
rect 70768 33856 70820 33862
rect 70768 33798 70820 33804
rect 70504 31726 70716 31754
rect 70780 31754 70808 33798
rect 70780 31726 70900 31754
rect 70504 22982 70532 31726
rect 70676 30796 70728 30802
rect 70676 30738 70728 30744
rect 70584 26444 70636 26450
rect 70584 26386 70636 26392
rect 70492 22976 70544 22982
rect 70492 22918 70544 22924
rect 70504 22166 70532 22918
rect 70492 22160 70544 22166
rect 70492 22102 70544 22108
rect 70596 20534 70624 26386
rect 70688 22094 70716 30738
rect 70768 30048 70820 30054
rect 70768 29990 70820 29996
rect 70780 29782 70808 29990
rect 70768 29776 70820 29782
rect 70768 29718 70820 29724
rect 70688 22066 70808 22094
rect 70584 20528 70636 20534
rect 70584 20470 70636 20476
rect 70780 20398 70808 22066
rect 70768 20392 70820 20398
rect 70768 20334 70820 20340
rect 70872 20262 70900 31726
rect 71700 30802 71728 37266
rect 73172 36922 73200 39200
rect 74000 37398 74028 39200
rect 74816 38480 74868 38486
rect 74816 38422 74868 38428
rect 74264 37732 74316 37738
rect 74264 37674 74316 37680
rect 73988 37392 74040 37398
rect 73988 37334 74040 37340
rect 74276 37330 74304 37674
rect 74264 37324 74316 37330
rect 74264 37266 74316 37272
rect 74724 37324 74776 37330
rect 74724 37266 74776 37272
rect 73252 37256 73304 37262
rect 73252 37198 73304 37204
rect 73528 37256 73580 37262
rect 73528 37198 73580 37204
rect 73264 36922 73292 37198
rect 73160 36916 73212 36922
rect 73160 36858 73212 36864
rect 73252 36916 73304 36922
rect 73252 36858 73304 36864
rect 73434 36816 73490 36825
rect 73434 36751 73490 36760
rect 72884 36644 72936 36650
rect 72884 36586 72936 36592
rect 72056 36576 72108 36582
rect 72056 36518 72108 36524
rect 72068 36417 72096 36518
rect 72054 36408 72110 36417
rect 72054 36343 72110 36352
rect 72896 36310 72924 36586
rect 73448 36582 73476 36751
rect 73436 36576 73488 36582
rect 73436 36518 73488 36524
rect 72884 36304 72936 36310
rect 72884 36246 72936 36252
rect 73540 36038 73568 37198
rect 73988 36712 74040 36718
rect 73988 36654 74040 36660
rect 73804 36576 73856 36582
rect 73804 36518 73856 36524
rect 73528 36032 73580 36038
rect 73528 35974 73580 35980
rect 73620 36032 73672 36038
rect 73620 35974 73672 35980
rect 72700 35760 72752 35766
rect 72700 35702 72752 35708
rect 72332 35148 72384 35154
rect 72332 35090 72384 35096
rect 72240 33584 72292 33590
rect 72240 33526 72292 33532
rect 71780 33040 71832 33046
rect 71780 32982 71832 32988
rect 71688 30796 71740 30802
rect 71688 30738 71740 30744
rect 71320 30388 71372 30394
rect 71320 30330 71372 30336
rect 71044 30252 71096 30258
rect 71044 30194 71096 30200
rect 71056 29306 71084 30194
rect 71332 30190 71360 30330
rect 71320 30184 71372 30190
rect 71320 30126 71372 30132
rect 71044 29300 71096 29306
rect 71044 29242 71096 29248
rect 71136 29096 71188 29102
rect 71136 29038 71188 29044
rect 71044 28960 71096 28966
rect 71044 28902 71096 28908
rect 71056 28694 71084 28902
rect 71044 28688 71096 28694
rect 71044 28630 71096 28636
rect 71044 23044 71096 23050
rect 71044 22986 71096 22992
rect 70860 20256 70912 20262
rect 70860 20198 70912 20204
rect 70688 18958 70900 18986
rect 70688 18834 70716 18958
rect 70766 18864 70822 18873
rect 70676 18828 70728 18834
rect 70766 18799 70768 18808
rect 70676 18770 70728 18776
rect 70820 18799 70822 18808
rect 70768 18770 70820 18776
rect 70780 18222 70808 18770
rect 70872 18426 70900 18958
rect 70952 18828 71004 18834
rect 71056 18816 71084 22986
rect 71148 20482 71176 29038
rect 71148 20454 71268 20482
rect 71136 20392 71188 20398
rect 71136 20334 71188 20340
rect 71148 20262 71176 20334
rect 71136 20256 71188 20262
rect 71136 20198 71188 20204
rect 71240 19718 71268 20454
rect 71228 19712 71280 19718
rect 71228 19654 71280 19660
rect 71004 18788 71084 18816
rect 71134 18864 71190 18873
rect 71134 18799 71136 18808
rect 70952 18770 71004 18776
rect 71188 18799 71190 18808
rect 71136 18770 71188 18776
rect 70860 18420 70912 18426
rect 70860 18362 70912 18368
rect 70768 18216 70820 18222
rect 70768 18158 70820 18164
rect 70768 16448 70820 16454
rect 70768 16390 70820 16396
rect 70780 15910 70808 16390
rect 70860 16176 70912 16182
rect 70860 16118 70912 16124
rect 70872 15910 70900 16118
rect 70768 15904 70820 15910
rect 70768 15846 70820 15852
rect 70860 15904 70912 15910
rect 70860 15846 70912 15852
rect 71044 14884 71096 14890
rect 71044 14826 71096 14832
rect 71056 14793 71084 14826
rect 71042 14784 71098 14793
rect 71042 14719 71098 14728
rect 70400 14544 70452 14550
rect 70400 14486 70452 14492
rect 70768 14476 70820 14482
rect 70768 14418 70820 14424
rect 70584 14272 70636 14278
rect 70584 14214 70636 14220
rect 70676 14272 70728 14278
rect 70676 14214 70728 14220
rect 70596 14074 70624 14214
rect 70584 14068 70636 14074
rect 70584 14010 70636 14016
rect 70124 13320 70176 13326
rect 70124 13262 70176 13268
rect 70216 12640 70268 12646
rect 70214 12608 70216 12617
rect 70268 12608 70270 12617
rect 70214 12543 70270 12552
rect 70124 11892 70176 11898
rect 70124 11834 70176 11840
rect 70308 11892 70360 11898
rect 70308 11834 70360 11840
rect 70032 3120 70084 3126
rect 70032 3062 70084 3068
rect 70136 3058 70164 11834
rect 70216 4140 70268 4146
rect 70216 4082 70268 4088
rect 70124 3052 70176 3058
rect 70124 2994 70176 3000
rect 70032 2100 70084 2106
rect 70032 2042 70084 2048
rect 70044 800 70072 2042
rect 70228 800 70256 4082
rect 70320 2582 70348 11834
rect 70400 3596 70452 3602
rect 70400 3538 70452 3544
rect 70308 2576 70360 2582
rect 70308 2518 70360 2524
rect 70412 800 70440 3538
rect 70584 2916 70636 2922
rect 70584 2858 70636 2864
rect 70596 800 70624 2858
rect 70688 1018 70716 14214
rect 70780 12374 70808 14418
rect 70768 12368 70820 12374
rect 70768 12310 70820 12316
rect 71228 7472 71280 7478
rect 71228 7414 71280 7420
rect 71044 5228 71096 5234
rect 71044 5170 71096 5176
rect 71056 4758 71084 5170
rect 71044 4752 71096 4758
rect 71044 4694 71096 4700
rect 70768 4684 70820 4690
rect 70768 4626 70820 4632
rect 70676 1012 70728 1018
rect 70676 954 70728 960
rect 70780 800 70808 4626
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 70860 2916 70912 2922
rect 70860 2858 70912 2864
rect 67454 504 67510 513
rect 67454 439 67510 448
rect 67546 0 67602 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70766 0 70822 800
rect 70872 66 70900 2858
rect 71056 800 71084 3538
rect 71240 2582 71268 7414
rect 71332 3670 71360 30126
rect 71412 24880 71464 24886
rect 71412 24822 71464 24828
rect 71424 22778 71452 24822
rect 71688 24132 71740 24138
rect 71688 24074 71740 24080
rect 71700 23050 71728 24074
rect 71688 23044 71740 23050
rect 71688 22986 71740 22992
rect 71412 22772 71464 22778
rect 71412 22714 71464 22720
rect 71792 20534 71820 32982
rect 72056 30864 72108 30870
rect 72056 30806 72108 30812
rect 72068 30666 72096 30806
rect 72056 30660 72108 30666
rect 72056 30602 72108 30608
rect 72068 27606 72096 30602
rect 72056 27600 72108 27606
rect 72056 27542 72108 27548
rect 72148 27464 72200 27470
rect 72148 27406 72200 27412
rect 71870 23760 71926 23769
rect 71870 23695 71872 23704
rect 71924 23695 71926 23704
rect 71872 23666 71924 23672
rect 72160 23254 72188 27406
rect 72252 23322 72280 33526
rect 72240 23316 72292 23322
rect 72240 23258 72292 23264
rect 72148 23248 72200 23254
rect 72148 23190 72200 23196
rect 72056 23180 72108 23186
rect 72056 23122 72108 23128
rect 71964 23112 72016 23118
rect 71964 23054 72016 23060
rect 71780 20528 71832 20534
rect 71780 20470 71832 20476
rect 71792 20262 71820 20470
rect 71780 20256 71832 20262
rect 71780 20198 71832 20204
rect 71688 19712 71740 19718
rect 71688 19654 71740 19660
rect 71780 19712 71832 19718
rect 71780 19654 71832 19660
rect 71700 12782 71728 19654
rect 71792 18154 71820 19654
rect 71872 19372 71924 19378
rect 71872 19314 71924 19320
rect 71780 18148 71832 18154
rect 71780 18090 71832 18096
rect 71780 14952 71832 14958
rect 71780 14894 71832 14900
rect 71792 13394 71820 14894
rect 71884 13938 71912 19314
rect 71976 17785 72004 23054
rect 71962 17776 72018 17785
rect 71962 17711 72018 17720
rect 71964 16720 72016 16726
rect 71964 16662 72016 16668
rect 71872 13932 71924 13938
rect 71872 13874 71924 13880
rect 71780 13388 71832 13394
rect 71780 13330 71832 13336
rect 71596 12776 71648 12782
rect 71596 12718 71648 12724
rect 71688 12776 71740 12782
rect 71688 12718 71740 12724
rect 71504 10532 71556 10538
rect 71504 10474 71556 10480
rect 71516 10062 71544 10474
rect 71504 10056 71556 10062
rect 71504 9998 71556 10004
rect 71608 5914 71636 12718
rect 71686 10160 71742 10169
rect 71686 10095 71742 10104
rect 71596 5908 71648 5914
rect 71596 5850 71648 5856
rect 71412 4072 71464 4078
rect 71412 4014 71464 4020
rect 71320 3664 71372 3670
rect 71320 3606 71372 3612
rect 71320 2984 71372 2990
rect 71320 2926 71372 2932
rect 71228 2576 71280 2582
rect 71228 2518 71280 2524
rect 71228 1420 71280 1426
rect 71228 1362 71280 1368
rect 71240 800 71268 1362
rect 70860 60 70912 66
rect 70860 2 70912 8
rect 71042 0 71098 800
rect 71226 0 71282 800
rect 71332 542 71360 2926
rect 71424 800 71452 4014
rect 71596 3596 71648 3602
rect 71596 3538 71648 3544
rect 71504 2984 71556 2990
rect 71504 2926 71556 2932
rect 71320 536 71372 542
rect 71320 478 71372 484
rect 71410 0 71466 800
rect 71516 610 71544 2926
rect 71608 800 71636 3538
rect 71700 2650 71728 10095
rect 71872 9376 71924 9382
rect 71872 9318 71924 9324
rect 71884 2990 71912 9318
rect 71976 6866 72004 16662
rect 72068 13938 72096 23122
rect 72240 23044 72292 23050
rect 72240 22986 72292 22992
rect 72148 21072 72200 21078
rect 72148 21014 72200 21020
rect 72160 20398 72188 21014
rect 72148 20392 72200 20398
rect 72148 20334 72200 20340
rect 72160 17746 72188 20334
rect 72148 17740 72200 17746
rect 72148 17682 72200 17688
rect 72148 17264 72200 17270
rect 72148 17206 72200 17212
rect 72056 13932 72108 13938
rect 72056 13874 72108 13880
rect 72160 6934 72188 17206
rect 72252 15706 72280 22986
rect 72240 15700 72292 15706
rect 72240 15642 72292 15648
rect 72344 11218 72372 35090
rect 72424 33992 72476 33998
rect 72424 33934 72476 33940
rect 72436 30802 72464 33934
rect 72424 30796 72476 30802
rect 72424 30738 72476 30744
rect 72436 23050 72464 30738
rect 72608 27396 72660 27402
rect 72608 27338 72660 27344
rect 72516 26376 72568 26382
rect 72514 26344 72516 26353
rect 72568 26344 72570 26353
rect 72514 26279 72570 26288
rect 72620 23186 72648 27338
rect 72712 24886 72740 35702
rect 72976 33924 73028 33930
rect 72976 33866 73028 33872
rect 72792 30796 72844 30802
rect 72792 30738 72844 30744
rect 72700 24880 72752 24886
rect 72700 24822 72752 24828
rect 72804 24750 72832 30738
rect 72988 28994 73016 33866
rect 73068 30796 73120 30802
rect 73068 30738 73120 30744
rect 72896 28966 73016 28994
rect 72896 26874 72924 28966
rect 72896 26846 73016 26874
rect 72884 26444 72936 26450
rect 72884 26386 72936 26392
rect 72792 24744 72844 24750
rect 72792 24686 72844 24692
rect 72700 24336 72752 24342
rect 72700 24278 72752 24284
rect 72792 24336 72844 24342
rect 72792 24278 72844 24284
rect 72712 23186 72740 24278
rect 72804 24206 72832 24278
rect 72792 24200 72844 24206
rect 72792 24142 72844 24148
rect 72608 23180 72660 23186
rect 72608 23122 72660 23128
rect 72700 23180 72752 23186
rect 72700 23122 72752 23128
rect 72424 23044 72476 23050
rect 72424 22986 72476 22992
rect 72700 20868 72752 20874
rect 72700 20810 72752 20816
rect 72712 20466 72740 20810
rect 72700 20460 72752 20466
rect 72700 20402 72752 20408
rect 72896 20398 72924 26386
rect 72988 20398 73016 26846
rect 73080 23662 73108 30738
rect 73632 30326 73660 35974
rect 73620 30320 73672 30326
rect 73620 30262 73672 30268
rect 73816 28014 73844 36518
rect 74000 30054 74028 36654
rect 74172 36032 74224 36038
rect 74172 35974 74224 35980
rect 74540 36032 74592 36038
rect 74540 35974 74592 35980
rect 73988 30048 74040 30054
rect 73988 29990 74040 29996
rect 74000 29102 74028 29990
rect 74078 29200 74134 29209
rect 74078 29135 74134 29144
rect 73988 29096 74040 29102
rect 73988 29038 74040 29044
rect 73804 28008 73856 28014
rect 73804 27950 73856 27956
rect 74092 26450 74120 29135
rect 73804 26444 73856 26450
rect 73724 26404 73804 26432
rect 73620 26376 73672 26382
rect 73620 26318 73672 26324
rect 73344 26308 73396 26314
rect 73344 26250 73396 26256
rect 73252 25832 73304 25838
rect 73252 25774 73304 25780
rect 73160 25220 73212 25226
rect 73160 25162 73212 25168
rect 73172 23798 73200 25162
rect 73160 23792 73212 23798
rect 73160 23734 73212 23740
rect 73068 23656 73120 23662
rect 73068 23598 73120 23604
rect 73080 20466 73108 23598
rect 73160 20528 73212 20534
rect 73160 20470 73212 20476
rect 73068 20460 73120 20466
rect 73068 20402 73120 20408
rect 72608 20392 72660 20398
rect 72884 20392 72936 20398
rect 72608 20334 72660 20340
rect 72712 20340 72884 20346
rect 72712 20334 72936 20340
rect 72976 20392 73028 20398
rect 72976 20334 73028 20340
rect 72620 19378 72648 20334
rect 72712 20318 72924 20334
rect 72608 19372 72660 19378
rect 72608 19314 72660 19320
rect 72424 18896 72476 18902
rect 72424 18838 72476 18844
rect 72436 18737 72464 18838
rect 72422 18728 72478 18737
rect 72422 18663 72478 18672
rect 72424 18148 72476 18154
rect 72424 18090 72476 18096
rect 72436 12782 72464 18090
rect 72712 16454 72740 20318
rect 72988 20210 73016 20334
rect 72804 20182 73016 20210
rect 72700 16448 72752 16454
rect 72700 16390 72752 16396
rect 72608 15904 72660 15910
rect 72608 15846 72660 15852
rect 72424 12776 72476 12782
rect 72424 12718 72476 12724
rect 72620 12306 72648 15846
rect 72700 14272 72752 14278
rect 72700 14214 72752 14220
rect 72712 14074 72740 14214
rect 72700 14068 72752 14074
rect 72700 14010 72752 14016
rect 72712 13870 72740 14010
rect 72700 13864 72752 13870
rect 72700 13806 72752 13812
rect 72804 13394 72832 20182
rect 73080 20074 73108 20402
rect 73172 20262 73200 20470
rect 73160 20256 73212 20262
rect 73160 20198 73212 20204
rect 72988 20046 73108 20074
rect 72988 19446 73016 20046
rect 73068 19984 73120 19990
rect 73068 19926 73120 19932
rect 72976 19440 73028 19446
rect 72976 19382 73028 19388
rect 72884 18828 72936 18834
rect 72884 18770 72936 18776
rect 72896 13954 72924 18770
rect 73080 18154 73108 19926
rect 73264 19310 73292 25774
rect 73356 23202 73384 26250
rect 73436 26240 73488 26246
rect 73436 26182 73488 26188
rect 73448 25974 73476 26182
rect 73436 25968 73488 25974
rect 73436 25910 73488 25916
rect 73356 23174 73568 23202
rect 73436 23112 73488 23118
rect 73436 23054 73488 23060
rect 73448 22098 73476 23054
rect 73436 22092 73488 22098
rect 73436 22034 73488 22040
rect 73252 19304 73304 19310
rect 73252 19246 73304 19252
rect 73160 18352 73212 18358
rect 73264 18340 73292 19246
rect 73212 18312 73292 18340
rect 73344 18352 73396 18358
rect 73160 18294 73212 18300
rect 73344 18294 73396 18300
rect 73068 18148 73120 18154
rect 73068 18090 73120 18096
rect 72976 17264 73028 17270
rect 72976 17206 73028 17212
rect 72988 16658 73016 17206
rect 72976 16652 73028 16658
rect 72976 16594 73028 16600
rect 72896 13926 73016 13954
rect 72884 13864 72936 13870
rect 72884 13806 72936 13812
rect 72792 13388 72844 13394
rect 72792 13330 72844 13336
rect 72608 12300 72660 12306
rect 72608 12242 72660 12248
rect 72332 11212 72384 11218
rect 72332 11154 72384 11160
rect 72148 6928 72200 6934
rect 72148 6870 72200 6876
rect 71964 6860 72016 6866
rect 71964 6802 72016 6808
rect 72608 6860 72660 6866
rect 72608 6802 72660 6808
rect 72620 6662 72648 6802
rect 72608 6656 72660 6662
rect 72608 6598 72660 6604
rect 72896 6458 72924 13806
rect 72988 13394 73016 13926
rect 72976 13388 73028 13394
rect 72976 13330 73028 13336
rect 73080 12434 73108 18090
rect 73356 16114 73384 18294
rect 73344 16108 73396 16114
rect 73344 16050 73396 16056
rect 73448 14890 73476 22034
rect 73436 14884 73488 14890
rect 73436 14826 73488 14832
rect 72988 12406 73108 12434
rect 72988 9586 73016 12406
rect 73068 9716 73120 9722
rect 73068 9658 73120 9664
rect 72976 9580 73028 9586
rect 72976 9522 73028 9528
rect 73080 7886 73108 9658
rect 73068 7880 73120 7886
rect 73068 7822 73120 7828
rect 72884 6452 72936 6458
rect 72884 6394 72936 6400
rect 72056 4072 72108 4078
rect 72056 4014 72108 4020
rect 72608 4072 72660 4078
rect 72608 4014 72660 4020
rect 73252 4072 73304 4078
rect 73252 4014 73304 4020
rect 71872 2984 71924 2990
rect 71872 2926 71924 2932
rect 71964 2848 72016 2854
rect 71964 2790 72016 2796
rect 71688 2644 71740 2650
rect 71688 2586 71740 2592
rect 71976 2553 72004 2790
rect 71962 2544 72018 2553
rect 71780 2508 71832 2514
rect 71780 2450 71832 2456
rect 71872 2508 71924 2514
rect 71962 2479 72018 2488
rect 71872 2450 71924 2456
rect 71688 2440 71740 2446
rect 71688 2382 71740 2388
rect 71700 2106 71728 2382
rect 71688 2100 71740 2106
rect 71688 2042 71740 2048
rect 71792 1970 71820 2450
rect 71780 1964 71832 1970
rect 71780 1906 71832 1912
rect 71884 1170 71912 2450
rect 71792 1142 71912 1170
rect 71792 800 71820 1142
rect 72068 800 72096 4014
rect 72240 2984 72292 2990
rect 72240 2926 72292 2932
rect 72148 2508 72200 2514
rect 72148 2450 72200 2456
rect 72160 2310 72188 2450
rect 72148 2304 72200 2310
rect 72148 2246 72200 2252
rect 72160 1222 72188 2246
rect 72148 1216 72200 1222
rect 72148 1158 72200 1164
rect 72252 800 72280 2926
rect 72424 2848 72476 2854
rect 72424 2790 72476 2796
rect 72330 2544 72386 2553
rect 72330 2479 72386 2488
rect 71504 604 71556 610
rect 71504 546 71556 552
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72344 474 72372 2479
rect 72436 800 72464 2790
rect 72516 2304 72568 2310
rect 72516 2246 72568 2252
rect 72528 2038 72556 2246
rect 72516 2032 72568 2038
rect 72516 1974 72568 1980
rect 72620 800 72648 4014
rect 72792 3596 72844 3602
rect 72792 3538 72844 3544
rect 72700 2372 72752 2378
rect 72700 2314 72752 2320
rect 72712 2038 72740 2314
rect 72700 2032 72752 2038
rect 72700 1974 72752 1980
rect 72804 800 72832 3538
rect 72884 2372 72936 2378
rect 72884 2314 72936 2320
rect 72896 1426 72924 2314
rect 73068 2304 73120 2310
rect 73068 2246 73120 2252
rect 72884 1420 72936 1426
rect 72884 1362 72936 1368
rect 73080 800 73108 2246
rect 73264 800 73292 4014
rect 73436 2984 73488 2990
rect 73436 2926 73488 2932
rect 73448 800 73476 2926
rect 73540 814 73568 23174
rect 73632 15434 73660 26318
rect 73724 21078 73752 26404
rect 73804 26386 73856 26392
rect 74080 26444 74132 26450
rect 74080 26386 74132 26392
rect 73988 26376 74040 26382
rect 73988 26318 74040 26324
rect 74000 25838 74028 26318
rect 73988 25832 74040 25838
rect 73988 25774 74040 25780
rect 74184 25401 74212 35974
rect 74448 30592 74500 30598
rect 74448 30534 74500 30540
rect 74356 28008 74408 28014
rect 74356 27950 74408 27956
rect 74264 27668 74316 27674
rect 74264 27610 74316 27616
rect 74276 26246 74304 27610
rect 74368 27334 74396 27950
rect 74356 27328 74408 27334
rect 74356 27270 74408 27276
rect 74356 26376 74408 26382
rect 74354 26344 74356 26353
rect 74408 26344 74410 26353
rect 74354 26279 74410 26288
rect 74264 26240 74316 26246
rect 74264 26182 74316 26188
rect 74170 25392 74226 25401
rect 74170 25327 74226 25336
rect 74356 25288 74408 25294
rect 74356 25230 74408 25236
rect 74368 23118 74396 25230
rect 74460 23594 74488 30534
rect 74448 23588 74500 23594
rect 74448 23530 74500 23536
rect 74356 23112 74408 23118
rect 74356 23054 74408 23060
rect 74448 22976 74500 22982
rect 74448 22918 74500 22924
rect 73804 22704 73856 22710
rect 73804 22646 73856 22652
rect 73712 21072 73764 21078
rect 73712 21014 73764 21020
rect 73712 18284 73764 18290
rect 73712 18226 73764 18232
rect 73620 15428 73672 15434
rect 73620 15370 73672 15376
rect 73620 1420 73672 1426
rect 73620 1362 73672 1368
rect 73528 808 73580 814
rect 72332 468 72384 474
rect 72332 410 72384 416
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73250 0 73306 800
rect 73434 0 73490 800
rect 73632 800 73660 1362
rect 73528 750 73580 756
rect 73618 0 73674 800
rect 73724 202 73752 18226
rect 73816 16046 73844 22646
rect 74460 22642 74488 22918
rect 74448 22636 74500 22642
rect 74448 22578 74500 22584
rect 73988 19916 74040 19922
rect 73988 19858 74040 19864
rect 74000 19514 74028 19858
rect 73988 19508 74040 19514
rect 73988 19450 74040 19456
rect 74264 17672 74316 17678
rect 74264 17614 74316 17620
rect 73804 16040 73856 16046
rect 73804 15982 73856 15988
rect 73896 11212 73948 11218
rect 73896 11154 73948 11160
rect 73908 9450 73936 11154
rect 73896 9444 73948 9450
rect 73896 9386 73948 9392
rect 73908 5914 73936 9386
rect 74276 9178 74304 17614
rect 74264 9172 74316 9178
rect 74264 9114 74316 9120
rect 74172 8968 74224 8974
rect 74172 8910 74224 8916
rect 74080 8288 74132 8294
rect 74080 8230 74132 8236
rect 73896 5908 73948 5914
rect 73896 5850 73948 5856
rect 74092 5778 74120 8230
rect 74184 7449 74212 8910
rect 74170 7440 74226 7449
rect 74170 7375 74226 7384
rect 74552 6769 74580 35974
rect 74736 28966 74764 37266
rect 74724 28960 74776 28966
rect 74724 28902 74776 28908
rect 74736 27878 74764 28902
rect 74724 27872 74776 27878
rect 74724 27814 74776 27820
rect 74632 26308 74684 26314
rect 74632 26250 74684 26256
rect 74644 24682 74672 26250
rect 74632 24676 74684 24682
rect 74632 24618 74684 24624
rect 74722 24168 74778 24177
rect 74722 24103 74724 24112
rect 74776 24103 74778 24112
rect 74724 24074 74776 24080
rect 74632 22568 74684 22574
rect 74632 22510 74684 22516
rect 74644 19922 74672 22510
rect 74632 19916 74684 19922
rect 74632 19858 74684 19864
rect 74538 6760 74594 6769
rect 74538 6695 74594 6704
rect 74080 5772 74132 5778
rect 74080 5714 74132 5720
rect 73988 5568 74040 5574
rect 73988 5510 74040 5516
rect 74000 5370 74028 5510
rect 74092 5370 74120 5714
rect 73988 5364 74040 5370
rect 73988 5306 74040 5312
rect 74080 5364 74132 5370
rect 74080 5306 74132 5312
rect 73804 4684 73856 4690
rect 73804 4626 73856 4632
rect 73816 800 73844 4626
rect 74172 4480 74224 4486
rect 74172 4422 74224 4428
rect 74080 3596 74132 3602
rect 74080 3538 74132 3544
rect 74092 800 74120 3538
rect 74184 2650 74212 4422
rect 74448 4072 74500 4078
rect 74448 4014 74500 4020
rect 74172 2644 74224 2650
rect 74172 2586 74224 2592
rect 74264 1488 74316 1494
rect 74264 1430 74316 1436
rect 74276 800 74304 1430
rect 74460 800 74488 4014
rect 74632 3596 74684 3602
rect 74632 3538 74684 3544
rect 74540 3392 74592 3398
rect 74540 3334 74592 3340
rect 74552 3194 74580 3334
rect 74540 3188 74592 3194
rect 74540 3130 74592 3136
rect 74644 800 74672 3538
rect 74828 3194 74856 38422
rect 74920 37330 74948 39200
rect 75736 38412 75788 38418
rect 75736 38354 75788 38360
rect 75368 37800 75420 37806
rect 75368 37742 75420 37748
rect 74908 37324 74960 37330
rect 74908 37266 74960 37272
rect 75274 36272 75330 36281
rect 75274 36207 75330 36216
rect 75184 34536 75236 34542
rect 75184 34478 75236 34484
rect 75092 27056 75144 27062
rect 75092 26998 75144 27004
rect 75104 26450 75132 26998
rect 75092 26444 75144 26450
rect 75092 26386 75144 26392
rect 75090 24440 75146 24449
rect 75000 24404 75052 24410
rect 75090 24375 75146 24384
rect 75000 24346 75052 24352
rect 75012 23526 75040 24346
rect 75104 24274 75132 24375
rect 75092 24268 75144 24274
rect 75092 24210 75144 24216
rect 75092 24132 75144 24138
rect 75092 24074 75144 24080
rect 75104 23662 75132 24074
rect 75092 23656 75144 23662
rect 75092 23598 75144 23604
rect 75000 23520 75052 23526
rect 75000 23462 75052 23468
rect 75196 22094 75224 34478
rect 75104 22066 75224 22094
rect 75104 15162 75132 22066
rect 75184 17604 75236 17610
rect 75184 17546 75236 17552
rect 75196 17338 75224 17546
rect 75184 17332 75236 17338
rect 75184 17274 75236 17280
rect 75092 15156 75144 15162
rect 75092 15098 75144 15104
rect 75288 12434 75316 36207
rect 75380 22098 75408 37742
rect 75460 37732 75512 37738
rect 75460 37674 75512 37680
rect 75472 30870 75500 37674
rect 75552 34536 75604 34542
rect 75552 34478 75604 34484
rect 75564 33930 75592 34478
rect 75552 33924 75604 33930
rect 75552 33866 75604 33872
rect 75460 30864 75512 30870
rect 75460 30806 75512 30812
rect 75472 23526 75500 30806
rect 75552 26920 75604 26926
rect 75552 26862 75604 26868
rect 75460 23520 75512 23526
rect 75460 23462 75512 23468
rect 75460 23316 75512 23322
rect 75460 23258 75512 23264
rect 75472 22642 75500 23258
rect 75460 22636 75512 22642
rect 75460 22578 75512 22584
rect 75368 22092 75420 22098
rect 75472 22094 75500 22578
rect 75564 22574 75592 26862
rect 75644 24676 75696 24682
rect 75644 24618 75696 24624
rect 75552 22568 75604 22574
rect 75552 22510 75604 22516
rect 75472 22066 75592 22094
rect 75368 22034 75420 22040
rect 75368 14544 75420 14550
rect 75368 14486 75420 14492
rect 75380 14414 75408 14486
rect 75368 14408 75420 14414
rect 75368 14350 75420 14356
rect 75368 13456 75420 13462
rect 75368 13398 75420 13404
rect 75380 12986 75408 13398
rect 75368 12980 75420 12986
rect 75368 12922 75420 12928
rect 75460 12980 75512 12986
rect 75460 12922 75512 12928
rect 75472 12782 75500 12922
rect 75460 12776 75512 12782
rect 75460 12718 75512 12724
rect 75460 12640 75512 12646
rect 75460 12582 75512 12588
rect 75288 12406 75408 12434
rect 75092 10600 75144 10606
rect 75092 10542 75144 10548
rect 75104 10130 75132 10542
rect 75276 10532 75328 10538
rect 75276 10474 75328 10480
rect 75184 10464 75236 10470
rect 75184 10406 75236 10412
rect 75196 10266 75224 10406
rect 75184 10260 75236 10266
rect 75184 10202 75236 10208
rect 75092 10124 75144 10130
rect 75092 10066 75144 10072
rect 75288 9994 75316 10474
rect 75276 9988 75328 9994
rect 75276 9930 75328 9936
rect 75092 4072 75144 4078
rect 75092 4014 75144 4020
rect 74908 3528 74960 3534
rect 74908 3470 74960 3476
rect 74816 3188 74868 3194
rect 74816 3130 74868 3136
rect 74828 2990 74856 3130
rect 74920 3058 74948 3470
rect 74908 3052 74960 3058
rect 74908 2994 74960 3000
rect 74816 2984 74868 2990
rect 74816 2926 74868 2932
rect 74908 2916 74960 2922
rect 74908 2858 74960 2864
rect 74724 2644 74776 2650
rect 74724 2586 74776 2592
rect 74736 1494 74764 2586
rect 74724 1488 74776 1494
rect 74724 1430 74776 1436
rect 74920 800 74948 2858
rect 75000 2440 75052 2446
rect 75000 2382 75052 2388
rect 75012 1426 75040 2382
rect 75000 1420 75052 1426
rect 75000 1362 75052 1368
rect 75104 800 75132 4014
rect 75276 2984 75328 2990
rect 75276 2926 75328 2932
rect 75288 800 75316 2926
rect 75380 2582 75408 12406
rect 75472 12374 75500 12582
rect 75460 12368 75512 12374
rect 75460 12310 75512 12316
rect 75472 11558 75500 12310
rect 75564 11762 75592 22066
rect 75656 21010 75684 24618
rect 75748 24313 75776 38354
rect 75840 36718 75868 39200
rect 76288 38888 76340 38894
rect 76288 38830 76340 38836
rect 76196 37256 76248 37262
rect 76196 37198 76248 37204
rect 76102 36952 76158 36961
rect 76102 36887 76158 36896
rect 75828 36712 75880 36718
rect 75828 36654 75880 36660
rect 75920 36644 75972 36650
rect 75920 36586 75972 36592
rect 75932 36106 75960 36586
rect 76012 36372 76064 36378
rect 76012 36314 76064 36320
rect 75920 36100 75972 36106
rect 75920 36042 75972 36048
rect 76024 35562 76052 36314
rect 76012 35556 76064 35562
rect 76012 35498 76064 35504
rect 76116 31754 76144 36887
rect 76208 36718 76236 37198
rect 76196 36712 76248 36718
rect 76196 36654 76248 36660
rect 76300 34950 76328 38830
rect 76668 37398 76696 39200
rect 76932 37664 76984 37670
rect 76932 37606 76984 37612
rect 76656 37392 76708 37398
rect 76840 37392 76892 37398
rect 76656 37334 76708 37340
rect 76838 37360 76840 37369
rect 76892 37360 76894 37369
rect 76838 37295 76894 37304
rect 76944 37262 76972 37606
rect 77588 37466 77616 39200
rect 77576 37460 77628 37466
rect 77576 37402 77628 37408
rect 77484 37324 77536 37330
rect 77484 37266 77536 37272
rect 76932 37256 76984 37262
rect 76932 37198 76984 37204
rect 76288 34944 76340 34950
rect 76288 34886 76340 34892
rect 77208 34944 77260 34950
rect 77208 34886 77260 34892
rect 76116 31726 76236 31754
rect 75920 25968 75972 25974
rect 75920 25910 75972 25916
rect 75828 24880 75880 24886
rect 75828 24822 75880 24828
rect 75840 24342 75868 24822
rect 75828 24336 75880 24342
rect 75734 24304 75790 24313
rect 75828 24278 75880 24284
rect 75734 24239 75736 24248
rect 75788 24239 75790 24248
rect 75736 24210 75788 24216
rect 75748 24179 75776 24210
rect 75840 24120 75868 24278
rect 75932 24274 75960 25910
rect 75920 24268 75972 24274
rect 75920 24210 75972 24216
rect 75748 24092 75868 24120
rect 75644 21004 75696 21010
rect 75644 20946 75696 20952
rect 75644 19916 75696 19922
rect 75644 19858 75696 19864
rect 75552 11756 75604 11762
rect 75552 11698 75604 11704
rect 75460 11552 75512 11558
rect 75460 11494 75512 11500
rect 75656 6225 75684 19858
rect 75748 19718 75776 24092
rect 76012 24064 76064 24070
rect 76012 24006 76064 24012
rect 76024 23848 76052 24006
rect 76104 23860 76156 23866
rect 76024 23820 76104 23848
rect 76104 23802 76156 23808
rect 76012 23520 76064 23526
rect 76012 23462 76064 23468
rect 75920 22092 75972 22098
rect 75920 22034 75972 22040
rect 75828 19916 75880 19922
rect 75828 19858 75880 19864
rect 75736 19712 75788 19718
rect 75736 19654 75788 19660
rect 75736 13320 75788 13326
rect 75736 13262 75788 13268
rect 75748 12714 75776 13262
rect 75736 12708 75788 12714
rect 75736 12650 75788 12656
rect 75642 6216 75698 6225
rect 75642 6151 75698 6160
rect 75840 4162 75868 19858
rect 75932 19174 75960 22034
rect 76024 22030 76052 23462
rect 76104 22568 76156 22574
rect 76104 22510 76156 22516
rect 76012 22024 76064 22030
rect 76012 21966 76064 21972
rect 75920 19168 75972 19174
rect 75920 19110 75972 19116
rect 76116 18970 76144 22510
rect 76104 18964 76156 18970
rect 76104 18906 76156 18912
rect 75920 15904 75972 15910
rect 75920 15846 75972 15852
rect 75932 15570 75960 15846
rect 75920 15564 75972 15570
rect 75920 15506 75972 15512
rect 76208 14074 76236 31726
rect 76748 27600 76800 27606
rect 76748 27542 76800 27548
rect 76472 25424 76524 25430
rect 76472 25366 76524 25372
rect 76378 24440 76434 24449
rect 76378 24375 76434 24384
rect 76286 24304 76342 24313
rect 76286 24239 76342 24248
rect 76300 24206 76328 24239
rect 76392 24206 76420 24375
rect 76288 24200 76340 24206
rect 76288 24142 76340 24148
rect 76380 24200 76432 24206
rect 76380 24142 76432 24148
rect 76288 24064 76340 24070
rect 76288 24006 76340 24012
rect 76300 23769 76328 24006
rect 76380 23792 76432 23798
rect 76286 23760 76342 23769
rect 76380 23734 76432 23740
rect 76286 23695 76342 23704
rect 76392 23322 76420 23734
rect 76380 23316 76432 23322
rect 76380 23258 76432 23264
rect 76484 22094 76512 25366
rect 76564 23588 76616 23594
rect 76564 23530 76616 23536
rect 76300 22066 76512 22094
rect 76300 19854 76328 22066
rect 76288 19848 76340 19854
rect 76288 19790 76340 19796
rect 76300 18630 76328 19790
rect 76288 18624 76340 18630
rect 76288 18566 76340 18572
rect 76196 14068 76248 14074
rect 76196 14010 76248 14016
rect 75920 12640 75972 12646
rect 75918 12608 75920 12617
rect 75972 12608 75974 12617
rect 75918 12543 75974 12552
rect 76576 5574 76604 23530
rect 76760 23322 76788 27542
rect 77024 26852 77076 26858
rect 77024 26794 77076 26800
rect 77036 26761 77064 26794
rect 77022 26752 77078 26761
rect 77022 26687 77078 26696
rect 77220 23662 77248 34886
rect 77392 26920 77444 26926
rect 77390 26888 77392 26897
rect 77444 26888 77446 26897
rect 77390 26823 77446 26832
rect 77496 26042 77524 37266
rect 78416 36802 78444 39200
rect 79048 37732 79100 37738
rect 79048 37674 79100 37680
rect 79060 37330 79088 37674
rect 79048 37324 79100 37330
rect 79048 37266 79100 37272
rect 78416 36774 78720 36802
rect 78692 36718 78720 36774
rect 79336 36718 79364 39200
rect 80164 37466 80192 39200
rect 81084 38162 81112 39200
rect 81084 38134 81388 38162
rect 80244 37664 80296 37670
rect 80244 37606 80296 37612
rect 80152 37460 80204 37466
rect 80152 37402 80204 37408
rect 80256 37330 80284 37606
rect 81020 37564 81316 37584
rect 81076 37562 81100 37564
rect 81156 37562 81180 37564
rect 81236 37562 81260 37564
rect 81098 37510 81100 37562
rect 81162 37510 81174 37562
rect 81236 37510 81238 37562
rect 81076 37508 81100 37510
rect 81156 37508 81180 37510
rect 81236 37508 81260 37510
rect 81020 37488 81316 37508
rect 81360 37466 81388 38134
rect 81808 37732 81860 37738
rect 81808 37674 81860 37680
rect 81348 37460 81400 37466
rect 81348 37402 81400 37408
rect 81820 37398 81848 37674
rect 81912 37398 81940 39200
rect 81992 38276 82044 38282
rect 81992 38218 82044 38224
rect 81808 37392 81860 37398
rect 81808 37334 81860 37340
rect 81900 37392 81952 37398
rect 81900 37334 81952 37340
rect 80244 37324 80296 37330
rect 80244 37266 80296 37272
rect 81440 37324 81492 37330
rect 81440 37266 81492 37272
rect 78680 36712 78732 36718
rect 78680 36654 78732 36660
rect 79324 36712 79376 36718
rect 79324 36654 79376 36660
rect 79416 36576 79468 36582
rect 79416 36518 79468 36524
rect 79140 35828 79192 35834
rect 79140 35770 79192 35776
rect 78864 35148 78916 35154
rect 78864 35090 78916 35096
rect 77760 34060 77812 34066
rect 77760 34002 77812 34008
rect 77852 34060 77904 34066
rect 77852 34002 77904 34008
rect 77668 27056 77720 27062
rect 77668 26998 77720 27004
rect 77484 26036 77536 26042
rect 77484 25978 77536 25984
rect 77116 23656 77168 23662
rect 77116 23598 77168 23604
rect 77208 23656 77260 23662
rect 77208 23598 77260 23604
rect 76748 23316 76800 23322
rect 76748 23258 76800 23264
rect 76656 23248 76708 23254
rect 76656 23190 76708 23196
rect 76668 20874 76696 23190
rect 76656 20868 76708 20874
rect 76656 20810 76708 20816
rect 77128 15910 77156 23598
rect 77576 18216 77628 18222
rect 77576 18158 77628 18164
rect 77116 15904 77168 15910
rect 77116 15846 77168 15852
rect 77300 15700 77352 15706
rect 77300 15642 77352 15648
rect 77312 15094 77340 15642
rect 77300 15088 77352 15094
rect 77300 15030 77352 15036
rect 77392 7744 77444 7750
rect 77392 7686 77444 7692
rect 76564 5568 76616 5574
rect 76564 5510 76616 5516
rect 76932 5160 76984 5166
rect 76932 5102 76984 5108
rect 76288 4684 76340 4690
rect 76288 4626 76340 4632
rect 75564 4134 75868 4162
rect 75368 2576 75420 2582
rect 75368 2518 75420 2524
rect 75460 2372 75512 2378
rect 75460 2314 75512 2320
rect 75472 800 75500 2314
rect 73712 196 73764 202
rect 73712 138 73764 144
rect 73802 0 73858 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74906 0 74962 800
rect 75090 0 75146 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75564 241 75592 4134
rect 75736 4072 75788 4078
rect 75736 4014 75788 4020
rect 75748 2774 75776 4014
rect 75920 3596 75972 3602
rect 75920 3538 75972 3544
rect 75656 2746 75776 2774
rect 75656 800 75684 2746
rect 75932 800 75960 3538
rect 76104 2576 76156 2582
rect 76104 2518 76156 2524
rect 76116 800 76144 2518
rect 76300 800 76328 4626
rect 76380 3732 76432 3738
rect 76380 3674 76432 3680
rect 76392 3194 76420 3674
rect 76472 3596 76524 3602
rect 76472 3538 76524 3544
rect 76380 3188 76432 3194
rect 76380 3130 76432 3136
rect 76380 2508 76432 2514
rect 76380 2450 76432 2456
rect 76392 2106 76420 2450
rect 76380 2100 76432 2106
rect 76380 2042 76432 2048
rect 76484 800 76512 3538
rect 76656 2916 76708 2922
rect 76656 2858 76708 2864
rect 76564 2508 76616 2514
rect 76564 2450 76616 2456
rect 76576 1902 76604 2450
rect 76564 1896 76616 1902
rect 76564 1838 76616 1844
rect 76668 800 76696 2858
rect 76944 800 76972 5102
rect 77116 4072 77168 4078
rect 77116 4014 77168 4020
rect 77128 800 77156 4014
rect 77300 1420 77352 1426
rect 77300 1362 77352 1368
rect 77312 800 77340 1362
rect 75550 232 75606 241
rect 75550 167 75606 176
rect 75642 0 75698 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76286 0 76342 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77404 377 77432 7686
rect 77484 5160 77536 5166
rect 77484 5102 77536 5108
rect 77496 800 77524 5102
rect 77588 2990 77616 18158
rect 77680 7562 77708 26998
rect 77772 7750 77800 34002
rect 77864 32502 77892 34002
rect 77852 32496 77904 32502
rect 77852 32438 77904 32444
rect 78876 32366 78904 35090
rect 78864 32360 78916 32366
rect 78864 32302 78916 32308
rect 79048 29164 79100 29170
rect 79048 29106 79100 29112
rect 78956 28620 79008 28626
rect 78956 28562 79008 28568
rect 78404 28484 78456 28490
rect 78404 28426 78456 28432
rect 78680 28484 78732 28490
rect 78680 28426 78732 28432
rect 78312 27464 78364 27470
rect 78312 27406 78364 27412
rect 78220 27056 78272 27062
rect 78220 26998 78272 27004
rect 78232 26926 78260 26998
rect 78220 26920 78272 26926
rect 78220 26862 78272 26868
rect 78128 26784 78180 26790
rect 78126 26752 78128 26761
rect 78180 26752 78182 26761
rect 78126 26687 78182 26696
rect 78324 24750 78352 27406
rect 78312 24744 78364 24750
rect 78312 24686 78364 24692
rect 78324 24274 78352 24686
rect 78312 24268 78364 24274
rect 78312 24210 78364 24216
rect 77944 21616 77996 21622
rect 77944 21558 77996 21564
rect 77956 17338 77984 21558
rect 78048 21554 78168 21570
rect 78036 21548 78180 21554
rect 78088 21542 78128 21548
rect 78036 21490 78088 21496
rect 78128 21490 78180 21496
rect 78036 20936 78088 20942
rect 78036 20878 78088 20884
rect 78048 17338 78076 20878
rect 78140 18834 78352 18850
rect 78128 18828 78352 18834
rect 78180 18822 78352 18828
rect 78128 18770 78180 18776
rect 78324 18698 78352 18822
rect 78220 18692 78272 18698
rect 78220 18634 78272 18640
rect 78312 18692 78364 18698
rect 78312 18634 78364 18640
rect 77944 17332 77996 17338
rect 77944 17274 77996 17280
rect 78036 17332 78088 17338
rect 78036 17274 78088 17280
rect 78048 17134 78076 17274
rect 78232 17134 78260 18634
rect 78416 18086 78444 28426
rect 78494 26888 78550 26897
rect 78494 26823 78496 26832
rect 78548 26823 78550 26832
rect 78496 26794 78548 26800
rect 78496 24268 78548 24274
rect 78496 24210 78548 24216
rect 78508 24177 78536 24210
rect 78494 24168 78550 24177
rect 78494 24103 78550 24112
rect 78692 20058 78720 28426
rect 78772 23656 78824 23662
rect 78772 23598 78824 23604
rect 78784 22982 78812 23598
rect 78772 22976 78824 22982
rect 78772 22918 78824 22924
rect 78680 20052 78732 20058
rect 78680 19994 78732 20000
rect 78404 18080 78456 18086
rect 78404 18022 78456 18028
rect 78036 17128 78088 17134
rect 78036 17070 78088 17076
rect 78220 17128 78272 17134
rect 78220 17070 78272 17076
rect 78312 17128 78364 17134
rect 78312 17070 78364 17076
rect 78220 15700 78272 15706
rect 78220 15642 78272 15648
rect 77944 10600 77996 10606
rect 77944 10542 77996 10548
rect 77760 7744 77812 7750
rect 77760 7686 77812 7692
rect 77852 7744 77904 7750
rect 77852 7686 77904 7692
rect 77680 7534 77800 7562
rect 77668 3596 77720 3602
rect 77668 3538 77720 3544
rect 77576 2984 77628 2990
rect 77576 2926 77628 2932
rect 77680 800 77708 3538
rect 77772 921 77800 7534
rect 77864 7478 77892 7686
rect 77852 7472 77904 7478
rect 77852 7414 77904 7420
rect 77956 7290 77984 10542
rect 77864 7262 77984 7290
rect 77864 2582 77892 7262
rect 77944 7200 77996 7206
rect 77944 7142 77996 7148
rect 77956 4690 77984 7142
rect 78232 4758 78260 15642
rect 78324 6458 78352 17070
rect 78416 6866 78444 18022
rect 78772 17672 78824 17678
rect 78772 17614 78824 17620
rect 78784 17270 78812 17614
rect 78772 17264 78824 17270
rect 78772 17206 78824 17212
rect 78496 17128 78548 17134
rect 78496 17070 78548 17076
rect 78508 16726 78536 17070
rect 78496 16720 78548 16726
rect 78496 16662 78548 16668
rect 78496 15156 78548 15162
rect 78496 15098 78548 15104
rect 78404 6860 78456 6866
rect 78404 6802 78456 6808
rect 78312 6452 78364 6458
rect 78312 6394 78364 6400
rect 78404 4820 78456 4826
rect 78404 4762 78456 4768
rect 78220 4752 78272 4758
rect 78220 4694 78272 4700
rect 77944 4684 77996 4690
rect 77944 4626 77996 4632
rect 78416 4554 78444 4762
rect 78404 4548 78456 4554
rect 78404 4490 78456 4496
rect 78312 4072 78364 4078
rect 78312 4014 78364 4020
rect 78128 3732 78180 3738
rect 78128 3674 78180 3680
rect 78036 3392 78088 3398
rect 78036 3334 78088 3340
rect 77944 2848 77996 2854
rect 77944 2790 77996 2796
rect 77852 2576 77904 2582
rect 77852 2518 77904 2524
rect 77758 912 77814 921
rect 77758 847 77814 856
rect 77956 800 77984 2790
rect 77390 368 77446 377
rect 77390 303 77446 312
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78048 678 78076 3334
rect 78140 800 78168 3674
rect 78324 800 78352 4014
rect 78508 3194 78536 15098
rect 78680 9580 78732 9586
rect 78680 9522 78732 9528
rect 78692 7546 78720 9522
rect 78968 8634 78996 28562
rect 79060 28490 79088 29106
rect 79048 28484 79100 28490
rect 79048 28426 79100 28432
rect 79152 22094 79180 35770
rect 79324 27464 79376 27470
rect 79324 27406 79376 27412
rect 79336 27062 79364 27406
rect 79324 27056 79376 27062
rect 79324 26998 79376 27004
rect 79428 26790 79456 36518
rect 81020 36476 81316 36496
rect 81076 36474 81100 36476
rect 81156 36474 81180 36476
rect 81236 36474 81260 36476
rect 81098 36422 81100 36474
rect 81162 36422 81174 36474
rect 81236 36422 81238 36474
rect 81076 36420 81100 36422
rect 81156 36420 81180 36422
rect 81236 36420 81260 36422
rect 81020 36400 81316 36420
rect 81020 35388 81316 35408
rect 81076 35386 81100 35388
rect 81156 35386 81180 35388
rect 81236 35386 81260 35388
rect 81098 35334 81100 35386
rect 81162 35334 81174 35386
rect 81236 35334 81238 35386
rect 81076 35332 81100 35334
rect 81156 35332 81180 35334
rect 81236 35332 81260 35334
rect 81020 35312 81316 35332
rect 81020 34300 81316 34320
rect 81076 34298 81100 34300
rect 81156 34298 81180 34300
rect 81236 34298 81260 34300
rect 81098 34246 81100 34298
rect 81162 34246 81174 34298
rect 81236 34246 81238 34298
rect 81076 34244 81100 34246
rect 81156 34244 81180 34246
rect 81236 34244 81260 34246
rect 81020 34224 81316 34244
rect 81020 33212 81316 33232
rect 81076 33210 81100 33212
rect 81156 33210 81180 33212
rect 81236 33210 81260 33212
rect 81098 33158 81100 33210
rect 81162 33158 81174 33210
rect 81236 33158 81238 33210
rect 81076 33156 81100 33158
rect 81156 33156 81180 33158
rect 81236 33156 81260 33158
rect 81020 33136 81316 33156
rect 79692 32360 79744 32366
rect 79692 32302 79744 32308
rect 79600 29028 79652 29034
rect 79600 28970 79652 28976
rect 79506 28520 79562 28529
rect 79506 28455 79562 28464
rect 79416 26784 79468 26790
rect 79416 26726 79468 26732
rect 79152 22066 79456 22094
rect 79046 20360 79102 20369
rect 79046 20295 79048 20304
rect 79100 20295 79102 20304
rect 79048 20266 79100 20272
rect 79428 12434 79456 22066
rect 79336 12406 79456 12434
rect 78956 8628 79008 8634
rect 78956 8570 79008 8576
rect 78680 7540 78732 7546
rect 78680 7482 78732 7488
rect 78680 4684 78732 4690
rect 78680 4626 78732 4632
rect 78772 4684 78824 4690
rect 78772 4626 78824 4632
rect 78692 3738 78720 4626
rect 78680 3732 78732 3738
rect 78680 3674 78732 3680
rect 78588 3664 78640 3670
rect 78588 3606 78640 3612
rect 78600 3194 78628 3606
rect 78496 3188 78548 3194
rect 78496 3130 78548 3136
rect 78588 3188 78640 3194
rect 78588 3130 78640 3136
rect 78496 2984 78548 2990
rect 78496 2926 78548 2932
rect 78508 800 78536 2926
rect 78680 2304 78732 2310
rect 78680 2246 78732 2252
rect 78692 2038 78720 2246
rect 78680 2032 78732 2038
rect 78680 1974 78732 1980
rect 78784 800 78812 4626
rect 78968 4622 78996 8570
rect 78956 4616 79008 4622
rect 78956 4558 79008 4564
rect 78956 4072 79008 4078
rect 78956 4014 79008 4020
rect 78968 800 78996 4014
rect 79336 3738 79364 12406
rect 79416 4684 79468 4690
rect 79416 4626 79468 4632
rect 79324 3732 79376 3738
rect 79324 3674 79376 3680
rect 79140 3460 79192 3466
rect 79140 3402 79192 3408
rect 79152 800 79180 3402
rect 79428 2774 79456 4626
rect 79336 2746 79456 2774
rect 79232 2508 79284 2514
rect 79232 2450 79284 2456
rect 79244 1426 79272 2450
rect 79232 1420 79284 1426
rect 79232 1362 79284 1368
rect 79336 800 79364 2746
rect 79520 2650 79548 28455
rect 79612 27470 79640 28970
rect 79600 27464 79652 27470
rect 79600 27406 79652 27412
rect 79704 17218 79732 32302
rect 81020 32124 81316 32144
rect 81076 32122 81100 32124
rect 81156 32122 81180 32124
rect 81236 32122 81260 32124
rect 81098 32070 81100 32122
rect 81162 32070 81174 32122
rect 81236 32070 81238 32122
rect 81076 32068 81100 32070
rect 81156 32068 81180 32070
rect 81236 32068 81260 32070
rect 81020 32048 81316 32068
rect 81020 31036 81316 31056
rect 81076 31034 81100 31036
rect 81156 31034 81180 31036
rect 81236 31034 81260 31036
rect 81098 30982 81100 31034
rect 81162 30982 81174 31034
rect 81236 30982 81238 31034
rect 81076 30980 81100 30982
rect 81156 30980 81180 30982
rect 81236 30980 81260 30982
rect 81020 30960 81316 30980
rect 80058 30696 80114 30705
rect 80058 30631 80114 30640
rect 79876 30116 79928 30122
rect 79876 30058 79928 30064
rect 79704 17190 79824 17218
rect 79692 12980 79744 12986
rect 79692 12922 79744 12928
rect 79704 11898 79732 12922
rect 79692 11892 79744 11898
rect 79692 11834 79744 11840
rect 79796 11218 79824 17190
rect 79888 13938 79916 30058
rect 80072 23866 80100 30631
rect 80520 30184 80572 30190
rect 80520 30126 80572 30132
rect 80428 25832 80480 25838
rect 80428 25774 80480 25780
rect 80060 23860 80112 23866
rect 80060 23802 80112 23808
rect 80060 20936 80112 20942
rect 80060 20878 80112 20884
rect 80072 16114 80100 20878
rect 80060 16108 80112 16114
rect 80060 16050 80112 16056
rect 79876 13932 79928 13938
rect 79876 13874 79928 13880
rect 79784 11212 79836 11218
rect 79784 11154 79836 11160
rect 80060 4684 80112 4690
rect 80060 4626 80112 4632
rect 79600 3596 79652 3602
rect 79600 3538 79652 3544
rect 79508 2644 79560 2650
rect 79508 2586 79560 2592
rect 79612 1442 79640 3538
rect 79784 2916 79836 2922
rect 79784 2858 79836 2864
rect 79520 1414 79640 1442
rect 79520 800 79548 1414
rect 79796 800 79824 2858
rect 80072 2802 80100 4626
rect 80244 3664 80296 3670
rect 80244 3606 80296 3612
rect 80152 3596 80204 3602
rect 80152 3538 80204 3544
rect 79980 2774 80100 2802
rect 79980 800 80008 2774
rect 80164 800 80192 3538
rect 80256 2650 80284 3606
rect 80336 2916 80388 2922
rect 80336 2858 80388 2864
rect 80244 2644 80296 2650
rect 80244 2586 80296 2592
rect 80348 800 80376 2858
rect 80440 2106 80468 25774
rect 80532 6798 80560 30126
rect 80888 30048 80940 30054
rect 80888 29990 80940 29996
rect 80900 28422 80928 29990
rect 81020 29948 81316 29968
rect 81076 29946 81100 29948
rect 81156 29946 81180 29948
rect 81236 29946 81260 29948
rect 81098 29894 81100 29946
rect 81162 29894 81174 29946
rect 81236 29894 81238 29946
rect 81076 29892 81100 29894
rect 81156 29892 81180 29894
rect 81236 29892 81260 29894
rect 81020 29872 81316 29892
rect 81020 28860 81316 28880
rect 81076 28858 81100 28860
rect 81156 28858 81180 28860
rect 81236 28858 81260 28860
rect 81098 28806 81100 28858
rect 81162 28806 81174 28858
rect 81236 28806 81238 28858
rect 81076 28804 81100 28806
rect 81156 28804 81180 28806
rect 81236 28804 81260 28806
rect 81020 28784 81316 28804
rect 80888 28416 80940 28422
rect 80888 28358 80940 28364
rect 80900 27062 80928 28358
rect 81020 27772 81316 27792
rect 81076 27770 81100 27772
rect 81156 27770 81180 27772
rect 81236 27770 81260 27772
rect 81098 27718 81100 27770
rect 81162 27718 81174 27770
rect 81236 27718 81238 27770
rect 81076 27716 81100 27718
rect 81156 27716 81180 27718
rect 81236 27716 81260 27718
rect 81020 27696 81316 27716
rect 80888 27056 80940 27062
rect 80888 26998 80940 27004
rect 80900 26926 80928 26998
rect 80888 26920 80940 26926
rect 80888 26862 80940 26868
rect 81020 26684 81316 26704
rect 81076 26682 81100 26684
rect 81156 26682 81180 26684
rect 81236 26682 81260 26684
rect 81098 26630 81100 26682
rect 81162 26630 81174 26682
rect 81236 26630 81238 26682
rect 81076 26628 81100 26630
rect 81156 26628 81180 26630
rect 81236 26628 81260 26630
rect 81020 26608 81316 26628
rect 81020 25596 81316 25616
rect 81076 25594 81100 25596
rect 81156 25594 81180 25596
rect 81236 25594 81260 25596
rect 81098 25542 81100 25594
rect 81162 25542 81174 25594
rect 81236 25542 81238 25594
rect 81076 25540 81100 25542
rect 81156 25540 81180 25542
rect 81236 25540 81260 25542
rect 81020 25520 81316 25540
rect 81020 24508 81316 24528
rect 81076 24506 81100 24508
rect 81156 24506 81180 24508
rect 81236 24506 81260 24508
rect 81098 24454 81100 24506
rect 81162 24454 81174 24506
rect 81236 24454 81238 24506
rect 81076 24452 81100 24454
rect 81156 24452 81180 24454
rect 81236 24452 81260 24454
rect 81020 24432 81316 24452
rect 81020 23420 81316 23440
rect 81076 23418 81100 23420
rect 81156 23418 81180 23420
rect 81236 23418 81260 23420
rect 81098 23366 81100 23418
rect 81162 23366 81174 23418
rect 81236 23366 81238 23418
rect 81076 23364 81100 23366
rect 81156 23364 81180 23366
rect 81236 23364 81260 23366
rect 81020 23344 81316 23364
rect 81020 22332 81316 22352
rect 81076 22330 81100 22332
rect 81156 22330 81180 22332
rect 81236 22330 81260 22332
rect 81098 22278 81100 22330
rect 81162 22278 81174 22330
rect 81236 22278 81238 22330
rect 81076 22276 81100 22278
rect 81156 22276 81180 22278
rect 81236 22276 81260 22278
rect 81020 22256 81316 22276
rect 80704 21616 80756 21622
rect 80704 21558 80756 21564
rect 80716 21486 80744 21558
rect 80704 21480 80756 21486
rect 80704 21422 80756 21428
rect 81020 21244 81316 21264
rect 81076 21242 81100 21244
rect 81156 21242 81180 21244
rect 81236 21242 81260 21244
rect 81098 21190 81100 21242
rect 81162 21190 81174 21242
rect 81236 21190 81238 21242
rect 81076 21188 81100 21190
rect 81156 21188 81180 21190
rect 81236 21188 81260 21190
rect 81020 21168 81316 21188
rect 80978 20496 81034 20505
rect 80978 20431 80980 20440
rect 81032 20431 81034 20440
rect 80980 20402 81032 20408
rect 81020 20156 81316 20176
rect 81076 20154 81100 20156
rect 81156 20154 81180 20156
rect 81236 20154 81260 20156
rect 81098 20102 81100 20154
rect 81162 20102 81174 20154
rect 81236 20102 81238 20154
rect 81076 20100 81100 20102
rect 81156 20100 81180 20102
rect 81236 20100 81260 20102
rect 81020 20080 81316 20100
rect 81020 19068 81316 19088
rect 81076 19066 81100 19068
rect 81156 19066 81180 19068
rect 81236 19066 81260 19068
rect 81098 19014 81100 19066
rect 81162 19014 81174 19066
rect 81236 19014 81238 19066
rect 81076 19012 81100 19014
rect 81156 19012 81180 19014
rect 81236 19012 81260 19014
rect 81020 18992 81316 19012
rect 81020 17980 81316 18000
rect 81076 17978 81100 17980
rect 81156 17978 81180 17980
rect 81236 17978 81260 17980
rect 81098 17926 81100 17978
rect 81162 17926 81174 17978
rect 81236 17926 81238 17978
rect 81076 17924 81100 17926
rect 81156 17924 81180 17926
rect 81236 17924 81260 17926
rect 81020 17904 81316 17924
rect 81020 16892 81316 16912
rect 81076 16890 81100 16892
rect 81156 16890 81180 16892
rect 81236 16890 81260 16892
rect 81098 16838 81100 16890
rect 81162 16838 81174 16890
rect 81236 16838 81238 16890
rect 81076 16836 81100 16838
rect 81156 16836 81180 16838
rect 81236 16836 81260 16838
rect 81020 16816 81316 16836
rect 81020 15804 81316 15824
rect 81076 15802 81100 15804
rect 81156 15802 81180 15804
rect 81236 15802 81260 15804
rect 81098 15750 81100 15802
rect 81162 15750 81174 15802
rect 81236 15750 81238 15802
rect 81076 15748 81100 15750
rect 81156 15748 81180 15750
rect 81236 15748 81260 15750
rect 81020 15728 81316 15748
rect 81020 14716 81316 14736
rect 81076 14714 81100 14716
rect 81156 14714 81180 14716
rect 81236 14714 81260 14716
rect 81098 14662 81100 14714
rect 81162 14662 81174 14714
rect 81236 14662 81238 14714
rect 81076 14660 81100 14662
rect 81156 14660 81180 14662
rect 81236 14660 81260 14662
rect 81020 14640 81316 14660
rect 81348 13728 81400 13734
rect 81348 13670 81400 13676
rect 81020 13628 81316 13648
rect 81076 13626 81100 13628
rect 81156 13626 81180 13628
rect 81236 13626 81260 13628
rect 81098 13574 81100 13626
rect 81162 13574 81174 13626
rect 81236 13574 81238 13626
rect 81076 13572 81100 13574
rect 81156 13572 81180 13574
rect 81236 13572 81260 13574
rect 81020 13552 81316 13572
rect 81360 13258 81388 13670
rect 81348 13252 81400 13258
rect 81348 13194 81400 13200
rect 81020 12540 81316 12560
rect 81076 12538 81100 12540
rect 81156 12538 81180 12540
rect 81236 12538 81260 12540
rect 81098 12486 81100 12538
rect 81162 12486 81174 12538
rect 81236 12486 81238 12538
rect 81076 12484 81100 12486
rect 81156 12484 81180 12486
rect 81236 12484 81260 12486
rect 81020 12464 81316 12484
rect 81020 11452 81316 11472
rect 81076 11450 81100 11452
rect 81156 11450 81180 11452
rect 81236 11450 81260 11452
rect 81098 11398 81100 11450
rect 81162 11398 81174 11450
rect 81236 11398 81238 11450
rect 81076 11396 81100 11398
rect 81156 11396 81180 11398
rect 81236 11396 81260 11398
rect 81020 11376 81316 11396
rect 81020 10364 81316 10384
rect 81076 10362 81100 10364
rect 81156 10362 81180 10364
rect 81236 10362 81260 10364
rect 81098 10310 81100 10362
rect 81162 10310 81174 10362
rect 81236 10310 81238 10362
rect 81076 10308 81100 10310
rect 81156 10308 81180 10310
rect 81236 10308 81260 10310
rect 81020 10288 81316 10308
rect 81020 9276 81316 9296
rect 81076 9274 81100 9276
rect 81156 9274 81180 9276
rect 81236 9274 81260 9276
rect 81098 9222 81100 9274
rect 81162 9222 81174 9274
rect 81236 9222 81238 9274
rect 81076 9220 81100 9222
rect 81156 9220 81180 9222
rect 81236 9220 81260 9222
rect 81020 9200 81316 9220
rect 81020 8188 81316 8208
rect 81076 8186 81100 8188
rect 81156 8186 81180 8188
rect 81236 8186 81260 8188
rect 81098 8134 81100 8186
rect 81162 8134 81174 8186
rect 81236 8134 81238 8186
rect 81076 8132 81100 8134
rect 81156 8132 81180 8134
rect 81236 8132 81260 8134
rect 81020 8112 81316 8132
rect 81020 7100 81316 7120
rect 81076 7098 81100 7100
rect 81156 7098 81180 7100
rect 81236 7098 81260 7100
rect 81098 7046 81100 7098
rect 81162 7046 81174 7098
rect 81236 7046 81238 7098
rect 81076 7044 81100 7046
rect 81156 7044 81180 7046
rect 81236 7044 81260 7046
rect 81020 7024 81316 7044
rect 80520 6792 80572 6798
rect 80520 6734 80572 6740
rect 81348 6656 81400 6662
rect 81348 6598 81400 6604
rect 81360 6322 81388 6598
rect 81348 6316 81400 6322
rect 81348 6258 81400 6264
rect 81452 6186 81480 37266
rect 81624 36236 81676 36242
rect 81624 36178 81676 36184
rect 81636 30122 81664 36178
rect 82004 35630 82032 38218
rect 82832 37466 82860 39200
rect 83660 37466 83688 39200
rect 82820 37460 82872 37466
rect 82820 37402 82872 37408
rect 83648 37460 83700 37466
rect 83648 37402 83700 37408
rect 82912 37324 82964 37330
rect 82912 37266 82964 37272
rect 84200 37324 84252 37330
rect 84200 37266 84252 37272
rect 82360 35692 82412 35698
rect 82360 35634 82412 35640
rect 81900 35624 81952 35630
rect 81900 35566 81952 35572
rect 81992 35624 82044 35630
rect 81992 35566 82044 35572
rect 82176 35624 82228 35630
rect 82176 35566 82228 35572
rect 81912 31754 81940 35566
rect 81820 31726 81940 31754
rect 81624 30116 81676 30122
rect 81624 30058 81676 30064
rect 81820 26246 81848 31726
rect 81900 30116 81952 30122
rect 81900 30058 81952 30064
rect 81808 26240 81860 26246
rect 81808 26182 81860 26188
rect 81820 25362 81848 26182
rect 81808 25356 81860 25362
rect 81808 25298 81860 25304
rect 81912 23186 81940 30058
rect 82188 25770 82216 35566
rect 82176 25764 82228 25770
rect 82176 25706 82228 25712
rect 82372 25498 82400 35634
rect 82924 29578 82952 37266
rect 83738 34640 83794 34649
rect 83464 34604 83516 34610
rect 83738 34575 83794 34584
rect 83464 34546 83516 34552
rect 83280 34536 83332 34542
rect 83280 34478 83332 34484
rect 82912 29572 82964 29578
rect 82912 29514 82964 29520
rect 83292 27402 83320 34478
rect 83280 27396 83332 27402
rect 83280 27338 83332 27344
rect 82728 25764 82780 25770
rect 82728 25706 82780 25712
rect 82360 25492 82412 25498
rect 82360 25434 82412 25440
rect 82740 25430 82768 25706
rect 82728 25424 82780 25430
rect 82728 25366 82780 25372
rect 83188 24268 83240 24274
rect 83188 24210 83240 24216
rect 81900 23180 81952 23186
rect 81900 23122 81952 23128
rect 82452 21480 82504 21486
rect 82452 21422 82504 21428
rect 81532 21140 81584 21146
rect 81532 21082 81584 21088
rect 81544 20398 81572 21082
rect 81624 20596 81676 20602
rect 81624 20538 81676 20544
rect 81532 20392 81584 20398
rect 81636 20380 81664 20538
rect 81716 20528 81768 20534
rect 81900 20528 81952 20534
rect 81768 20476 81900 20482
rect 81716 20470 81952 20476
rect 82266 20496 82322 20505
rect 81728 20454 81940 20470
rect 82266 20431 82268 20440
rect 82320 20431 82322 20440
rect 82268 20402 82320 20408
rect 81716 20392 81768 20398
rect 81636 20352 81716 20380
rect 81532 20334 81584 20340
rect 81716 20334 81768 20340
rect 81900 20392 81952 20398
rect 81900 20334 81952 20340
rect 82084 20392 82136 20398
rect 82176 20392 82228 20398
rect 82084 20334 82136 20340
rect 82174 20360 82176 20369
rect 82360 20392 82412 20398
rect 82228 20360 82230 20369
rect 81808 20256 81860 20262
rect 81912 20210 81940 20334
rect 81860 20204 81940 20210
rect 81808 20198 81940 20204
rect 81820 20182 81940 20198
rect 81912 14618 81940 20182
rect 82096 18902 82124 20334
rect 82360 20334 82412 20340
rect 82174 20295 82230 20304
rect 82084 18896 82136 18902
rect 82084 18838 82136 18844
rect 81900 14612 81952 14618
rect 81900 14554 81952 14560
rect 81716 14340 81768 14346
rect 81716 14282 81768 14288
rect 81728 10130 81756 14282
rect 81900 14272 81952 14278
rect 81900 14214 81952 14220
rect 81912 12782 81940 14214
rect 82084 13184 82136 13190
rect 82084 13126 82136 13132
rect 81900 12776 81952 12782
rect 81900 12718 81952 12724
rect 81716 10124 81768 10130
rect 81716 10066 81768 10072
rect 81728 7954 81756 10066
rect 81716 7948 81768 7954
rect 81716 7890 81768 7896
rect 81900 7948 81952 7954
rect 81900 7890 81952 7896
rect 81912 6254 81940 7890
rect 81900 6248 81952 6254
rect 81900 6190 81952 6196
rect 81440 6180 81492 6186
rect 81440 6122 81492 6128
rect 81020 6012 81316 6032
rect 81076 6010 81100 6012
rect 81156 6010 81180 6012
rect 81236 6010 81260 6012
rect 81098 5958 81100 6010
rect 81162 5958 81174 6010
rect 81236 5958 81238 6010
rect 81076 5956 81100 5958
rect 81156 5956 81180 5958
rect 81236 5956 81260 5958
rect 81020 5936 81316 5956
rect 81020 4924 81316 4944
rect 81076 4922 81100 4924
rect 81156 4922 81180 4924
rect 81236 4922 81260 4924
rect 81098 4870 81100 4922
rect 81162 4870 81174 4922
rect 81236 4870 81238 4922
rect 81076 4868 81100 4870
rect 81156 4868 81180 4870
rect 81236 4868 81260 4870
rect 81020 4848 81316 4868
rect 80520 4616 80572 4622
rect 80520 4558 80572 4564
rect 80428 2100 80480 2106
rect 80428 2042 80480 2048
rect 80532 800 80560 4558
rect 80796 4072 80848 4078
rect 80796 4014 80848 4020
rect 81348 4072 81400 4078
rect 81348 4014 81400 4020
rect 81992 4072 82044 4078
rect 81992 4014 82044 4020
rect 80808 800 80836 4014
rect 80888 4004 80940 4010
rect 80888 3946 80940 3952
rect 80900 3194 80928 3946
rect 81020 3836 81316 3856
rect 81076 3834 81100 3836
rect 81156 3834 81180 3836
rect 81236 3834 81260 3836
rect 81098 3782 81100 3834
rect 81162 3782 81174 3834
rect 81236 3782 81238 3834
rect 81076 3780 81100 3782
rect 81156 3780 81180 3782
rect 81236 3780 81260 3782
rect 81020 3760 81316 3780
rect 80888 3188 80940 3194
rect 80888 3130 80940 3136
rect 80888 2984 80940 2990
rect 80888 2926 80940 2932
rect 80900 898 80928 2926
rect 81020 2748 81316 2768
rect 81076 2746 81100 2748
rect 81156 2746 81180 2748
rect 81236 2746 81260 2748
rect 81098 2694 81100 2746
rect 81162 2694 81174 2746
rect 81236 2694 81238 2746
rect 81076 2692 81100 2694
rect 81156 2692 81180 2694
rect 81236 2692 81260 2694
rect 81020 2672 81316 2692
rect 81164 2100 81216 2106
rect 81164 2042 81216 2048
rect 80900 870 81020 898
rect 80992 800 81020 870
rect 81176 800 81204 2042
rect 81360 800 81388 4014
rect 81532 3460 81584 3466
rect 81532 3402 81584 3408
rect 81544 800 81572 3402
rect 81808 3188 81860 3194
rect 81808 3130 81860 3136
rect 81820 800 81848 3130
rect 82004 800 82032 4014
rect 78036 672 78088 678
rect 78036 614 78088 620
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78770 0 78826 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81346 0 81402 800
rect 81530 0 81586 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82096 649 82124 13126
rect 82372 9586 82400 20334
rect 82360 9580 82412 9586
rect 82360 9522 82412 9528
rect 82464 7562 82492 21422
rect 82728 18692 82780 18698
rect 82728 18634 82780 18640
rect 82740 18222 82768 18634
rect 82728 18216 82780 18222
rect 82728 18158 82780 18164
rect 82740 13870 82768 18158
rect 83096 17604 83148 17610
rect 83096 17546 83148 17552
rect 82728 13864 82780 13870
rect 82728 13806 82780 13812
rect 83108 13394 83136 17546
rect 83096 13388 83148 13394
rect 83096 13330 83148 13336
rect 82636 11212 82688 11218
rect 82636 11154 82688 11160
rect 82648 10606 82676 11154
rect 83096 11008 83148 11014
rect 83096 10950 83148 10956
rect 82636 10600 82688 10606
rect 82636 10542 82688 10548
rect 82280 7534 82492 7562
rect 82176 5364 82228 5370
rect 82176 5306 82228 5312
rect 82188 5234 82216 5306
rect 82176 5228 82228 5234
rect 82176 5170 82228 5176
rect 82188 5098 82216 5170
rect 82176 5092 82228 5098
rect 82176 5034 82228 5040
rect 82176 2848 82228 2854
rect 82176 2790 82228 2796
rect 82188 800 82216 2790
rect 82280 1970 82308 7534
rect 82452 7472 82504 7478
rect 82452 7414 82504 7420
rect 82360 3732 82412 3738
rect 82360 3674 82412 3680
rect 82268 1964 82320 1970
rect 82268 1906 82320 1912
rect 82372 800 82400 3674
rect 82464 2582 82492 7414
rect 82648 5234 82676 10542
rect 82636 5228 82688 5234
rect 82636 5170 82688 5176
rect 82912 4684 82964 4690
rect 82912 4626 82964 4632
rect 82728 4072 82780 4078
rect 82728 4014 82780 4020
rect 82636 2984 82688 2990
rect 82636 2926 82688 2932
rect 82648 2774 82676 2926
rect 82556 2746 82676 2774
rect 82452 2576 82504 2582
rect 82452 2518 82504 2524
rect 82556 800 82584 2746
rect 82740 2106 82768 4014
rect 82924 3194 82952 4626
rect 83004 3596 83056 3602
rect 83004 3538 83056 3544
rect 82912 3188 82964 3194
rect 82912 3130 82964 3136
rect 82820 2372 82872 2378
rect 82820 2314 82872 2320
rect 82728 2100 82780 2106
rect 82728 2042 82780 2048
rect 82832 800 82860 2314
rect 83016 800 83044 3538
rect 83108 2582 83136 10950
rect 83200 6730 83228 24210
rect 83292 17134 83320 27338
rect 83280 17128 83332 17134
rect 83280 17070 83332 17076
rect 83292 7954 83320 17070
rect 83372 13320 83424 13326
rect 83372 13262 83424 13268
rect 83280 7948 83332 7954
rect 83280 7890 83332 7896
rect 83384 7750 83412 13262
rect 83372 7744 83424 7750
rect 83372 7686 83424 7692
rect 83188 6724 83240 6730
rect 83188 6666 83240 6672
rect 83476 3194 83504 34546
rect 83556 27464 83608 27470
rect 83556 27406 83608 27412
rect 83568 26314 83596 27406
rect 83556 26308 83608 26314
rect 83556 26250 83608 26256
rect 83648 26308 83700 26314
rect 83648 26250 83700 26256
rect 83556 24268 83608 24274
rect 83556 24210 83608 24216
rect 83568 23730 83596 24210
rect 83556 23724 83608 23730
rect 83556 23666 83608 23672
rect 83660 17610 83688 26250
rect 83648 17604 83700 17610
rect 83648 17546 83700 17552
rect 83752 15434 83780 34575
rect 83832 33312 83884 33318
rect 83832 33254 83884 33260
rect 83844 23798 83872 33254
rect 84212 31754 84240 37266
rect 84580 36718 84608 39200
rect 85212 37664 85264 37670
rect 85212 37606 85264 37612
rect 85224 37398 85252 37606
rect 85408 37398 85436 39200
rect 86224 38208 86276 38214
rect 86224 38150 86276 38156
rect 86040 37936 86092 37942
rect 86040 37878 86092 37884
rect 85212 37392 85264 37398
rect 85212 37334 85264 37340
rect 85396 37392 85448 37398
rect 85396 37334 85448 37340
rect 85488 37392 85540 37398
rect 85488 37334 85540 37340
rect 84568 36712 84620 36718
rect 84568 36654 84620 36660
rect 84658 36136 84714 36145
rect 84658 36071 84714 36080
rect 84200 31748 84252 31754
rect 84200 31690 84252 31696
rect 84212 31482 84240 31690
rect 84200 31476 84252 31482
rect 84200 31418 84252 31424
rect 84476 30048 84528 30054
rect 84476 29990 84528 29996
rect 84488 29646 84516 29990
rect 84476 29640 84528 29646
rect 84476 29582 84528 29588
rect 84108 29572 84160 29578
rect 84108 29514 84160 29520
rect 84120 29238 84148 29514
rect 83924 29232 83976 29238
rect 83924 29174 83976 29180
rect 84108 29232 84160 29238
rect 84108 29174 84160 29180
rect 83832 23792 83884 23798
rect 83832 23734 83884 23740
rect 83936 15570 83964 29174
rect 84200 28076 84252 28082
rect 84200 28018 84252 28024
rect 84016 24200 84068 24206
rect 84016 24142 84068 24148
rect 84028 23866 84056 24142
rect 84016 23860 84068 23866
rect 84016 23802 84068 23808
rect 84212 21146 84240 28018
rect 84200 21140 84252 21146
rect 84200 21082 84252 21088
rect 83924 15564 83976 15570
rect 83924 15506 83976 15512
rect 83740 15428 83792 15434
rect 83740 15370 83792 15376
rect 83936 7206 83964 15506
rect 84200 7336 84252 7342
rect 84200 7278 84252 7284
rect 83924 7200 83976 7206
rect 83924 7142 83976 7148
rect 84212 6322 84240 7278
rect 84200 6316 84252 6322
rect 84200 6258 84252 6264
rect 83740 5704 83792 5710
rect 83740 5646 83792 5652
rect 83556 4684 83608 4690
rect 83556 4626 83608 4632
rect 83568 3738 83596 4626
rect 83648 4072 83700 4078
rect 83648 4014 83700 4020
rect 83556 3732 83608 3738
rect 83556 3674 83608 3680
rect 83464 3188 83516 3194
rect 83464 3130 83516 3136
rect 83280 2984 83332 2990
rect 83280 2926 83332 2932
rect 83292 2774 83320 2926
rect 83200 2746 83320 2774
rect 83096 2576 83148 2582
rect 83096 2518 83148 2524
rect 83200 800 83228 2746
rect 83372 2304 83424 2310
rect 83372 2246 83424 2252
rect 83384 800 83412 2246
rect 83660 800 83688 4014
rect 83752 3466 83780 5646
rect 84292 4752 84344 4758
rect 84292 4694 84344 4700
rect 84200 4072 84252 4078
rect 84200 4014 84252 4020
rect 83832 3596 83884 3602
rect 83832 3538 83884 3544
rect 83740 3460 83792 3466
rect 83740 3402 83792 3408
rect 83844 800 83872 3538
rect 84016 2304 84068 2310
rect 84016 2246 84068 2252
rect 84028 800 84056 2246
rect 84212 800 84240 4014
rect 84304 2514 84332 4694
rect 84384 3596 84436 3602
rect 84384 3538 84436 3544
rect 84292 2508 84344 2514
rect 84292 2450 84344 2456
rect 84396 800 84424 3538
rect 84672 2514 84700 36071
rect 85500 34202 85528 37334
rect 84844 34196 84896 34202
rect 84844 34138 84896 34144
rect 85488 34196 85540 34202
rect 85488 34138 85540 34144
rect 84856 33454 84884 34138
rect 84844 33448 84896 33454
rect 84844 33390 84896 33396
rect 84752 32360 84804 32366
rect 84752 32302 84804 32308
rect 84764 31958 84792 32302
rect 84752 31952 84804 31958
rect 84752 31894 84804 31900
rect 84856 31754 84884 33390
rect 85764 32564 85816 32570
rect 85764 32506 85816 32512
rect 84856 31726 84976 31754
rect 84844 27328 84896 27334
rect 84844 27270 84896 27276
rect 84856 27130 84884 27270
rect 84844 27124 84896 27130
rect 84844 27066 84896 27072
rect 84948 23662 84976 31726
rect 85580 27872 85632 27878
rect 85580 27814 85632 27820
rect 84936 23656 84988 23662
rect 84936 23598 84988 23604
rect 84948 22094 84976 23598
rect 84856 22066 84976 22094
rect 85488 22092 85540 22098
rect 84752 15904 84804 15910
rect 84752 15846 84804 15852
rect 84764 15706 84792 15846
rect 84752 15700 84804 15706
rect 84752 15642 84804 15648
rect 84856 6254 84884 22066
rect 85488 22034 85540 22040
rect 85304 22024 85356 22030
rect 85302 21992 85304 22001
rect 85356 21992 85358 22001
rect 85302 21927 85358 21936
rect 85120 21888 85172 21894
rect 85120 21830 85172 21836
rect 84844 6248 84896 6254
rect 84844 6190 84896 6196
rect 84844 4072 84896 4078
rect 84844 4014 84896 4020
rect 84660 2508 84712 2514
rect 84660 2450 84712 2456
rect 84752 2440 84804 2446
rect 84752 2382 84804 2388
rect 84764 1170 84792 2382
rect 84672 1142 84792 1170
rect 84672 800 84700 1142
rect 84856 800 84884 4014
rect 85028 3596 85080 3602
rect 85028 3538 85080 3544
rect 85040 800 85068 3538
rect 85132 1057 85160 21830
rect 85500 21690 85528 22034
rect 85488 21684 85540 21690
rect 85488 21626 85540 21632
rect 85592 21078 85620 27814
rect 85580 21072 85632 21078
rect 85580 21014 85632 21020
rect 85488 16448 85540 16454
rect 85488 16390 85540 16396
rect 85500 16114 85528 16390
rect 85488 16108 85540 16114
rect 85488 16050 85540 16056
rect 85396 12640 85448 12646
rect 85396 12582 85448 12588
rect 85408 12374 85436 12582
rect 85396 12368 85448 12374
rect 85396 12310 85448 12316
rect 85500 11830 85528 16050
rect 85672 13456 85724 13462
rect 85672 13398 85724 13404
rect 85580 12912 85632 12918
rect 85578 12880 85580 12889
rect 85632 12880 85634 12889
rect 85578 12815 85634 12824
rect 85580 12776 85632 12782
rect 85580 12718 85632 12724
rect 85488 11824 85540 11830
rect 85488 11766 85540 11772
rect 85500 4758 85528 11766
rect 85592 7313 85620 12718
rect 85684 12646 85712 13398
rect 85672 12640 85724 12646
rect 85672 12582 85724 12588
rect 85672 12368 85724 12374
rect 85672 12310 85724 12316
rect 85578 7304 85634 7313
rect 85578 7239 85634 7248
rect 85488 4752 85540 4758
rect 85488 4694 85540 4700
rect 85396 4684 85448 4690
rect 85396 4626 85448 4632
rect 85304 2508 85356 2514
rect 85304 2450 85356 2456
rect 85316 1170 85344 2450
rect 85224 1142 85344 1170
rect 85118 1048 85174 1057
rect 85118 983 85174 992
rect 85224 800 85252 1142
rect 85408 800 85436 4626
rect 85684 4010 85712 12310
rect 85672 4004 85724 4010
rect 85672 3946 85724 3952
rect 85672 2984 85724 2990
rect 85672 2926 85724 2932
rect 85684 800 85712 2926
rect 85776 2650 85804 32506
rect 86052 30938 86080 37878
rect 86236 37346 86264 38150
rect 86328 37466 86356 39200
rect 86960 37732 87012 37738
rect 86960 37674 87012 37680
rect 86316 37460 86368 37466
rect 86316 37402 86368 37408
rect 86236 37318 86356 37346
rect 86328 35154 86356 37318
rect 86972 36922 87000 37674
rect 87052 37664 87104 37670
rect 87052 37606 87104 37612
rect 86960 36916 87012 36922
rect 86960 36858 87012 36864
rect 86316 35148 86368 35154
rect 86316 35090 86368 35096
rect 86408 35080 86460 35086
rect 86408 35022 86460 35028
rect 86040 30932 86092 30938
rect 86040 30874 86092 30880
rect 86316 30864 86368 30870
rect 86420 30818 86448 35022
rect 86684 35012 86736 35018
rect 86684 34954 86736 34960
rect 86592 31680 86644 31686
rect 86592 31622 86644 31628
rect 86368 30812 86448 30818
rect 86316 30806 86448 30812
rect 86328 30790 86448 30806
rect 86604 30802 86632 31622
rect 86696 31142 86724 34954
rect 86868 34944 86920 34950
rect 86868 34886 86920 34892
rect 86880 34678 86908 34886
rect 86868 34672 86920 34678
rect 86868 34614 86920 34620
rect 87064 34610 87092 37606
rect 87156 36718 87184 39200
rect 87880 37664 87932 37670
rect 87880 37606 87932 37612
rect 87892 37398 87920 37606
rect 88076 37398 88104 39200
rect 88996 38418 89024 39200
rect 88984 38412 89036 38418
rect 88984 38354 89036 38360
rect 89456 37398 89484 39238
rect 89810 39200 89866 40000
rect 90730 39200 90786 40000
rect 91558 39200 91614 40000
rect 92478 39200 92534 40000
rect 93306 39200 93362 40000
rect 94226 39200 94282 40000
rect 95054 39200 95110 40000
rect 95974 39200 96030 40000
rect 96802 39200 96858 40000
rect 97722 39200 97778 40000
rect 98550 39200 98606 40000
rect 99470 39200 99526 40000
rect 89628 38412 89680 38418
rect 89628 38354 89680 38360
rect 89640 37482 89668 38354
rect 89640 37466 89760 37482
rect 89640 37460 89772 37466
rect 89640 37454 89720 37460
rect 89720 37402 89772 37408
rect 87880 37392 87932 37398
rect 87880 37334 87932 37340
rect 88064 37392 88116 37398
rect 88064 37334 88116 37340
rect 89444 37392 89496 37398
rect 89444 37334 89496 37340
rect 88984 36848 89036 36854
rect 88984 36790 89036 36796
rect 87144 36712 87196 36718
rect 87144 36654 87196 36660
rect 88340 35760 88392 35766
rect 88340 35702 88392 35708
rect 87052 34604 87104 34610
rect 87052 34546 87104 34552
rect 87328 32224 87380 32230
rect 87328 32166 87380 32172
rect 87788 32224 87840 32230
rect 87788 32166 87840 32172
rect 87236 31272 87288 31278
rect 87236 31214 87288 31220
rect 87248 31142 87276 31214
rect 86684 31136 86736 31142
rect 86684 31078 86736 31084
rect 87236 31136 87288 31142
rect 87236 31078 87288 31084
rect 86224 30184 86276 30190
rect 86224 30126 86276 30132
rect 86236 29238 86264 30126
rect 86224 29232 86276 29238
rect 86224 29174 86276 29180
rect 86236 26994 86264 29174
rect 86224 26988 86276 26994
rect 86224 26930 86276 26936
rect 86420 26874 86448 30790
rect 86592 30796 86644 30802
rect 86592 30738 86644 30744
rect 86776 30592 86828 30598
rect 86776 30534 86828 30540
rect 86592 29096 86644 29102
rect 86592 29038 86644 29044
rect 86500 26988 86552 26994
rect 86500 26930 86552 26936
rect 86236 26846 86448 26874
rect 86132 26376 86184 26382
rect 86130 26344 86132 26353
rect 86184 26344 86186 26353
rect 86130 26279 86186 26288
rect 86236 14074 86264 26846
rect 86316 26444 86368 26450
rect 86408 26444 86460 26450
rect 86368 26404 86408 26432
rect 86316 26386 86368 26392
rect 86408 26386 86460 26392
rect 86316 26308 86368 26314
rect 86316 26250 86368 26256
rect 86328 21622 86356 26250
rect 86316 21616 86368 21622
rect 86316 21558 86368 21564
rect 86224 14068 86276 14074
rect 86224 14010 86276 14016
rect 86038 12880 86094 12889
rect 86038 12815 86094 12824
rect 86052 12782 86080 12815
rect 85856 12776 85908 12782
rect 85856 12718 85908 12724
rect 86040 12776 86092 12782
rect 86040 12718 86092 12724
rect 85868 12646 85896 12718
rect 85856 12640 85908 12646
rect 85856 12582 85908 12588
rect 86512 11082 86540 26930
rect 86604 26330 86632 29038
rect 86684 26920 86736 26926
rect 86684 26862 86736 26868
rect 86696 26450 86724 26862
rect 86684 26444 86736 26450
rect 86684 26386 86736 26392
rect 86604 26302 86724 26330
rect 86592 25900 86644 25906
rect 86592 25842 86644 25848
rect 86500 11076 86552 11082
rect 86500 11018 86552 11024
rect 85948 10668 86000 10674
rect 85948 10610 86000 10616
rect 85960 9382 85988 10610
rect 85948 9376 86000 9382
rect 85948 9318 86000 9324
rect 85960 6254 85988 9318
rect 86604 6322 86632 25842
rect 86696 7274 86724 26302
rect 86788 10198 86816 30534
rect 86960 29164 87012 29170
rect 86960 29106 87012 29112
rect 86868 27464 86920 27470
rect 86868 27406 86920 27412
rect 86880 26926 86908 27406
rect 86868 26920 86920 26926
rect 86868 26862 86920 26868
rect 86868 26444 86920 26450
rect 86868 26386 86920 26392
rect 86880 24410 86908 26386
rect 86868 24404 86920 24410
rect 86868 24346 86920 24352
rect 86972 19922 87000 29106
rect 87052 27396 87104 27402
rect 87052 27338 87104 27344
rect 87064 26450 87092 27338
rect 87052 26444 87104 26450
rect 87052 26386 87104 26392
rect 86960 19916 87012 19922
rect 86960 19858 87012 19864
rect 86776 10192 86828 10198
rect 86776 10134 86828 10140
rect 86960 9512 87012 9518
rect 86960 9454 87012 9460
rect 86972 7290 87000 9454
rect 87052 9104 87104 9110
rect 87052 9046 87104 9052
rect 87064 7410 87092 9046
rect 87248 7478 87276 31078
rect 87236 7472 87288 7478
rect 87236 7414 87288 7420
rect 87052 7404 87104 7410
rect 87052 7346 87104 7352
rect 86684 7268 86736 7274
rect 86972 7262 87092 7290
rect 86684 7210 86736 7216
rect 86592 6316 86644 6322
rect 86592 6258 86644 6264
rect 85948 6248 86000 6254
rect 85948 6190 86000 6196
rect 86040 4684 86092 4690
rect 86040 4626 86092 4632
rect 86960 4684 87012 4690
rect 86960 4626 87012 4632
rect 85948 3188 86000 3194
rect 85948 3130 86000 3136
rect 85960 2922 85988 3130
rect 85856 2916 85908 2922
rect 85856 2858 85908 2864
rect 85948 2916 86000 2922
rect 85948 2858 86000 2864
rect 85764 2644 85816 2650
rect 85764 2586 85816 2592
rect 85868 800 85896 2858
rect 86052 800 86080 4626
rect 86972 3754 87000 4626
rect 86696 3726 87000 3754
rect 86224 3596 86276 3602
rect 86224 3538 86276 3544
rect 86236 800 86264 3538
rect 86408 2644 86460 2650
rect 86408 2586 86460 2592
rect 86420 800 86448 2586
rect 86696 800 86724 3726
rect 87064 3652 87092 7262
rect 87340 5166 87368 32166
rect 87800 31754 87828 32166
rect 87708 31726 87828 31754
rect 87708 28014 87736 31726
rect 88352 29782 88380 35702
rect 88892 34604 88944 34610
rect 88892 34546 88944 34552
rect 88800 34468 88852 34474
rect 88800 34410 88852 34416
rect 88616 30592 88668 30598
rect 88616 30534 88668 30540
rect 88340 29776 88392 29782
rect 88340 29718 88392 29724
rect 88628 28218 88656 30534
rect 88708 29572 88760 29578
rect 88708 29514 88760 29520
rect 88720 29170 88748 29514
rect 88708 29164 88760 29170
rect 88708 29106 88760 29112
rect 88616 28212 88668 28218
rect 88616 28154 88668 28160
rect 87604 28008 87656 28014
rect 87604 27950 87656 27956
rect 87696 28008 87748 28014
rect 87696 27950 87748 27956
rect 87512 27056 87564 27062
rect 87512 26998 87564 27004
rect 87420 26988 87472 26994
rect 87420 26930 87472 26936
rect 87432 25906 87460 26930
rect 87524 26790 87552 26998
rect 87512 26784 87564 26790
rect 87512 26726 87564 26732
rect 87524 26586 87552 26726
rect 87512 26580 87564 26586
rect 87512 26522 87564 26528
rect 87420 25900 87472 25906
rect 87420 25842 87472 25848
rect 87512 17128 87564 17134
rect 87512 17070 87564 17076
rect 87524 8090 87552 17070
rect 87512 8084 87564 8090
rect 87512 8026 87564 8032
rect 87616 6662 87644 27950
rect 87708 19786 87736 27950
rect 87788 26784 87840 26790
rect 87788 26726 87840 26732
rect 87800 26518 87828 26726
rect 87788 26512 87840 26518
rect 87788 26454 87840 26460
rect 87972 26376 88024 26382
rect 88248 26376 88300 26382
rect 87972 26318 88024 26324
rect 88246 26344 88248 26353
rect 88300 26344 88302 26353
rect 87984 24818 88012 26318
rect 88246 26279 88302 26288
rect 87972 24812 88024 24818
rect 87972 24754 88024 24760
rect 88248 23316 88300 23322
rect 88248 23258 88300 23264
rect 88260 21962 88288 23258
rect 88812 22094 88840 34410
rect 88904 31754 88932 34546
rect 88996 32026 89024 36790
rect 89824 36718 89852 39200
rect 90456 38752 90508 38758
rect 90456 38694 90508 38700
rect 89812 36712 89864 36718
rect 89812 36654 89864 36660
rect 90362 33552 90418 33561
rect 90362 33487 90418 33496
rect 89902 33416 89958 33425
rect 89902 33351 89958 33360
rect 89168 32292 89220 32298
rect 89168 32234 89220 32240
rect 88984 32020 89036 32026
rect 88984 31962 89036 31968
rect 89180 31890 89208 32234
rect 89536 32020 89588 32026
rect 89536 31962 89588 31968
rect 89548 31890 89576 31962
rect 89168 31884 89220 31890
rect 89168 31826 89220 31832
rect 89536 31884 89588 31890
rect 89536 31826 89588 31832
rect 89812 31816 89864 31822
rect 89812 31758 89864 31764
rect 88904 31726 89024 31754
rect 88812 22066 88932 22094
rect 88248 21956 88300 21962
rect 88248 21898 88300 21904
rect 87696 19780 87748 19786
rect 87696 19722 87748 19728
rect 88524 13728 88576 13734
rect 88524 13670 88576 13676
rect 87788 10736 87840 10742
rect 87788 10678 87840 10684
rect 87604 6656 87656 6662
rect 87604 6598 87656 6604
rect 87328 5160 87380 5166
rect 87328 5102 87380 5108
rect 87604 5160 87656 5166
rect 87604 5102 87656 5108
rect 87236 5024 87288 5030
rect 87236 4966 87288 4972
rect 87144 4140 87196 4146
rect 87144 4082 87196 4088
rect 86972 3624 87092 3652
rect 86868 3596 86920 3602
rect 86868 3538 86920 3544
rect 86880 800 86908 3538
rect 86972 2582 87000 3624
rect 87052 2848 87104 2854
rect 87052 2790 87104 2796
rect 86960 2576 87012 2582
rect 86960 2518 87012 2524
rect 87064 800 87092 2790
rect 82082 640 82138 649
rect 82082 575 82138 584
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83002 0 83058 800
rect 83186 0 83242 800
rect 83370 0 83426 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85026 0 85082 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87156 134 87184 4082
rect 87248 800 87276 4966
rect 87616 4758 87644 5102
rect 87604 4752 87656 4758
rect 87604 4694 87656 4700
rect 87616 4078 87644 4694
rect 87604 4072 87656 4078
rect 87604 4014 87656 4020
rect 87512 3596 87564 3602
rect 87512 3538 87564 3544
rect 87524 800 87552 3538
rect 87616 2990 87644 4014
rect 87604 2984 87656 2990
rect 87604 2926 87656 2932
rect 87800 2582 87828 10678
rect 88536 9110 88564 13670
rect 88524 9104 88576 9110
rect 88524 9046 88576 9052
rect 88432 8968 88484 8974
rect 88432 8910 88484 8916
rect 88340 4616 88392 4622
rect 88340 4558 88392 4564
rect 87880 3732 87932 3738
rect 87880 3674 87932 3680
rect 87788 2576 87840 2582
rect 87788 2518 87840 2524
rect 87696 2372 87748 2378
rect 87696 2314 87748 2320
rect 87708 800 87736 2314
rect 87892 800 87920 3674
rect 88064 3528 88116 3534
rect 88064 3470 88116 3476
rect 87972 2984 88024 2990
rect 87972 2926 88024 2932
rect 87984 1329 88012 2926
rect 87970 1320 88026 1329
rect 87970 1255 88026 1264
rect 88076 800 88104 3470
rect 88352 3194 88380 4558
rect 88340 3188 88392 3194
rect 88340 3130 88392 3136
rect 88248 2440 88300 2446
rect 88248 2382 88300 2388
rect 88260 800 88288 2382
rect 88340 2304 88392 2310
rect 88340 2246 88392 2252
rect 88352 882 88380 2246
rect 88444 1193 88472 8910
rect 88524 5160 88576 5166
rect 88524 5102 88576 5108
rect 88430 1184 88486 1193
rect 88430 1119 88486 1128
rect 88340 876 88392 882
rect 88340 818 88392 824
rect 88536 800 88564 5102
rect 88800 4684 88852 4690
rect 88800 4626 88852 4632
rect 88812 3738 88840 4626
rect 88800 3732 88852 3738
rect 88800 3674 88852 3680
rect 88708 3664 88760 3670
rect 88708 3606 88760 3612
rect 88616 2508 88668 2514
rect 88616 2450 88668 2456
rect 88628 2310 88656 2450
rect 88616 2304 88668 2310
rect 88616 2246 88668 2252
rect 88720 800 88748 3606
rect 88800 2848 88852 2854
rect 88800 2790 88852 2796
rect 88812 2514 88840 2790
rect 88904 2650 88932 22066
rect 88996 9042 89024 31726
rect 89628 30184 89680 30190
rect 89628 30126 89680 30132
rect 89640 29510 89668 30126
rect 89628 29504 89680 29510
rect 89628 29446 89680 29452
rect 89536 25356 89588 25362
rect 89536 25298 89588 25304
rect 89352 23180 89404 23186
rect 89352 23122 89404 23128
rect 89260 15496 89312 15502
rect 89260 15438 89312 15444
rect 89272 11257 89300 15438
rect 89258 11248 89314 11257
rect 89258 11183 89314 11192
rect 89364 9042 89392 23122
rect 89548 20398 89576 25298
rect 89536 20392 89588 20398
rect 89536 20334 89588 20340
rect 89548 18290 89576 20334
rect 89536 18284 89588 18290
rect 89536 18226 89588 18232
rect 89824 16574 89852 31758
rect 89732 16546 89852 16574
rect 89916 16574 89944 33351
rect 90088 32768 90140 32774
rect 90088 32710 90140 32716
rect 90100 23254 90128 32710
rect 90376 32026 90404 33487
rect 90364 32020 90416 32026
rect 90364 31962 90416 31968
rect 90468 26586 90496 38694
rect 90548 37664 90600 37670
rect 90548 37606 90600 37612
rect 90560 37398 90588 37606
rect 90744 37398 90772 39200
rect 90916 38344 90968 38350
rect 90916 38286 90968 38292
rect 90548 37392 90600 37398
rect 90548 37334 90600 37340
rect 90732 37392 90784 37398
rect 90732 37334 90784 37340
rect 90640 34400 90692 34406
rect 90640 34342 90692 34348
rect 90652 33114 90680 34342
rect 90640 33108 90692 33114
rect 90640 33050 90692 33056
rect 90824 32972 90876 32978
rect 90824 32914 90876 32920
rect 90640 31816 90692 31822
rect 90640 31758 90692 31764
rect 90456 26580 90508 26586
rect 90456 26522 90508 26528
rect 90456 25288 90508 25294
rect 90456 25230 90508 25236
rect 90180 24336 90232 24342
rect 90180 24278 90232 24284
rect 90192 23594 90220 24278
rect 90180 23588 90232 23594
rect 90180 23530 90232 23536
rect 90088 23248 90140 23254
rect 90088 23190 90140 23196
rect 89916 16546 90036 16574
rect 89732 9654 89760 16546
rect 89812 15360 89864 15366
rect 89812 15302 89864 15308
rect 89824 14278 89852 15302
rect 89812 14272 89864 14278
rect 89812 14214 89864 14220
rect 89720 9648 89772 9654
rect 89720 9590 89772 9596
rect 88984 9036 89036 9042
rect 88984 8978 89036 8984
rect 89352 9036 89404 9042
rect 89352 8978 89404 8984
rect 89364 5642 89392 8978
rect 89732 8838 89760 9590
rect 89720 8832 89772 8838
rect 89720 8774 89772 8780
rect 89352 5636 89404 5642
rect 89352 5578 89404 5584
rect 89812 5024 89864 5030
rect 89812 4966 89864 4972
rect 89076 4684 89128 4690
rect 89076 4626 89128 4632
rect 89720 4684 89772 4690
rect 89720 4626 89772 4632
rect 88892 2644 88944 2650
rect 88892 2586 88944 2592
rect 88800 2508 88852 2514
rect 88800 2450 88852 2456
rect 88892 2304 88944 2310
rect 88892 2246 88944 2252
rect 88904 800 88932 2246
rect 89088 800 89116 4626
rect 89352 4480 89404 4486
rect 89352 4422 89404 4428
rect 89364 3738 89392 4422
rect 89352 3732 89404 3738
rect 89352 3674 89404 3680
rect 89260 3460 89312 3466
rect 89260 3402 89312 3408
rect 89272 800 89300 3402
rect 89536 2100 89588 2106
rect 89536 2042 89588 2048
rect 89548 800 89576 2042
rect 89732 800 89760 4626
rect 89824 950 89852 4966
rect 89904 3664 89956 3670
rect 89904 3606 89956 3612
rect 89812 944 89864 950
rect 89812 886 89864 892
rect 89916 800 89944 3606
rect 90008 3194 90036 16546
rect 90192 15570 90220 23530
rect 90180 15564 90232 15570
rect 90180 15506 90232 15512
rect 90180 8016 90232 8022
rect 90180 7958 90232 7964
rect 89996 3188 90048 3194
rect 89996 3130 90048 3136
rect 90088 2916 90140 2922
rect 90088 2858 90140 2864
rect 90100 800 90128 2858
rect 90192 2650 90220 7958
rect 90468 5273 90496 25230
rect 90652 21418 90680 31758
rect 90836 24342 90864 32914
rect 90824 24336 90876 24342
rect 90824 24278 90876 24284
rect 90640 21412 90692 21418
rect 90640 21354 90692 21360
rect 90732 17536 90784 17542
rect 90732 17478 90784 17484
rect 90640 12640 90692 12646
rect 90640 12582 90692 12588
rect 90454 5264 90510 5273
rect 90454 5199 90510 5208
rect 90272 4684 90324 4690
rect 90272 4626 90324 4632
rect 90180 2644 90232 2650
rect 90180 2586 90232 2592
rect 90284 800 90312 4626
rect 90652 4146 90680 12582
rect 90744 9518 90772 17478
rect 90732 9512 90784 9518
rect 90732 9454 90784 9460
rect 90824 9512 90876 9518
rect 90824 9454 90876 9460
rect 90836 5370 90864 9454
rect 90824 5364 90876 5370
rect 90824 5306 90876 5312
rect 90822 5264 90878 5273
rect 90822 5199 90878 5208
rect 90836 5166 90864 5199
rect 90732 5160 90784 5166
rect 90732 5102 90784 5108
rect 90824 5160 90876 5166
rect 90824 5102 90876 5108
rect 90744 4554 90772 5102
rect 90732 4548 90784 4554
rect 90732 4490 90784 4496
rect 90640 4140 90692 4146
rect 90640 4082 90692 4088
rect 90548 3528 90600 3534
rect 90548 3470 90600 3476
rect 90560 800 90588 3470
rect 90824 2848 90876 2854
rect 90824 2790 90876 2796
rect 90836 1442 90864 2790
rect 90928 2650 90956 38286
rect 91572 35834 91600 39200
rect 92492 36718 92520 39200
rect 93124 38684 93176 38690
rect 93124 38626 93176 38632
rect 92480 36712 92532 36718
rect 92480 36654 92532 36660
rect 91560 35828 91612 35834
rect 91560 35770 91612 35776
rect 92112 34740 92164 34746
rect 92112 34682 92164 34688
rect 91744 31204 91796 31210
rect 91744 31146 91796 31152
rect 91836 31204 91888 31210
rect 91836 31146 91888 31152
rect 91466 27976 91522 27985
rect 91466 27911 91522 27920
rect 91284 25288 91336 25294
rect 91284 25230 91336 25236
rect 91296 24954 91324 25230
rect 91284 24948 91336 24954
rect 91284 24890 91336 24896
rect 91100 23112 91152 23118
rect 91100 23054 91152 23060
rect 91112 16574 91140 23054
rect 91192 18080 91244 18086
rect 91192 18022 91244 18028
rect 91204 17626 91232 18022
rect 91204 17598 91324 17626
rect 91112 16546 91232 16574
rect 91008 12436 91060 12442
rect 91008 12378 91060 12384
rect 91020 11830 91048 12378
rect 91008 11824 91060 11830
rect 91008 11766 91060 11772
rect 91100 4684 91152 4690
rect 91100 4626 91152 4632
rect 91112 3618 91140 4626
rect 91204 4078 91232 16546
rect 91296 7818 91324 17598
rect 91480 16574 91508 27911
rect 91652 27532 91704 27538
rect 91652 27474 91704 27480
rect 91664 26450 91692 27474
rect 91652 26444 91704 26450
rect 91652 26386 91704 26392
rect 91560 26376 91612 26382
rect 91560 26318 91612 26324
rect 91572 25974 91600 26318
rect 91560 25968 91612 25974
rect 91560 25910 91612 25916
rect 91480 16546 91692 16574
rect 91560 10804 91612 10810
rect 91560 10746 91612 10752
rect 91284 7812 91336 7818
rect 91284 7754 91336 7760
rect 91468 6860 91520 6866
rect 91468 6802 91520 6808
rect 91480 5710 91508 6802
rect 91468 5704 91520 5710
rect 91468 5646 91520 5652
rect 91480 5166 91508 5646
rect 91468 5160 91520 5166
rect 91468 5102 91520 5108
rect 91192 4072 91244 4078
rect 91192 4014 91244 4020
rect 91376 4072 91428 4078
rect 91376 4014 91428 4020
rect 91020 3590 91140 3618
rect 90916 2644 90968 2650
rect 90916 2586 90968 2592
rect 91020 2394 91048 3590
rect 91100 3528 91152 3534
rect 91100 3470 91152 3476
rect 90744 1414 90864 1442
rect 90928 2366 91048 2394
rect 90744 800 90772 1414
rect 90928 800 90956 2366
rect 91112 800 91140 3470
rect 91284 2440 91336 2446
rect 91284 2382 91336 2388
rect 91296 800 91324 2382
rect 91388 1358 91416 4014
rect 91572 2990 91600 10746
rect 91664 6914 91692 16546
rect 91756 15910 91784 31146
rect 91848 26450 91876 31146
rect 91836 26444 91888 26450
rect 91836 26386 91888 26392
rect 91928 26308 91980 26314
rect 91928 26250 91980 26256
rect 91940 24410 91968 26250
rect 91928 24404 91980 24410
rect 91928 24346 91980 24352
rect 91836 20052 91888 20058
rect 91836 19994 91888 20000
rect 91744 15904 91796 15910
rect 91744 15846 91796 15852
rect 91664 6886 91784 6914
rect 91652 4684 91704 4690
rect 91652 4626 91704 4632
rect 91560 2984 91612 2990
rect 91560 2926 91612 2932
rect 91664 2394 91692 4626
rect 91756 4162 91784 6886
rect 91848 5914 91876 19994
rect 91940 14550 91968 24346
rect 92020 16448 92072 16454
rect 92020 16390 92072 16396
rect 92032 14890 92060 16390
rect 92020 14884 92072 14890
rect 92020 14826 92072 14832
rect 91928 14544 91980 14550
rect 91928 14486 91980 14492
rect 91836 5908 91888 5914
rect 91836 5850 91888 5856
rect 91848 5098 91876 5850
rect 91836 5092 91888 5098
rect 91836 5034 91888 5040
rect 91756 4146 92060 4162
rect 91756 4140 92072 4146
rect 91756 4134 92020 4140
rect 91756 4010 91784 4134
rect 92020 4082 92072 4088
rect 91744 4004 91796 4010
rect 91744 3946 91796 3952
rect 91744 3664 91796 3670
rect 91744 3606 91796 3612
rect 91572 2366 91692 2394
rect 91376 1352 91428 1358
rect 91376 1294 91428 1300
rect 91572 800 91600 2366
rect 91756 800 91784 3606
rect 91928 2848 91980 2854
rect 91928 2790 91980 2796
rect 91940 800 91968 2790
rect 92124 2650 92152 34682
rect 92572 32020 92624 32026
rect 92572 31962 92624 31968
rect 92480 31884 92532 31890
rect 92480 31826 92532 31832
rect 92204 29844 92256 29850
rect 92204 29786 92256 29792
rect 92216 15162 92244 29786
rect 92492 28082 92520 31826
rect 92584 28150 92612 31962
rect 92664 30116 92716 30122
rect 92664 30058 92716 30064
rect 92676 28966 92704 30058
rect 92664 28960 92716 28966
rect 92664 28902 92716 28908
rect 92572 28144 92624 28150
rect 92572 28086 92624 28092
rect 92480 28076 92532 28082
rect 92480 28018 92532 28024
rect 92296 20256 92348 20262
rect 92296 20198 92348 20204
rect 92204 15156 92256 15162
rect 92204 15098 92256 15104
rect 92204 3120 92256 3126
rect 92204 3062 92256 3068
rect 92112 2644 92164 2650
rect 92112 2586 92164 2592
rect 92216 2530 92244 3062
rect 92308 2990 92336 20198
rect 92492 18766 92520 28018
rect 92480 18760 92532 18766
rect 92480 18702 92532 18708
rect 92492 18442 92520 18702
rect 92584 18578 92612 28086
rect 92676 20262 92704 28902
rect 92848 21956 92900 21962
rect 92848 21898 92900 21904
rect 92756 20800 92808 20806
rect 92756 20742 92808 20748
rect 92664 20256 92716 20262
rect 92664 20198 92716 20204
rect 92584 18550 92704 18578
rect 92492 18414 92612 18442
rect 92676 18426 92704 18550
rect 92480 18284 92532 18290
rect 92480 18226 92532 18232
rect 92492 18170 92520 18226
rect 92400 18142 92520 18170
rect 92400 16454 92428 18142
rect 92584 18034 92612 18414
rect 92664 18420 92716 18426
rect 92664 18362 92716 18368
rect 92492 18006 92612 18034
rect 92492 16574 92520 18006
rect 92492 16546 92612 16574
rect 92388 16448 92440 16454
rect 92388 16390 92440 16396
rect 92388 15156 92440 15162
rect 92388 15098 92440 15104
rect 92400 14906 92428 15098
rect 92480 14952 92532 14958
rect 92400 14900 92480 14906
rect 92400 14894 92532 14900
rect 92400 14878 92520 14894
rect 92584 11558 92612 16546
rect 92572 11552 92624 11558
rect 92572 11494 92624 11500
rect 92676 11082 92704 18362
rect 92664 11076 92716 11082
rect 92664 11018 92716 11024
rect 92768 6914 92796 20742
rect 92860 20330 92888 21898
rect 92940 20936 92992 20942
rect 92940 20878 92992 20884
rect 92848 20324 92900 20330
rect 92848 20266 92900 20272
rect 92952 18290 92980 20878
rect 92940 18284 92992 18290
rect 92940 18226 92992 18232
rect 93136 15978 93164 38626
rect 93320 37398 93348 39200
rect 93584 38140 93636 38146
rect 93584 38082 93636 38088
rect 93308 37392 93360 37398
rect 93308 37334 93360 37340
rect 93492 37324 93544 37330
rect 93492 37266 93544 37272
rect 93216 33856 93268 33862
rect 93216 33798 93268 33804
rect 93228 25702 93256 33798
rect 93400 31272 93452 31278
rect 93400 31214 93452 31220
rect 93308 30184 93360 30190
rect 93308 30126 93360 30132
rect 93216 25696 93268 25702
rect 93216 25638 93268 25644
rect 93320 20602 93348 30126
rect 93412 23050 93440 31214
rect 93400 23044 93452 23050
rect 93400 22986 93452 22992
rect 93308 20596 93360 20602
rect 93308 20538 93360 20544
rect 93124 15972 93176 15978
rect 93124 15914 93176 15920
rect 92492 6886 92796 6914
rect 92388 4072 92440 4078
rect 92388 4014 92440 4020
rect 92296 2984 92348 2990
rect 92296 2926 92348 2932
rect 92124 2502 92244 2530
rect 92124 800 92152 2502
rect 92400 800 92428 4014
rect 87144 128 87196 134
rect 87144 70 87196 76
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88522 0 88578 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89258 0 89314 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92386 0 92442 800
rect 92492 406 92520 6886
rect 93504 6458 93532 37266
rect 93596 31142 93624 38082
rect 94136 37324 94188 37330
rect 94136 37266 94188 37272
rect 93860 36780 93912 36786
rect 93860 36722 93912 36728
rect 93872 36242 93900 36722
rect 93860 36236 93912 36242
rect 93860 36178 93912 36184
rect 94044 36168 94096 36174
rect 94044 36110 94096 36116
rect 93860 31748 93912 31754
rect 93860 31690 93912 31696
rect 93872 31346 93900 31690
rect 93860 31340 93912 31346
rect 93860 31282 93912 31288
rect 93952 31340 94004 31346
rect 93952 31282 94004 31288
rect 93964 31226 93992 31282
rect 93872 31210 93992 31226
rect 93860 31204 93992 31210
rect 93912 31198 93992 31204
rect 93860 31146 93912 31152
rect 93584 31136 93636 31142
rect 93584 31078 93636 31084
rect 94056 29646 94084 36110
rect 94044 29640 94096 29646
rect 94044 29582 94096 29588
rect 93860 21548 93912 21554
rect 93860 21490 93912 21496
rect 93584 21004 93636 21010
rect 93584 20946 93636 20952
rect 93596 20806 93624 20946
rect 93584 20800 93636 20806
rect 93584 20742 93636 20748
rect 93676 20392 93728 20398
rect 93676 20334 93728 20340
rect 93688 12238 93716 20334
rect 93872 15162 93900 21490
rect 93952 20528 94004 20534
rect 93952 20470 94004 20476
rect 93964 20398 93992 20470
rect 93952 20392 94004 20398
rect 93952 20334 94004 20340
rect 93952 18624 94004 18630
rect 93952 18566 94004 18572
rect 93964 17338 93992 18566
rect 93952 17332 94004 17338
rect 93952 17274 94004 17280
rect 94044 16516 94096 16522
rect 94044 16458 94096 16464
rect 93860 15156 93912 15162
rect 93860 15098 93912 15104
rect 93952 13184 94004 13190
rect 93952 13126 94004 13132
rect 93676 12232 93728 12238
rect 93676 12174 93728 12180
rect 93492 6452 93544 6458
rect 93492 6394 93544 6400
rect 92940 5160 92992 5166
rect 92940 5102 92992 5108
rect 92756 4684 92808 4690
rect 92756 4626 92808 4632
rect 92664 2508 92716 2514
rect 92664 2450 92716 2456
rect 92572 2372 92624 2378
rect 92572 2314 92624 2320
rect 92584 800 92612 2314
rect 92676 1086 92704 2450
rect 92664 1080 92716 1086
rect 92664 1022 92716 1028
rect 92768 800 92796 4626
rect 92952 3126 92980 5102
rect 93860 4684 93912 4690
rect 93860 4626 93912 4632
rect 93584 4072 93636 4078
rect 93584 4014 93636 4020
rect 93032 3528 93084 3534
rect 93032 3470 93084 3476
rect 92940 3120 92992 3126
rect 92940 3062 92992 3068
rect 92848 2848 92900 2854
rect 92848 2790 92900 2796
rect 92480 400 92532 406
rect 92480 342 92532 348
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 92860 338 92888 2790
rect 93044 1850 93072 3470
rect 93124 2916 93176 2922
rect 93124 2858 93176 2864
rect 93400 2916 93452 2922
rect 93400 2858 93452 2864
rect 92952 1822 93072 1850
rect 92952 800 92980 1822
rect 93136 800 93164 2858
rect 93308 2304 93360 2310
rect 93308 2246 93360 2252
rect 93320 2106 93348 2246
rect 93308 2100 93360 2106
rect 93308 2042 93360 2048
rect 93412 800 93440 2858
rect 93596 800 93624 4014
rect 93872 2922 93900 4626
rect 93964 2990 93992 13126
rect 93952 2984 94004 2990
rect 93952 2926 94004 2932
rect 93860 2916 93912 2922
rect 93860 2858 93912 2864
rect 93768 2848 93820 2854
rect 93768 2790 93820 2796
rect 93780 800 93808 2790
rect 94056 2582 94084 16458
rect 94148 16153 94176 37266
rect 94240 36854 94268 39200
rect 94228 36848 94280 36854
rect 94228 36790 94280 36796
rect 95068 36242 95096 39200
rect 95988 37466 96016 39200
rect 96068 37800 96120 37806
rect 96068 37742 96120 37748
rect 95976 37460 96028 37466
rect 95976 37402 96028 37408
rect 96080 37398 96108 37742
rect 96068 37392 96120 37398
rect 96068 37334 96120 37340
rect 95240 37324 95292 37330
rect 95240 37266 95292 37272
rect 94596 36236 94648 36242
rect 94596 36178 94648 36184
rect 95056 36236 95108 36242
rect 95056 36178 95108 36184
rect 94228 34536 94280 34542
rect 94228 34478 94280 34484
rect 94240 16574 94268 34478
rect 94504 31476 94556 31482
rect 94504 31418 94556 31424
rect 94320 31204 94372 31210
rect 94320 31146 94372 31152
rect 94332 27062 94360 31146
rect 94412 27328 94464 27334
rect 94412 27270 94464 27276
rect 94320 27056 94372 27062
rect 94320 26998 94372 27004
rect 94320 17536 94372 17542
rect 94320 17478 94372 17484
rect 94332 17338 94360 17478
rect 94320 17332 94372 17338
rect 94320 17274 94372 17280
rect 94424 16574 94452 27270
rect 94516 26926 94544 31418
rect 94504 26920 94556 26926
rect 94504 26862 94556 26868
rect 94608 20534 94636 36178
rect 95252 35834 95280 37266
rect 96380 37020 96676 37040
rect 96436 37018 96460 37020
rect 96516 37018 96540 37020
rect 96596 37018 96620 37020
rect 96458 36966 96460 37018
rect 96522 36966 96534 37018
rect 96596 36966 96598 37018
rect 96436 36964 96460 36966
rect 96516 36964 96540 36966
rect 96596 36964 96620 36966
rect 96380 36944 96676 36964
rect 96816 36854 96844 39200
rect 97632 37732 97684 37738
rect 97632 37674 97684 37680
rect 97644 37466 97672 37674
rect 97632 37460 97684 37466
rect 97632 37402 97684 37408
rect 96804 36848 96856 36854
rect 96804 36790 96856 36796
rect 97630 36680 97686 36689
rect 97630 36615 97632 36624
rect 97684 36615 97686 36624
rect 97632 36586 97684 36592
rect 96620 36576 96672 36582
rect 96620 36518 96672 36524
rect 96632 36378 96660 36518
rect 96620 36372 96672 36378
rect 96620 36314 96672 36320
rect 97736 36242 97764 39200
rect 98564 37398 98592 39200
rect 98552 37392 98604 37398
rect 98552 37334 98604 37340
rect 99484 36854 99512 39200
rect 99472 36848 99524 36854
rect 99472 36790 99524 36796
rect 97724 36236 97776 36242
rect 97724 36178 97776 36184
rect 96380 35932 96676 35952
rect 96436 35930 96460 35932
rect 96516 35930 96540 35932
rect 96596 35930 96620 35932
rect 96458 35878 96460 35930
rect 96522 35878 96534 35930
rect 96596 35878 96598 35930
rect 96436 35876 96460 35878
rect 96516 35876 96540 35878
rect 96596 35876 96620 35878
rect 96380 35856 96676 35876
rect 95240 35828 95292 35834
rect 95240 35770 95292 35776
rect 96712 35284 96764 35290
rect 96712 35226 96764 35232
rect 94964 35148 95016 35154
rect 94964 35090 95016 35096
rect 94688 30252 94740 30258
rect 94688 30194 94740 30200
rect 94700 23662 94728 30194
rect 94780 28484 94832 28490
rect 94780 28426 94832 28432
rect 94792 27062 94820 28426
rect 94780 27056 94832 27062
rect 94780 26998 94832 27004
rect 94688 23656 94740 23662
rect 94688 23598 94740 23604
rect 94596 20528 94648 20534
rect 94596 20470 94648 20476
rect 94240 16546 94360 16574
rect 94424 16546 94544 16574
rect 94134 16144 94190 16153
rect 94134 16079 94190 16088
rect 94136 9104 94188 9110
rect 94136 9046 94188 9052
rect 94148 8634 94176 9046
rect 94136 8628 94188 8634
rect 94136 8570 94188 8576
rect 94148 8362 94176 8570
rect 94136 8356 94188 8362
rect 94136 8298 94188 8304
rect 94228 4684 94280 4690
rect 94228 4626 94280 4632
rect 94136 4072 94188 4078
rect 94136 4014 94188 4020
rect 94044 2576 94096 2582
rect 94044 2518 94096 2524
rect 93952 2440 94004 2446
rect 93952 2382 94004 2388
rect 93964 800 93992 2382
rect 94148 800 94176 4014
rect 94240 2446 94268 4626
rect 94332 2446 94360 16546
rect 94412 6384 94464 6390
rect 94412 6326 94464 6332
rect 94424 3194 94452 6326
rect 94412 3188 94464 3194
rect 94412 3130 94464 3136
rect 94412 2984 94464 2990
rect 94412 2926 94464 2932
rect 94228 2440 94280 2446
rect 94228 2382 94280 2388
rect 94320 2440 94372 2446
rect 94320 2382 94372 2388
rect 94424 800 94452 2926
rect 94516 2650 94544 16546
rect 94976 14822 95004 35090
rect 95424 35080 95476 35086
rect 95424 35022 95476 35028
rect 95332 34944 95384 34950
rect 95332 34886 95384 34892
rect 95148 33992 95200 33998
rect 95148 33934 95200 33940
rect 95056 32360 95108 32366
rect 95056 32302 95108 32308
rect 94964 14816 95016 14822
rect 94964 14758 95016 14764
rect 94872 8832 94924 8838
rect 94872 8774 94924 8780
rect 94884 8566 94912 8774
rect 94872 8560 94924 8566
rect 94872 8502 94924 8508
rect 95068 3602 95096 32302
rect 95160 30258 95188 33934
rect 95148 30252 95200 30258
rect 95148 30194 95200 30200
rect 95148 29640 95200 29646
rect 95148 29582 95200 29588
rect 95160 26926 95188 29582
rect 95148 26920 95200 26926
rect 95148 26862 95200 26868
rect 95344 24274 95372 34886
rect 95436 34066 95464 35022
rect 95516 34944 95568 34950
rect 95516 34886 95568 34892
rect 95424 34060 95476 34066
rect 95424 34002 95476 34008
rect 95528 33046 95556 34886
rect 96380 34844 96676 34864
rect 96436 34842 96460 34844
rect 96516 34842 96540 34844
rect 96596 34842 96620 34844
rect 96458 34790 96460 34842
rect 96522 34790 96534 34842
rect 96596 34790 96598 34842
rect 96436 34788 96460 34790
rect 96516 34788 96540 34790
rect 96596 34788 96620 34790
rect 96380 34768 96676 34788
rect 96380 33756 96676 33776
rect 96436 33754 96460 33756
rect 96516 33754 96540 33756
rect 96596 33754 96620 33756
rect 96458 33702 96460 33754
rect 96522 33702 96534 33754
rect 96596 33702 96598 33754
rect 96436 33700 96460 33702
rect 96516 33700 96540 33702
rect 96596 33700 96620 33702
rect 96380 33680 96676 33700
rect 95516 33040 95568 33046
rect 95516 32982 95568 32988
rect 96380 32668 96676 32688
rect 96436 32666 96460 32668
rect 96516 32666 96540 32668
rect 96596 32666 96620 32668
rect 96458 32614 96460 32666
rect 96522 32614 96534 32666
rect 96596 32614 96598 32666
rect 96436 32612 96460 32614
rect 96516 32612 96540 32614
rect 96596 32612 96620 32614
rect 96380 32592 96676 32612
rect 95884 32224 95936 32230
rect 95884 32166 95936 32172
rect 95896 31890 95924 32166
rect 95884 31884 95936 31890
rect 95884 31826 95936 31832
rect 96068 31816 96120 31822
rect 96068 31758 96120 31764
rect 95884 29300 95936 29306
rect 95884 29242 95936 29248
rect 95332 24268 95384 24274
rect 95332 24210 95384 24216
rect 95792 22772 95844 22778
rect 95792 22714 95844 22720
rect 95148 20528 95200 20534
rect 95148 20470 95200 20476
rect 95160 9042 95188 20470
rect 95516 9580 95568 9586
rect 95516 9522 95568 9528
rect 95528 9110 95556 9522
rect 95516 9104 95568 9110
rect 95516 9046 95568 9052
rect 95148 9036 95200 9042
rect 95148 8978 95200 8984
rect 95332 5772 95384 5778
rect 95332 5714 95384 5720
rect 95344 5574 95372 5714
rect 95332 5568 95384 5574
rect 95332 5510 95384 5516
rect 95700 5160 95752 5166
rect 95700 5102 95752 5108
rect 95240 5092 95292 5098
rect 95240 5034 95292 5040
rect 95056 3596 95108 3602
rect 95056 3538 95108 3544
rect 94780 3528 94832 3534
rect 94780 3470 94832 3476
rect 94596 2848 94648 2854
rect 94596 2790 94648 2796
rect 94504 2644 94556 2650
rect 94504 2586 94556 2592
rect 94608 800 94636 2790
rect 94792 800 94820 3470
rect 94964 3460 95016 3466
rect 94964 3402 95016 3408
rect 94976 800 95004 3402
rect 95252 2802 95280 5034
rect 95332 4684 95384 4690
rect 95332 4626 95384 4632
rect 95344 2854 95372 4626
rect 95424 4072 95476 4078
rect 95424 4014 95476 4020
rect 95160 2774 95280 2802
rect 95332 2848 95384 2854
rect 95332 2790 95384 2796
rect 95160 800 95188 2774
rect 95436 800 95464 4014
rect 95608 2916 95660 2922
rect 95608 2858 95660 2864
rect 95620 800 95648 2858
rect 95712 1034 95740 5102
rect 95804 3194 95832 22714
rect 95896 22234 95924 29242
rect 95884 22228 95936 22234
rect 95884 22170 95936 22176
rect 95896 21078 95924 22170
rect 95884 21072 95936 21078
rect 95884 21014 95936 21020
rect 96080 16574 96108 31758
rect 96380 31580 96676 31600
rect 96436 31578 96460 31580
rect 96516 31578 96540 31580
rect 96596 31578 96620 31580
rect 96458 31526 96460 31578
rect 96522 31526 96534 31578
rect 96596 31526 96598 31578
rect 96436 31524 96460 31526
rect 96516 31524 96540 31526
rect 96596 31524 96620 31526
rect 96380 31504 96676 31524
rect 96380 30492 96676 30512
rect 96436 30490 96460 30492
rect 96516 30490 96540 30492
rect 96596 30490 96620 30492
rect 96458 30438 96460 30490
rect 96522 30438 96534 30490
rect 96596 30438 96598 30490
rect 96436 30436 96460 30438
rect 96516 30436 96540 30438
rect 96596 30436 96620 30438
rect 96380 30416 96676 30436
rect 96380 29404 96676 29424
rect 96436 29402 96460 29404
rect 96516 29402 96540 29404
rect 96596 29402 96620 29404
rect 96458 29350 96460 29402
rect 96522 29350 96534 29402
rect 96596 29350 96598 29402
rect 96436 29348 96460 29350
rect 96516 29348 96540 29350
rect 96596 29348 96620 29350
rect 96380 29328 96676 29348
rect 96380 28316 96676 28336
rect 96436 28314 96460 28316
rect 96516 28314 96540 28316
rect 96596 28314 96620 28316
rect 96458 28262 96460 28314
rect 96522 28262 96534 28314
rect 96596 28262 96598 28314
rect 96436 28260 96460 28262
rect 96516 28260 96540 28262
rect 96596 28260 96620 28262
rect 96380 28240 96676 28260
rect 96380 27228 96676 27248
rect 96436 27226 96460 27228
rect 96516 27226 96540 27228
rect 96596 27226 96620 27228
rect 96458 27174 96460 27226
rect 96522 27174 96534 27226
rect 96596 27174 96598 27226
rect 96436 27172 96460 27174
rect 96516 27172 96540 27174
rect 96596 27172 96620 27174
rect 96380 27152 96676 27172
rect 96380 26140 96676 26160
rect 96436 26138 96460 26140
rect 96516 26138 96540 26140
rect 96596 26138 96620 26140
rect 96458 26086 96460 26138
rect 96522 26086 96534 26138
rect 96596 26086 96598 26138
rect 96436 26084 96460 26086
rect 96516 26084 96540 26086
rect 96596 26084 96620 26086
rect 96380 26064 96676 26084
rect 96380 25052 96676 25072
rect 96436 25050 96460 25052
rect 96516 25050 96540 25052
rect 96596 25050 96620 25052
rect 96458 24998 96460 25050
rect 96522 24998 96534 25050
rect 96596 24998 96598 25050
rect 96436 24996 96460 24998
rect 96516 24996 96540 24998
rect 96596 24996 96620 24998
rect 96380 24976 96676 24996
rect 96380 23964 96676 23984
rect 96436 23962 96460 23964
rect 96516 23962 96540 23964
rect 96596 23962 96620 23964
rect 96458 23910 96460 23962
rect 96522 23910 96534 23962
rect 96596 23910 96598 23962
rect 96436 23908 96460 23910
rect 96516 23908 96540 23910
rect 96596 23908 96620 23910
rect 96380 23888 96676 23908
rect 96380 22876 96676 22896
rect 96436 22874 96460 22876
rect 96516 22874 96540 22876
rect 96596 22874 96620 22876
rect 96458 22822 96460 22874
rect 96522 22822 96534 22874
rect 96596 22822 96598 22874
rect 96436 22820 96460 22822
rect 96516 22820 96540 22822
rect 96596 22820 96620 22822
rect 96380 22800 96676 22820
rect 96380 21788 96676 21808
rect 96436 21786 96460 21788
rect 96516 21786 96540 21788
rect 96596 21786 96620 21788
rect 96458 21734 96460 21786
rect 96522 21734 96534 21786
rect 96596 21734 96598 21786
rect 96436 21732 96460 21734
rect 96516 21732 96540 21734
rect 96596 21732 96620 21734
rect 96380 21712 96676 21732
rect 96380 20700 96676 20720
rect 96436 20698 96460 20700
rect 96516 20698 96540 20700
rect 96596 20698 96620 20700
rect 96458 20646 96460 20698
rect 96522 20646 96534 20698
rect 96596 20646 96598 20698
rect 96436 20644 96460 20646
rect 96516 20644 96540 20646
rect 96596 20644 96620 20646
rect 96380 20624 96676 20644
rect 96380 19612 96676 19632
rect 96436 19610 96460 19612
rect 96516 19610 96540 19612
rect 96596 19610 96620 19612
rect 96458 19558 96460 19610
rect 96522 19558 96534 19610
rect 96596 19558 96598 19610
rect 96436 19556 96460 19558
rect 96516 19556 96540 19558
rect 96596 19556 96620 19558
rect 96380 19536 96676 19556
rect 96380 18524 96676 18544
rect 96436 18522 96460 18524
rect 96516 18522 96540 18524
rect 96596 18522 96620 18524
rect 96458 18470 96460 18522
rect 96522 18470 96534 18522
rect 96596 18470 96598 18522
rect 96436 18468 96460 18470
rect 96516 18468 96540 18470
rect 96596 18468 96620 18470
rect 96380 18448 96676 18468
rect 96380 17436 96676 17456
rect 96436 17434 96460 17436
rect 96516 17434 96540 17436
rect 96596 17434 96620 17436
rect 96458 17382 96460 17434
rect 96522 17382 96534 17434
rect 96596 17382 96598 17434
rect 96436 17380 96460 17382
rect 96516 17380 96540 17382
rect 96596 17380 96620 17382
rect 96380 17360 96676 17380
rect 95988 16546 96108 16574
rect 96724 16574 96752 35226
rect 97538 31240 97594 31249
rect 97538 31175 97594 31184
rect 96896 26920 96948 26926
rect 96896 26862 96948 26868
rect 97448 26920 97500 26926
rect 97448 26862 97500 26868
rect 96908 22506 96936 26862
rect 97460 25226 97488 26862
rect 97448 25220 97500 25226
rect 97448 25162 97500 25168
rect 96896 22500 96948 22506
rect 96896 22442 96948 22448
rect 97552 19990 97580 31175
rect 98092 29028 98144 29034
rect 98092 28970 98144 28976
rect 97908 28756 97960 28762
rect 97908 28698 97960 28704
rect 97816 26784 97868 26790
rect 97816 26726 97868 26732
rect 97630 20088 97686 20097
rect 97630 20023 97632 20032
rect 97684 20023 97686 20032
rect 97632 19994 97684 20000
rect 97540 19984 97592 19990
rect 97540 19926 97592 19932
rect 96986 18184 97042 18193
rect 96986 18119 97042 18128
rect 97000 16574 97028 18119
rect 96724 16546 96844 16574
rect 97000 16546 97120 16574
rect 95988 9081 96016 16546
rect 96380 16348 96676 16368
rect 96436 16346 96460 16348
rect 96516 16346 96540 16348
rect 96596 16346 96620 16348
rect 96458 16294 96460 16346
rect 96522 16294 96534 16346
rect 96596 16294 96598 16346
rect 96436 16292 96460 16294
rect 96516 16292 96540 16294
rect 96596 16292 96620 16294
rect 96380 16272 96676 16292
rect 96380 15260 96676 15280
rect 96436 15258 96460 15260
rect 96516 15258 96540 15260
rect 96596 15258 96620 15260
rect 96458 15206 96460 15258
rect 96522 15206 96534 15258
rect 96596 15206 96598 15258
rect 96436 15204 96460 15206
rect 96516 15204 96540 15206
rect 96596 15204 96620 15206
rect 96380 15184 96676 15204
rect 96252 14408 96304 14414
rect 96252 14350 96304 14356
rect 96712 14408 96764 14414
rect 96712 14350 96764 14356
rect 96264 14006 96292 14350
rect 96380 14172 96676 14192
rect 96436 14170 96460 14172
rect 96516 14170 96540 14172
rect 96596 14170 96620 14172
rect 96458 14118 96460 14170
rect 96522 14118 96534 14170
rect 96596 14118 96598 14170
rect 96436 14116 96460 14118
rect 96516 14116 96540 14118
rect 96596 14116 96620 14118
rect 96380 14096 96676 14116
rect 96252 14000 96304 14006
rect 96252 13942 96304 13948
rect 96724 13530 96752 14350
rect 96712 13524 96764 13530
rect 96712 13466 96764 13472
rect 96380 13084 96676 13104
rect 96436 13082 96460 13084
rect 96516 13082 96540 13084
rect 96596 13082 96620 13084
rect 96458 13030 96460 13082
rect 96522 13030 96534 13082
rect 96596 13030 96598 13082
rect 96436 13028 96460 13030
rect 96516 13028 96540 13030
rect 96596 13028 96620 13030
rect 96380 13008 96676 13028
rect 96380 11996 96676 12016
rect 96436 11994 96460 11996
rect 96516 11994 96540 11996
rect 96596 11994 96620 11996
rect 96458 11942 96460 11994
rect 96522 11942 96534 11994
rect 96596 11942 96598 11994
rect 96436 11940 96460 11942
rect 96516 11940 96540 11942
rect 96596 11940 96620 11942
rect 96380 11920 96676 11940
rect 96712 11552 96764 11558
rect 96712 11494 96764 11500
rect 96724 11218 96752 11494
rect 96712 11212 96764 11218
rect 96712 11154 96764 11160
rect 96380 10908 96676 10928
rect 96436 10906 96460 10908
rect 96516 10906 96540 10908
rect 96596 10906 96620 10908
rect 96458 10854 96460 10906
rect 96522 10854 96534 10906
rect 96596 10854 96598 10906
rect 96436 10852 96460 10854
rect 96516 10852 96540 10854
rect 96596 10852 96620 10854
rect 96380 10832 96676 10852
rect 96068 10464 96120 10470
rect 96068 10406 96120 10412
rect 95974 9072 96030 9081
rect 95974 9007 96030 9016
rect 95884 6792 95936 6798
rect 95884 6734 95936 6740
rect 95896 5914 95924 6734
rect 95884 5908 95936 5914
rect 95884 5850 95936 5856
rect 95976 4684 96028 4690
rect 95976 4626 96028 4632
rect 95792 3188 95844 3194
rect 95792 3130 95844 3136
rect 95804 2990 95832 3130
rect 95792 2984 95844 2990
rect 95792 2926 95844 2932
rect 95792 2508 95844 2514
rect 95792 2450 95844 2456
rect 95804 1154 95832 2450
rect 95792 1148 95844 1154
rect 95792 1090 95844 1096
rect 95712 1006 95832 1034
rect 95804 800 95832 1006
rect 95988 800 96016 4626
rect 96080 3194 96108 10406
rect 96380 9820 96676 9840
rect 96436 9818 96460 9820
rect 96516 9818 96540 9820
rect 96596 9818 96620 9820
rect 96458 9766 96460 9818
rect 96522 9766 96534 9818
rect 96596 9766 96598 9818
rect 96436 9764 96460 9766
rect 96516 9764 96540 9766
rect 96596 9764 96620 9766
rect 96380 9744 96676 9764
rect 96380 8732 96676 8752
rect 96436 8730 96460 8732
rect 96516 8730 96540 8732
rect 96596 8730 96620 8732
rect 96458 8678 96460 8730
rect 96522 8678 96534 8730
rect 96596 8678 96598 8730
rect 96436 8676 96460 8678
rect 96516 8676 96540 8678
rect 96596 8676 96620 8678
rect 96380 8656 96676 8676
rect 96380 7644 96676 7664
rect 96436 7642 96460 7644
rect 96516 7642 96540 7644
rect 96596 7642 96620 7644
rect 96458 7590 96460 7642
rect 96522 7590 96534 7642
rect 96596 7590 96598 7642
rect 96436 7588 96460 7590
rect 96516 7588 96540 7590
rect 96596 7588 96620 7590
rect 96380 7568 96676 7588
rect 96380 6556 96676 6576
rect 96436 6554 96460 6556
rect 96516 6554 96540 6556
rect 96596 6554 96620 6556
rect 96458 6502 96460 6554
rect 96522 6502 96534 6554
rect 96596 6502 96598 6554
rect 96436 6500 96460 6502
rect 96516 6500 96540 6502
rect 96596 6500 96620 6502
rect 96380 6480 96676 6500
rect 96252 5772 96304 5778
rect 96252 5714 96304 5720
rect 96160 5024 96212 5030
rect 96160 4966 96212 4972
rect 96172 3534 96200 4966
rect 96160 3528 96212 3534
rect 96160 3470 96212 3476
rect 96068 3188 96120 3194
rect 96068 3130 96120 3136
rect 96160 3052 96212 3058
rect 96160 2994 96212 3000
rect 96172 1442 96200 2994
rect 96264 1986 96292 5714
rect 96380 5468 96676 5488
rect 96436 5466 96460 5468
rect 96516 5466 96540 5468
rect 96596 5466 96620 5468
rect 96458 5414 96460 5466
rect 96522 5414 96534 5466
rect 96596 5414 96598 5466
rect 96436 5412 96460 5414
rect 96516 5412 96540 5414
rect 96596 5412 96620 5414
rect 96380 5392 96676 5412
rect 96712 4684 96764 4690
rect 96712 4626 96764 4632
rect 96380 4380 96676 4400
rect 96436 4378 96460 4380
rect 96516 4378 96540 4380
rect 96596 4378 96620 4380
rect 96458 4326 96460 4378
rect 96522 4326 96534 4378
rect 96596 4326 96598 4378
rect 96436 4324 96460 4326
rect 96516 4324 96540 4326
rect 96596 4324 96620 4326
rect 96380 4304 96676 4324
rect 96380 3292 96676 3312
rect 96436 3290 96460 3292
rect 96516 3290 96540 3292
rect 96596 3290 96620 3292
rect 96458 3238 96460 3290
rect 96522 3238 96534 3290
rect 96596 3238 96598 3290
rect 96436 3236 96460 3238
rect 96516 3236 96540 3238
rect 96596 3236 96620 3238
rect 96380 3216 96676 3236
rect 96380 2204 96676 2224
rect 96436 2202 96460 2204
rect 96516 2202 96540 2204
rect 96596 2202 96620 2204
rect 96458 2150 96460 2202
rect 96522 2150 96534 2202
rect 96596 2150 96598 2202
rect 96436 2148 96460 2150
rect 96516 2148 96540 2150
rect 96596 2148 96620 2150
rect 96380 2128 96676 2148
rect 96724 1986 96752 4626
rect 96816 3670 96844 16546
rect 96896 9988 96948 9994
rect 96896 9930 96948 9936
rect 96804 3664 96856 3670
rect 96804 3606 96856 3612
rect 96804 2984 96856 2990
rect 96804 2926 96856 2932
rect 96264 1958 96476 1986
rect 96172 1414 96292 1442
rect 96264 800 96292 1414
rect 96448 800 96476 1958
rect 96632 1958 96752 1986
rect 96632 800 96660 1958
rect 96816 800 96844 2926
rect 96908 2922 96936 9930
rect 96988 6248 97040 6254
rect 96988 6190 97040 6196
rect 96896 2916 96948 2922
rect 96896 2858 96948 2864
rect 97000 800 97028 6190
rect 97092 4146 97120 16546
rect 97172 15972 97224 15978
rect 97172 15914 97224 15920
rect 97184 14482 97212 15914
rect 97356 15904 97408 15910
rect 97356 15846 97408 15852
rect 97172 14476 97224 14482
rect 97172 14418 97224 14424
rect 97264 14272 97316 14278
rect 97264 14214 97316 14220
rect 97276 13938 97304 14214
rect 97264 13932 97316 13938
rect 97264 13874 97316 13880
rect 97368 13870 97396 15846
rect 97448 15020 97500 15026
rect 97448 14962 97500 14968
rect 97460 14074 97488 14962
rect 97448 14068 97500 14074
rect 97448 14010 97500 14016
rect 97356 13864 97408 13870
rect 97356 13806 97408 13812
rect 97540 12096 97592 12102
rect 97540 12038 97592 12044
rect 97552 11354 97580 12038
rect 97540 11348 97592 11354
rect 97540 11290 97592 11296
rect 97724 7336 97776 7342
rect 97724 7278 97776 7284
rect 97632 6248 97684 6254
rect 97632 6190 97684 6196
rect 97540 4820 97592 4826
rect 97540 4762 97592 4768
rect 97264 4684 97316 4690
rect 97264 4626 97316 4632
rect 97080 4140 97132 4146
rect 97080 4082 97132 4088
rect 97276 800 97304 4626
rect 97448 3392 97500 3398
rect 97448 3334 97500 3340
rect 97460 800 97488 3334
rect 97552 2514 97580 4762
rect 97540 2508 97592 2514
rect 97540 2450 97592 2456
rect 97644 800 97672 6190
rect 97736 3058 97764 7278
rect 97828 6322 97856 26726
rect 97816 6316 97868 6322
rect 97816 6258 97868 6264
rect 97816 5160 97868 5166
rect 97816 5102 97868 5108
rect 97724 3052 97776 3058
rect 97724 2994 97776 3000
rect 97724 2848 97776 2854
rect 97724 2790 97776 2796
rect 97736 2582 97764 2790
rect 97724 2576 97776 2582
rect 97724 2518 97776 2524
rect 97828 800 97856 5102
rect 97920 4078 97948 28698
rect 98104 15065 98132 28970
rect 98368 19372 98420 19378
rect 98368 19314 98420 19320
rect 98090 15056 98146 15065
rect 98090 14991 98146 15000
rect 98276 6860 98328 6866
rect 98276 6802 98328 6808
rect 97908 4072 97960 4078
rect 97908 4014 97960 4020
rect 98000 3936 98052 3942
rect 98000 3878 98052 3884
rect 98012 800 98040 3878
rect 98288 800 98316 6802
rect 98380 2922 98408 19314
rect 99012 5772 99064 5778
rect 99012 5714 99064 5720
rect 98460 5092 98512 5098
rect 98460 5034 98512 5040
rect 98368 2916 98420 2922
rect 98368 2858 98420 2864
rect 98472 800 98500 5034
rect 98644 3460 98696 3466
rect 98644 3402 98696 3408
rect 98656 800 98684 3402
rect 98828 3052 98880 3058
rect 98828 2994 98880 3000
rect 98840 800 98868 2994
rect 99024 800 99052 5714
rect 99288 4004 99340 4010
rect 99288 3946 99340 3952
rect 99300 800 99328 3946
rect 99472 3528 99524 3534
rect 99472 3470 99524 3476
rect 99484 800 99512 3470
rect 99840 2848 99892 2854
rect 99840 2790 99892 2796
rect 99656 2372 99708 2378
rect 99656 2314 99708 2320
rect 99668 800 99696 2314
rect 99852 800 99880 2790
rect 92848 332 92900 338
rect 92848 274 92900 280
rect 92938 0 92994 800
rect 93122 0 93178 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95146 0 95202 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< via2 >>
rect 2502 29572 2558 29608
rect 2502 29552 2504 29572
rect 2504 29552 2556 29572
rect 2556 29552 2558 29572
rect 1398 20032 1454 20088
rect 2134 17720 2190 17776
rect 2686 7828 2688 7848
rect 2688 7828 2740 7848
rect 2740 7828 2742 7848
rect 2686 7792 2742 7828
rect 2226 720 2282 776
rect 3238 36780 3294 36816
rect 3238 36760 3240 36780
rect 3240 36760 3292 36780
rect 3292 36760 3294 36780
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 3238 9460 3240 9480
rect 3240 9460 3292 9480
rect 3292 9460 3294 9480
rect 3238 9424 3294 9460
rect 3054 6160 3110 6216
rect 2410 176 2466 232
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 5078 5516 5080 5536
rect 5080 5516 5132 5536
rect 5132 5516 5134 5536
rect 5078 5480 5134 5516
rect 5446 6296 5502 6352
rect 7654 5636 7710 5672
rect 7654 5616 7656 5636
rect 7656 5616 7708 5636
rect 7708 5616 7710 5636
rect 8758 5652 8760 5672
rect 8760 5652 8812 5672
rect 8812 5652 8814 5672
rect 8758 5616 8814 5652
rect 8482 5516 8484 5536
rect 8484 5516 8536 5536
rect 8536 5516 8538 5536
rect 8482 5480 8538 5516
rect 9954 21936 10010 21992
rect 10046 7928 10102 7984
rect 10874 18128 10930 18184
rect 11794 9036 11850 9072
rect 11794 9016 11796 9036
rect 11796 9016 11848 9036
rect 11848 9016 11850 9036
rect 13266 34584 13322 34640
rect 12346 11212 12402 11248
rect 12346 11192 12348 11212
rect 12348 11192 12400 11212
rect 12400 11192 12402 11212
rect 12530 11056 12586 11112
rect 12806 11192 12862 11248
rect 13082 11212 13138 11248
rect 13082 11192 13084 11212
rect 13084 11192 13136 11212
rect 13136 11192 13138 11212
rect 12162 7384 12218 7440
rect 15014 33904 15070 33960
rect 13818 25200 13874 25256
rect 14278 25200 14334 25256
rect 15658 28736 15714 28792
rect 16026 28736 16082 28792
rect 16026 11056 16082 11112
rect 17130 27956 17132 27976
rect 17132 27956 17184 27976
rect 17184 27956 17186 27976
rect 17130 27920 17186 27956
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 17590 33516 17646 33552
rect 17590 33496 17592 33516
rect 17592 33496 17644 33516
rect 17644 33496 17646 33516
rect 17222 3440 17278 3496
rect 17590 3612 17592 3632
rect 17592 3612 17644 3632
rect 17644 3612 17646 3632
rect 17590 3576 17646 3612
rect 17866 3304 17922 3360
rect 17498 1128 17554 1184
rect 18602 27956 18604 27976
rect 18604 27956 18656 27976
rect 18656 27956 18658 27976
rect 18602 27920 18658 27956
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 18970 31340 19026 31376
rect 18970 31320 18972 31340
rect 18972 31320 19024 31340
rect 19024 31320 19026 31340
rect 19614 31340 19670 31376
rect 19614 31320 19616 31340
rect 19616 31320 19668 31340
rect 19668 31320 19670 31340
rect 18878 28056 18934 28112
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19062 28056 19118 28112
rect 19154 27920 19210 27976
rect 18142 3612 18144 3632
rect 18144 3612 18196 3632
rect 18196 3612 18198 3632
rect 18142 3576 18198 3612
rect 18234 3460 18290 3496
rect 18234 3440 18236 3460
rect 18236 3440 18288 3460
rect 18288 3440 18290 3460
rect 18142 3340 18144 3360
rect 18144 3340 18196 3360
rect 18196 3340 18198 3360
rect 18142 3304 18198 3340
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19338 15000 19394 15056
rect 19522 15036 19524 15056
rect 19524 15036 19576 15056
rect 19576 15036 19578 15056
rect 19522 15000 19578 15036
rect 19430 14884 19486 14920
rect 19706 15000 19762 15056
rect 19430 14864 19432 14884
rect 19432 14864 19484 14884
rect 19484 14864 19486 14884
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19338 14592 19394 14648
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 20074 31048 20130 31104
rect 20350 28192 20406 28248
rect 20718 26460 20720 26480
rect 20720 26460 20772 26480
rect 20772 26460 20774 26480
rect 20718 26424 20774 26460
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 20534 14864 20590 14920
rect 20718 18536 20774 18592
rect 20718 15136 20774 15192
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 18878 5208 18934 5264
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19062 2896 19118 2952
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 20166 3712 20222 3768
rect 20074 2896 20130 2952
rect 20166 2624 20222 2680
rect 20350 6024 20406 6080
rect 21178 27784 21234 27840
rect 20626 3576 20682 3632
rect 20718 856 20774 912
rect 21546 27004 21548 27024
rect 21548 27004 21600 27024
rect 21600 27004 21602 27024
rect 21546 26968 21602 27004
rect 21546 26424 21602 26480
rect 22006 32972 22062 33008
rect 22006 32952 22008 32972
rect 22008 32952 22060 32972
rect 22060 32952 22062 32972
rect 22190 32988 22192 33008
rect 22192 32988 22244 33008
rect 22244 32988 22246 33008
rect 22190 32952 22246 32988
rect 22374 32292 22430 32328
rect 22374 32272 22376 32292
rect 22376 32272 22428 32292
rect 22428 32272 22430 32292
rect 21638 19236 21694 19272
rect 21638 19216 21640 19236
rect 21640 19216 21692 19236
rect 21692 19216 21694 19236
rect 21822 17856 21878 17912
rect 22282 27004 22284 27024
rect 22284 27004 22336 27024
rect 22336 27004 22338 27024
rect 22282 26968 22338 27004
rect 22466 20596 22522 20632
rect 22466 20576 22468 20596
rect 22468 20576 22520 20596
rect 22520 20576 22522 20596
rect 22466 20460 22522 20496
rect 22466 20440 22468 20460
rect 22468 20440 22520 20460
rect 22520 20440 22522 20460
rect 22466 19116 22468 19136
rect 22468 19116 22520 19136
rect 22520 19116 22522 19136
rect 22466 19080 22522 19116
rect 22466 13404 22468 13424
rect 22468 13404 22520 13424
rect 22520 13404 22522 13424
rect 22466 13368 22522 13404
rect 22742 19216 22798 19272
rect 23018 20596 23074 20632
rect 23018 20576 23020 20596
rect 23020 20576 23072 20596
rect 23072 20576 23074 20596
rect 23018 20460 23074 20496
rect 23018 20440 23020 20460
rect 23020 20440 23072 20460
rect 23072 20440 23074 20460
rect 23018 19080 23074 19136
rect 23018 18536 23074 18592
rect 21822 6704 21878 6760
rect 21822 6024 21878 6080
rect 21730 3440 21786 3496
rect 21178 2624 21234 2680
rect 21546 992 21602 1048
rect 22006 3304 22062 3360
rect 22282 3576 22338 3632
rect 24030 31628 24032 31648
rect 24032 31628 24084 31648
rect 24084 31628 24086 31648
rect 24030 31592 24086 31628
rect 24122 16532 24124 16552
rect 24124 16532 24176 16552
rect 24176 16532 24178 16552
rect 24122 16496 24178 16532
rect 24122 7112 24178 7168
rect 25042 19080 25098 19136
rect 24674 17856 24730 17912
rect 24766 7248 24822 7304
rect 25318 22888 25374 22944
rect 25226 18264 25282 18320
rect 25134 10240 25190 10296
rect 25594 17312 25650 17368
rect 26514 23296 26570 23352
rect 26330 23024 26386 23080
rect 25686 7284 25688 7304
rect 25688 7284 25740 7304
rect 25740 7284 25742 7304
rect 25686 7248 25742 7284
rect 25962 7284 25964 7304
rect 25964 7284 26016 7304
rect 26016 7284 26018 7304
rect 25962 7248 26018 7284
rect 25962 7148 25964 7168
rect 25964 7148 26016 7168
rect 26016 7148 26018 7168
rect 25962 7112 26018 7148
rect 25594 2760 25650 2816
rect 26514 16532 26516 16552
rect 26516 16532 26568 16552
rect 26568 16532 26570 16552
rect 26514 16496 26570 16532
rect 26330 10260 26386 10296
rect 26330 10240 26332 10260
rect 26332 10240 26384 10260
rect 26384 10240 26386 10260
rect 26974 32272 27030 32328
rect 26882 30776 26938 30832
rect 26882 23060 26884 23080
rect 26884 23060 26936 23080
rect 26936 23060 26938 23080
rect 26882 23024 26938 23060
rect 26882 17584 26938 17640
rect 27158 27396 27214 27432
rect 27158 27376 27160 27396
rect 27160 27376 27212 27396
rect 27212 27376 27214 27396
rect 27526 31592 27582 31648
rect 27526 31320 27582 31376
rect 26146 2896 26202 2952
rect 26422 3712 26478 3768
rect 28722 36116 28724 36136
rect 28724 36116 28776 36136
rect 28776 36116 28778 36136
rect 28722 36080 28778 36116
rect 27894 28192 27950 28248
rect 27802 26832 27858 26888
rect 28354 31356 28356 31376
rect 28356 31356 28408 31376
rect 28408 31356 28410 31376
rect 28354 31320 28410 31356
rect 28078 31184 28134 31240
rect 28170 31048 28226 31104
rect 28354 30812 28356 30832
rect 28356 30812 28408 30832
rect 28408 30812 28410 30832
rect 28354 30776 28410 30812
rect 27710 13404 27712 13424
rect 27712 13404 27764 13424
rect 27764 13404 27766 13424
rect 27710 13368 27766 13404
rect 28630 17620 28632 17640
rect 28632 17620 28684 17640
rect 28684 17620 28686 17640
rect 28630 17584 28686 17620
rect 29090 17992 29146 18048
rect 29090 17856 29146 17912
rect 30010 33380 30066 33416
rect 30010 33360 30012 33380
rect 30012 33360 30064 33380
rect 30064 33360 30066 33380
rect 30010 28600 30066 28656
rect 30194 33632 30250 33688
rect 30470 33260 30472 33280
rect 30472 33260 30524 33280
rect 30524 33260 30526 33280
rect 30470 33224 30526 33260
rect 30470 27376 30526 27432
rect 30470 26968 30526 27024
rect 30378 26580 30434 26616
rect 30378 26560 30380 26580
rect 30380 26560 30432 26580
rect 30432 26560 30434 26580
rect 30930 33360 30986 33416
rect 30378 24556 30380 24576
rect 30380 24556 30432 24576
rect 30432 24556 30434 24576
rect 30378 24520 30434 24556
rect 31298 30640 31354 30696
rect 31022 15988 31024 16008
rect 31024 15988 31076 16008
rect 31076 15988 31078 16008
rect 31022 15952 31078 15988
rect 31206 15680 31262 15736
rect 31390 16244 31446 16280
rect 31390 16224 31392 16244
rect 31392 16224 31444 16244
rect 31444 16224 31446 16244
rect 31390 16108 31446 16144
rect 31390 16088 31392 16108
rect 31392 16088 31444 16108
rect 31444 16088 31446 16108
rect 31482 15408 31538 15464
rect 31758 28056 31814 28112
rect 31758 16396 31760 16416
rect 31760 16396 31812 16416
rect 31812 16396 31814 16416
rect 31758 16360 31814 16396
rect 31758 16224 31814 16280
rect 31758 15952 31814 16008
rect 32034 16108 32090 16144
rect 32034 16088 32036 16108
rect 32036 16088 32088 16108
rect 32088 16088 32090 16108
rect 32034 15680 32090 15736
rect 32034 15408 32090 15464
rect 32494 22208 32550 22264
rect 33046 22108 33048 22128
rect 33048 22108 33100 22128
rect 33100 22108 33102 22128
rect 33046 22072 33102 22108
rect 33046 18264 33102 18320
rect 33322 26696 33378 26752
rect 33598 27784 33654 27840
rect 33230 10104 33286 10160
rect 33690 26460 33692 26480
rect 33692 26460 33744 26480
rect 33744 26460 33746 26480
rect 33690 26424 33746 26460
rect 33690 26324 33692 26344
rect 33692 26324 33744 26344
rect 33744 26324 33746 26344
rect 33690 26288 33746 26324
rect 33598 22636 33654 22672
rect 33598 22616 33600 22636
rect 33600 22616 33652 22636
rect 33652 22616 33654 22636
rect 33874 34448 33930 34504
rect 33874 30776 33930 30832
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34242 33652 34298 33688
rect 34242 33632 34244 33652
rect 34244 33632 34296 33652
rect 34296 33632 34298 33652
rect 33874 22636 33930 22672
rect 33874 22616 33876 22636
rect 33876 22616 33928 22636
rect 33928 22616 33930 22636
rect 33966 22344 34022 22400
rect 33690 20304 33746 20360
rect 33690 20032 33746 20088
rect 33690 19372 33746 19408
rect 33690 19352 33692 19372
rect 33692 19352 33744 19372
rect 33744 19352 33746 19372
rect 33598 18828 33654 18864
rect 33598 18808 33600 18828
rect 33600 18808 33652 18828
rect 33652 18808 33654 18828
rect 33414 18672 33470 18728
rect 33506 18400 33562 18456
rect 33598 18264 33654 18320
rect 33506 17176 33562 17232
rect 33690 14864 33746 14920
rect 34058 19896 34114 19952
rect 27434 448 27490 504
rect 34242 18944 34298 19000
rect 34150 18400 34206 18456
rect 34058 16124 34060 16144
rect 34060 16124 34112 16144
rect 34112 16124 34114 16144
rect 34058 16088 34114 16124
rect 34426 19080 34482 19136
rect 34426 17076 34428 17096
rect 34428 17076 34480 17096
rect 34480 17076 34482 17096
rect 34426 17040 34482 17076
rect 35990 35400 36046 35456
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34702 20324 34758 20360
rect 34702 20304 34704 20324
rect 34704 20304 34756 20324
rect 34756 20304 34758 20324
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34702 19080 34758 19136
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 35162 18264 35218 18320
rect 35346 18264 35402 18320
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 35162 17212 35164 17232
rect 35164 17212 35216 17232
rect 35216 17212 35218 17232
rect 35162 17176 35218 17212
rect 34702 16360 34758 16416
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34794 11464 34850 11520
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 33046 584 33102 640
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 35346 12416 35402 12472
rect 35714 29416 35770 29472
rect 35898 27548 35900 27568
rect 35900 27548 35952 27568
rect 35952 27548 35954 27568
rect 35898 27512 35954 27548
rect 36266 30776 36322 30832
rect 36174 28192 36230 28248
rect 36082 26832 36138 26888
rect 35806 25744 35862 25800
rect 35530 12280 35586 12336
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 35898 17040 35954 17096
rect 36358 26968 36414 27024
rect 36450 26560 36506 26616
rect 36082 19252 36084 19272
rect 36084 19252 36136 19272
rect 36136 19252 36138 19272
rect 36082 19216 36138 19252
rect 36726 26460 36728 26480
rect 36728 26460 36780 26480
rect 36780 26460 36782 26480
rect 36726 26424 36782 26460
rect 36726 26324 36728 26344
rect 36728 26324 36780 26344
rect 36780 26324 36782 26344
rect 36726 26288 36782 26324
rect 36634 19372 36690 19408
rect 36634 19352 36636 19372
rect 36636 19352 36688 19372
rect 36688 19352 36690 19372
rect 36726 19236 36782 19272
rect 36726 19216 36728 19236
rect 36728 19216 36780 19236
rect 36780 19216 36782 19236
rect 36266 14864 36322 14920
rect 35990 9560 36046 9616
rect 36726 19080 36782 19136
rect 36634 18672 36690 18728
rect 36726 17992 36782 18048
rect 36450 10376 36506 10432
rect 37002 28464 37058 28520
rect 37278 35400 37334 35456
rect 37554 28620 37610 28656
rect 37554 28600 37556 28620
rect 37556 28600 37608 28620
rect 37608 28600 37610 28620
rect 37002 24520 37058 24576
rect 37738 28500 37740 28520
rect 37740 28500 37792 28520
rect 37792 28500 37794 28520
rect 37738 28464 37794 28500
rect 37186 10376 37242 10432
rect 37278 9560 37334 9616
rect 38014 33260 38016 33280
rect 38016 33260 38068 33280
rect 38068 33260 38070 33280
rect 38014 33224 38070 33260
rect 38198 34176 38254 34232
rect 37830 26560 37886 26616
rect 37646 22108 37648 22128
rect 37648 22108 37700 22128
rect 37700 22108 37702 22128
rect 37646 22072 37702 22108
rect 37830 21528 37886 21584
rect 37738 19896 37794 19952
rect 38658 34448 38714 34504
rect 38934 33088 38990 33144
rect 38658 32716 38660 32736
rect 38660 32716 38712 32736
rect 38712 32716 38714 32736
rect 38658 32680 38714 32716
rect 38566 29416 38622 29472
rect 39946 36488 40002 36544
rect 39670 35672 39726 35728
rect 39302 35572 39304 35592
rect 39304 35572 39356 35592
rect 39356 35572 39358 35592
rect 39302 35536 39358 35572
rect 39486 35128 39542 35184
rect 39578 32952 39634 33008
rect 39394 32852 39396 32872
rect 39396 32852 39448 32872
rect 39448 32852 39450 32872
rect 39394 32816 39450 32852
rect 38566 22344 38622 22400
rect 38474 22208 38530 22264
rect 38566 21528 38622 21584
rect 38198 19080 38254 19136
rect 37922 12144 37978 12200
rect 38014 11328 38070 11384
rect 37922 10920 37978 10976
rect 38198 10104 38254 10160
rect 38934 26696 38990 26752
rect 38566 20052 38622 20088
rect 38566 20032 38568 20052
rect 38568 20032 38620 20052
rect 38620 20032 38622 20052
rect 38658 19780 38714 19816
rect 38658 19760 38660 19780
rect 38660 19760 38712 19780
rect 38712 19760 38714 19780
rect 38750 19624 38806 19680
rect 38566 17856 38622 17912
rect 38658 12280 38714 12336
rect 38842 11872 38898 11928
rect 38566 11464 38622 11520
rect 39302 27648 39358 27704
rect 39946 33632 40002 33688
rect 40130 33360 40186 33416
rect 39946 32308 39948 32328
rect 39948 32308 40000 32328
rect 40000 32308 40002 32328
rect 39946 32272 40002 32308
rect 40038 27784 40094 27840
rect 39578 27532 39634 27568
rect 39578 27512 39580 27532
rect 39580 27512 39632 27532
rect 39632 27512 39634 27532
rect 39854 25880 39910 25936
rect 39118 19760 39174 19816
rect 38474 11328 38530 11384
rect 38658 11328 38714 11384
rect 38934 11328 38990 11384
rect 38750 11056 38806 11112
rect 38842 8064 38898 8120
rect 39302 17992 39358 18048
rect 39394 12144 39450 12200
rect 39854 18944 39910 19000
rect 40038 18944 40094 19000
rect 39762 18536 39818 18592
rect 40038 16668 40040 16688
rect 40040 16668 40092 16688
rect 40092 16668 40094 16688
rect 40038 16632 40094 16668
rect 39394 11328 39450 11384
rect 39578 10920 39634 10976
rect 40682 32680 40738 32736
rect 40590 28056 40646 28112
rect 40498 27240 40554 27296
rect 40498 26460 40500 26480
rect 40500 26460 40552 26480
rect 40552 26460 40554 26480
rect 40498 26424 40554 26460
rect 40498 25472 40554 25528
rect 40498 24692 40500 24712
rect 40500 24692 40552 24712
rect 40552 24692 40554 24712
rect 40498 24656 40554 24692
rect 40314 15580 40316 15600
rect 40316 15580 40368 15600
rect 40368 15580 40370 15600
rect 39486 8064 39542 8120
rect 38566 312 38622 368
rect 40314 15544 40370 15580
rect 40406 14320 40462 14376
rect 40406 13796 40462 13832
rect 40406 13776 40408 13796
rect 40408 13776 40460 13796
rect 40460 13776 40462 13796
rect 40866 33768 40922 33824
rect 41510 36488 41566 36544
rect 41418 36216 41474 36272
rect 41418 35536 41474 35592
rect 41326 35264 41382 35320
rect 41326 34992 41382 35048
rect 41510 34196 41566 34232
rect 41510 34176 41512 34196
rect 41512 34176 41564 34196
rect 41564 34176 41566 34196
rect 41326 33632 41382 33688
rect 41234 33088 41290 33144
rect 42154 36896 42210 36952
rect 42154 33088 42210 33144
rect 41970 32544 42026 32600
rect 41050 26288 41106 26344
rect 40958 26152 41014 26208
rect 40958 23976 41014 24032
rect 40958 18692 41014 18728
rect 40958 18672 40960 18692
rect 40960 18672 41012 18692
rect 41012 18672 41014 18692
rect 41510 28192 41566 28248
rect 41510 27532 41566 27568
rect 41510 27512 41512 27532
rect 41512 27512 41564 27532
rect 41564 27512 41566 27532
rect 42062 28464 42118 28520
rect 41510 26696 41566 26752
rect 41510 25472 41566 25528
rect 41418 25200 41474 25256
rect 41510 21412 41566 21448
rect 41510 21392 41512 21412
rect 41512 21392 41564 21412
rect 41564 21392 41566 21412
rect 41418 18400 41474 18456
rect 41050 15700 41106 15736
rect 41050 15680 41052 15700
rect 41052 15680 41104 15700
rect 41104 15680 41106 15700
rect 41142 13948 41144 13968
rect 41144 13948 41196 13968
rect 41196 13948 41198 13968
rect 41142 13912 41198 13948
rect 41418 17856 41474 17912
rect 41510 15564 41566 15600
rect 41510 15544 41512 15564
rect 41512 15544 41564 15564
rect 41564 15544 41566 15564
rect 41786 24384 41842 24440
rect 41786 17992 41842 18048
rect 41786 15700 41842 15736
rect 41786 15680 41788 15700
rect 41788 15680 41840 15700
rect 41840 15680 41842 15700
rect 42706 32544 42762 32600
rect 42430 28328 42486 28384
rect 42614 27512 42670 27568
rect 42522 27240 42578 27296
rect 42338 26288 42394 26344
rect 41694 12164 41750 12200
rect 41694 12144 41696 12164
rect 41696 12144 41748 12164
rect 41748 12144 41750 12164
rect 41142 10668 41198 10704
rect 41142 10648 41144 10668
rect 41144 10648 41196 10668
rect 41196 10648 41198 10668
rect 41694 10648 41750 10704
rect 41786 10548 41788 10568
rect 41788 10548 41840 10568
rect 41840 10548 41842 10568
rect 41786 10512 41842 10548
rect 42890 26324 42892 26344
rect 42892 26324 42944 26344
rect 42944 26324 42946 26344
rect 42890 26288 42946 26324
rect 42982 23724 43038 23760
rect 42982 23704 42984 23724
rect 42984 23704 43036 23724
rect 43036 23704 43038 23724
rect 42798 18672 42854 18728
rect 43350 36488 43406 36544
rect 43442 36352 43498 36408
rect 43626 35128 43682 35184
rect 43350 34856 43406 34912
rect 43718 33360 43774 33416
rect 43534 30504 43590 30560
rect 43350 29960 43406 30016
rect 43350 29416 43406 29472
rect 43350 26560 43406 26616
rect 43258 25608 43314 25664
rect 43166 18944 43222 19000
rect 43534 28600 43590 28656
rect 43718 25608 43774 25664
rect 43626 25356 43682 25392
rect 43626 25336 43628 25356
rect 43628 25336 43680 25356
rect 43680 25336 43682 25356
rect 43718 25200 43774 25256
rect 43442 24792 43498 24848
rect 43534 24520 43590 24576
rect 43442 19624 43498 19680
rect 43442 19080 43498 19136
rect 43442 18300 43444 18320
rect 43444 18300 43496 18320
rect 43496 18300 43498 18320
rect 43442 18264 43498 18300
rect 44270 34992 44326 35048
rect 43994 33360 44050 33416
rect 44178 32272 44234 32328
rect 44086 27104 44142 27160
rect 43994 19760 44050 19816
rect 43902 19660 43904 19680
rect 43904 19660 43956 19680
rect 43956 19660 43958 19680
rect 43902 19624 43958 19660
rect 44086 19488 44142 19544
rect 44086 13932 44142 13968
rect 44086 13912 44088 13932
rect 44088 13912 44140 13932
rect 44140 13912 44142 13932
rect 43534 12724 43536 12744
rect 43536 12724 43588 12744
rect 43588 12724 43590 12744
rect 43534 12688 43590 12724
rect 44270 13776 44326 13832
rect 44270 10648 44326 10704
rect 44086 10376 44142 10432
rect 43994 9988 44050 10024
rect 43994 9968 43996 9988
rect 43996 9968 44048 9988
rect 44048 9968 44050 9988
rect 44638 24828 44640 24848
rect 44640 24828 44692 24848
rect 44692 24828 44694 24848
rect 44638 24792 44694 24828
rect 47766 36488 47822 36544
rect 47398 36352 47454 36408
rect 46754 35708 46756 35728
rect 46756 35708 46808 35728
rect 46808 35708 46810 35728
rect 46754 35672 46810 35708
rect 45466 34040 45522 34096
rect 45466 32952 45522 33008
rect 44546 21392 44602 21448
rect 44638 18944 44694 19000
rect 44546 18536 44602 18592
rect 44822 19488 44878 19544
rect 44730 18672 44786 18728
rect 44638 10512 44694 10568
rect 45098 19388 45100 19408
rect 45100 19388 45152 19408
rect 45152 19388 45154 19408
rect 45098 19352 45154 19388
rect 46294 30776 46350 30832
rect 45926 29824 45982 29880
rect 45834 29688 45890 29744
rect 45374 23740 45376 23760
rect 45376 23740 45428 23760
rect 45428 23740 45430 23760
rect 45374 23704 45430 23740
rect 45466 17856 45522 17912
rect 46110 30096 46166 30152
rect 46018 27648 46074 27704
rect 46294 27124 46350 27160
rect 46294 27104 46296 27124
rect 46296 27104 46348 27124
rect 46348 27104 46350 27124
rect 45926 19624 45982 19680
rect 47306 35264 47362 35320
rect 46478 33768 46534 33824
rect 46570 32836 46626 32872
rect 46570 32816 46572 32836
rect 46572 32816 46624 32836
rect 46624 32816 46626 32836
rect 46662 30504 46718 30560
rect 46662 30096 46718 30152
rect 46662 26288 46718 26344
rect 46662 24384 46718 24440
rect 46110 19388 46112 19408
rect 46112 19388 46164 19408
rect 46164 19388 46166 19408
rect 46110 19352 46166 19388
rect 46110 18808 46166 18864
rect 46110 17992 46166 18048
rect 46294 18964 46350 19000
rect 46294 18944 46296 18964
rect 46296 18944 46348 18964
rect 46348 18944 46350 18964
rect 46386 17992 46442 18048
rect 46386 17856 46442 17912
rect 46202 12688 46258 12744
rect 46662 24112 46718 24168
rect 46570 16360 46626 16416
rect 46938 29960 46994 30016
rect 46846 28056 46902 28112
rect 47030 24656 47086 24712
rect 46938 24520 46994 24576
rect 46846 24384 46902 24440
rect 46938 23976 46994 24032
rect 47306 34076 47308 34096
rect 47308 34076 47360 34096
rect 47360 34076 47362 34096
rect 47306 34040 47362 34076
rect 47306 33088 47362 33144
rect 47214 32952 47270 33008
rect 47214 30776 47270 30832
rect 47306 29688 47362 29744
rect 47214 29452 47216 29472
rect 47216 29452 47268 29472
rect 47268 29452 47270 29472
rect 47214 29416 47270 29452
rect 47306 23044 47362 23080
rect 47306 23024 47308 23044
rect 47308 23024 47360 23044
rect 47360 23024 47362 23044
rect 46938 19488 46994 19544
rect 46938 18400 46994 18456
rect 46938 16652 46994 16688
rect 46938 16632 46940 16652
rect 46940 16632 46992 16652
rect 46992 16632 46994 16652
rect 46846 16360 46902 16416
rect 47122 19080 47178 19136
rect 47214 14320 47270 14376
rect 46570 10668 46626 10704
rect 46570 10648 46572 10668
rect 46572 10648 46624 10668
rect 46624 10648 46626 10668
rect 46662 9968 46718 10024
rect 46478 1264 46534 1320
rect 47582 29824 47638 29880
rect 48502 36896 48558 36952
rect 48410 36216 48466 36272
rect 49698 36624 49754 36680
rect 48594 35980 48596 36000
rect 48596 35980 48648 36000
rect 48648 35980 48650 36000
rect 48594 35944 48650 35980
rect 49882 34992 49938 35048
rect 49054 32952 49110 33008
rect 48410 31728 48466 31784
rect 48042 26152 48098 26208
rect 48686 27376 48742 27432
rect 48318 26424 48374 26480
rect 48042 23060 48044 23080
rect 48044 23060 48096 23080
rect 48096 23060 48098 23080
rect 48042 23024 48098 23060
rect 47398 7792 47454 7848
rect 48318 20304 48374 20360
rect 48318 19916 48374 19952
rect 48318 19896 48320 19916
rect 48320 19896 48372 19916
rect 48372 19896 48374 19916
rect 48042 12180 48044 12200
rect 48044 12180 48096 12200
rect 48096 12180 48098 12200
rect 48042 12144 48098 12180
rect 48686 18536 48742 18592
rect 48778 15564 48834 15600
rect 48778 15544 48780 15564
rect 48780 15544 48832 15564
rect 48832 15544 48834 15564
rect 49238 27240 49294 27296
rect 49422 28600 49478 28656
rect 49514 15952 49570 16008
rect 48870 7112 48926 7168
rect 49974 28092 49976 28112
rect 49976 28092 50028 28112
rect 50028 28092 50030 28112
rect 49974 28056 50030 28092
rect 50300 37562 50356 37564
rect 50380 37562 50436 37564
rect 50460 37562 50516 37564
rect 50540 37562 50596 37564
rect 50300 37510 50326 37562
rect 50326 37510 50356 37562
rect 50380 37510 50390 37562
rect 50390 37510 50436 37562
rect 50460 37510 50506 37562
rect 50506 37510 50516 37562
rect 50540 37510 50570 37562
rect 50570 37510 50596 37562
rect 50300 37508 50356 37510
rect 50380 37508 50436 37510
rect 50460 37508 50516 37510
rect 50540 37508 50596 37510
rect 50300 36474 50356 36476
rect 50380 36474 50436 36476
rect 50460 36474 50516 36476
rect 50540 36474 50596 36476
rect 50300 36422 50326 36474
rect 50326 36422 50356 36474
rect 50380 36422 50390 36474
rect 50390 36422 50436 36474
rect 50460 36422 50506 36474
rect 50506 36422 50516 36474
rect 50540 36422 50570 36474
rect 50570 36422 50596 36474
rect 50300 36420 50356 36422
rect 50380 36420 50436 36422
rect 50460 36420 50516 36422
rect 50540 36420 50596 36422
rect 50300 35386 50356 35388
rect 50380 35386 50436 35388
rect 50460 35386 50516 35388
rect 50540 35386 50596 35388
rect 50300 35334 50326 35386
rect 50326 35334 50356 35386
rect 50380 35334 50390 35386
rect 50390 35334 50436 35386
rect 50460 35334 50506 35386
rect 50506 35334 50516 35386
rect 50540 35334 50570 35386
rect 50570 35334 50596 35386
rect 50300 35332 50356 35334
rect 50380 35332 50436 35334
rect 50460 35332 50516 35334
rect 50540 35332 50596 35334
rect 50300 34298 50356 34300
rect 50380 34298 50436 34300
rect 50460 34298 50516 34300
rect 50540 34298 50596 34300
rect 50300 34246 50326 34298
rect 50326 34246 50356 34298
rect 50380 34246 50390 34298
rect 50390 34246 50436 34298
rect 50460 34246 50506 34298
rect 50506 34246 50516 34298
rect 50540 34246 50570 34298
rect 50570 34246 50596 34298
rect 50300 34244 50356 34246
rect 50380 34244 50436 34246
rect 50460 34244 50516 34246
rect 50540 34244 50596 34246
rect 50300 33210 50356 33212
rect 50380 33210 50436 33212
rect 50460 33210 50516 33212
rect 50540 33210 50596 33212
rect 50300 33158 50326 33210
rect 50326 33158 50356 33210
rect 50380 33158 50390 33210
rect 50390 33158 50436 33210
rect 50460 33158 50506 33210
rect 50506 33158 50516 33210
rect 50540 33158 50570 33210
rect 50570 33158 50596 33210
rect 50300 33156 50356 33158
rect 50380 33156 50436 33158
rect 50460 33156 50516 33158
rect 50540 33156 50596 33158
rect 50618 32680 50674 32736
rect 50300 32122 50356 32124
rect 50380 32122 50436 32124
rect 50460 32122 50516 32124
rect 50540 32122 50596 32124
rect 50300 32070 50326 32122
rect 50326 32070 50356 32122
rect 50380 32070 50390 32122
rect 50390 32070 50436 32122
rect 50460 32070 50506 32122
rect 50506 32070 50516 32122
rect 50540 32070 50570 32122
rect 50570 32070 50596 32122
rect 50300 32068 50356 32070
rect 50380 32068 50436 32070
rect 50460 32068 50516 32070
rect 50540 32068 50596 32070
rect 50986 34448 51042 34504
rect 51170 34448 51226 34504
rect 50894 34060 50950 34096
rect 50894 34040 50896 34060
rect 50896 34040 50948 34060
rect 50948 34040 50950 34060
rect 51078 33224 51134 33280
rect 51078 32680 51134 32736
rect 50986 32172 50988 32192
rect 50988 32172 51040 32192
rect 51040 32172 51042 32192
rect 50986 32136 51042 32172
rect 50300 31034 50356 31036
rect 50380 31034 50436 31036
rect 50460 31034 50516 31036
rect 50540 31034 50596 31036
rect 50300 30982 50326 31034
rect 50326 30982 50356 31034
rect 50380 30982 50390 31034
rect 50390 30982 50436 31034
rect 50460 30982 50506 31034
rect 50506 30982 50516 31034
rect 50540 30982 50570 31034
rect 50570 30982 50596 31034
rect 50300 30980 50356 30982
rect 50380 30980 50436 30982
rect 50460 30980 50516 30982
rect 50540 30980 50596 30982
rect 50300 29946 50356 29948
rect 50380 29946 50436 29948
rect 50460 29946 50516 29948
rect 50540 29946 50596 29948
rect 50300 29894 50326 29946
rect 50326 29894 50356 29946
rect 50380 29894 50390 29946
rect 50390 29894 50436 29946
rect 50460 29894 50506 29946
rect 50506 29894 50516 29946
rect 50540 29894 50570 29946
rect 50570 29894 50596 29946
rect 50300 29892 50356 29894
rect 50380 29892 50436 29894
rect 50460 29892 50516 29894
rect 50540 29892 50596 29894
rect 50300 28858 50356 28860
rect 50380 28858 50436 28860
rect 50460 28858 50516 28860
rect 50540 28858 50596 28860
rect 50300 28806 50326 28858
rect 50326 28806 50356 28858
rect 50380 28806 50390 28858
rect 50390 28806 50436 28858
rect 50460 28806 50506 28858
rect 50506 28806 50516 28858
rect 50540 28806 50570 28858
rect 50570 28806 50596 28858
rect 50300 28804 50356 28806
rect 50380 28804 50436 28806
rect 50460 28804 50516 28806
rect 50540 28804 50596 28806
rect 50300 27770 50356 27772
rect 50380 27770 50436 27772
rect 50460 27770 50516 27772
rect 50540 27770 50596 27772
rect 50300 27718 50326 27770
rect 50326 27718 50356 27770
rect 50380 27718 50390 27770
rect 50390 27718 50436 27770
rect 50460 27718 50506 27770
rect 50506 27718 50516 27770
rect 50540 27718 50570 27770
rect 50570 27718 50596 27770
rect 50300 27716 50356 27718
rect 50380 27716 50436 27718
rect 50460 27716 50516 27718
rect 50540 27716 50596 27718
rect 50710 27548 50712 27568
rect 50712 27548 50764 27568
rect 50764 27548 50766 27568
rect 50300 26682 50356 26684
rect 50380 26682 50436 26684
rect 50460 26682 50516 26684
rect 50540 26682 50596 26684
rect 50300 26630 50326 26682
rect 50326 26630 50356 26682
rect 50380 26630 50390 26682
rect 50390 26630 50436 26682
rect 50460 26630 50506 26682
rect 50506 26630 50516 26682
rect 50540 26630 50570 26682
rect 50570 26630 50596 26682
rect 50300 26628 50356 26630
rect 50380 26628 50436 26630
rect 50460 26628 50516 26630
rect 50540 26628 50596 26630
rect 50710 27512 50766 27548
rect 50710 27104 50766 27160
rect 49790 3712 49846 3768
rect 49790 3440 49846 3496
rect 50300 25594 50356 25596
rect 50380 25594 50436 25596
rect 50460 25594 50516 25596
rect 50540 25594 50596 25596
rect 50300 25542 50326 25594
rect 50326 25542 50356 25594
rect 50380 25542 50390 25594
rect 50390 25542 50436 25594
rect 50460 25542 50506 25594
rect 50506 25542 50516 25594
rect 50540 25542 50570 25594
rect 50570 25542 50596 25594
rect 50300 25540 50356 25542
rect 50380 25540 50436 25542
rect 50460 25540 50516 25542
rect 50540 25540 50596 25542
rect 50526 24812 50582 24848
rect 50526 24792 50528 24812
rect 50528 24792 50580 24812
rect 50580 24792 50582 24812
rect 50526 24676 50582 24712
rect 50526 24656 50528 24676
rect 50528 24656 50580 24676
rect 50580 24656 50582 24676
rect 50300 24506 50356 24508
rect 50380 24506 50436 24508
rect 50460 24506 50516 24508
rect 50540 24506 50596 24508
rect 50300 24454 50326 24506
rect 50326 24454 50356 24506
rect 50380 24454 50390 24506
rect 50390 24454 50436 24506
rect 50460 24454 50506 24506
rect 50506 24454 50516 24506
rect 50540 24454 50570 24506
rect 50570 24454 50596 24506
rect 50300 24452 50356 24454
rect 50380 24452 50436 24454
rect 50460 24452 50516 24454
rect 50540 24452 50596 24454
rect 50300 23418 50356 23420
rect 50380 23418 50436 23420
rect 50460 23418 50516 23420
rect 50540 23418 50596 23420
rect 50300 23366 50326 23418
rect 50326 23366 50356 23418
rect 50380 23366 50390 23418
rect 50390 23366 50436 23418
rect 50460 23366 50506 23418
rect 50506 23366 50516 23418
rect 50540 23366 50570 23418
rect 50570 23366 50596 23418
rect 50300 23364 50356 23366
rect 50380 23364 50436 23366
rect 50460 23364 50516 23366
rect 50540 23364 50596 23366
rect 50300 22330 50356 22332
rect 50380 22330 50436 22332
rect 50460 22330 50516 22332
rect 50540 22330 50596 22332
rect 50300 22278 50326 22330
rect 50326 22278 50356 22330
rect 50380 22278 50390 22330
rect 50390 22278 50436 22330
rect 50460 22278 50506 22330
rect 50506 22278 50516 22330
rect 50540 22278 50570 22330
rect 50570 22278 50596 22330
rect 50300 22276 50356 22278
rect 50380 22276 50436 22278
rect 50460 22276 50516 22278
rect 50540 22276 50596 22278
rect 50300 21242 50356 21244
rect 50380 21242 50436 21244
rect 50460 21242 50516 21244
rect 50540 21242 50596 21244
rect 50300 21190 50326 21242
rect 50326 21190 50356 21242
rect 50380 21190 50390 21242
rect 50390 21190 50436 21242
rect 50460 21190 50506 21242
rect 50506 21190 50516 21242
rect 50540 21190 50570 21242
rect 50570 21190 50596 21242
rect 50300 21188 50356 21190
rect 50380 21188 50436 21190
rect 50460 21188 50516 21190
rect 50540 21188 50596 21190
rect 50300 20154 50356 20156
rect 50380 20154 50436 20156
rect 50460 20154 50516 20156
rect 50540 20154 50596 20156
rect 50300 20102 50326 20154
rect 50326 20102 50356 20154
rect 50380 20102 50390 20154
rect 50390 20102 50436 20154
rect 50460 20102 50506 20154
rect 50506 20102 50516 20154
rect 50540 20102 50570 20154
rect 50570 20102 50596 20154
rect 50300 20100 50356 20102
rect 50380 20100 50436 20102
rect 50460 20100 50516 20102
rect 50540 20100 50596 20102
rect 50894 28600 50950 28656
rect 50986 28328 51042 28384
rect 51170 28328 51226 28384
rect 51078 27668 51134 27704
rect 51078 27648 51080 27668
rect 51080 27648 51132 27668
rect 51132 27648 51134 27668
rect 51446 27104 51502 27160
rect 50986 25608 51042 25664
rect 51262 25220 51318 25256
rect 51262 25200 51264 25220
rect 51264 25200 51316 25220
rect 51316 25200 51318 25220
rect 51354 24812 51410 24848
rect 51354 24792 51356 24812
rect 51356 24792 51408 24812
rect 51408 24792 51410 24812
rect 51170 23160 51226 23216
rect 50894 21528 50950 21584
rect 50894 20868 50950 20904
rect 50894 20848 50896 20868
rect 50896 20848 50948 20868
rect 50948 20848 50950 20868
rect 51170 20848 51226 20904
rect 50300 19066 50356 19068
rect 50380 19066 50436 19068
rect 50460 19066 50516 19068
rect 50540 19066 50596 19068
rect 50300 19014 50326 19066
rect 50326 19014 50356 19066
rect 50380 19014 50390 19066
rect 50390 19014 50436 19066
rect 50460 19014 50506 19066
rect 50506 19014 50516 19066
rect 50540 19014 50570 19066
rect 50570 19014 50596 19066
rect 50300 19012 50356 19014
rect 50380 19012 50436 19014
rect 50460 19012 50516 19014
rect 50540 19012 50596 19014
rect 50710 18808 50766 18864
rect 50802 18672 50858 18728
rect 50300 17978 50356 17980
rect 50380 17978 50436 17980
rect 50460 17978 50516 17980
rect 50540 17978 50596 17980
rect 50300 17926 50326 17978
rect 50326 17926 50356 17978
rect 50380 17926 50390 17978
rect 50390 17926 50436 17978
rect 50460 17926 50506 17978
rect 50506 17926 50516 17978
rect 50540 17926 50570 17978
rect 50570 17926 50596 17978
rect 50300 17924 50356 17926
rect 50380 17924 50436 17926
rect 50460 17924 50516 17926
rect 50540 17924 50596 17926
rect 50300 16890 50356 16892
rect 50380 16890 50436 16892
rect 50460 16890 50516 16892
rect 50540 16890 50596 16892
rect 50300 16838 50326 16890
rect 50326 16838 50356 16890
rect 50380 16838 50390 16890
rect 50390 16838 50436 16890
rect 50460 16838 50506 16890
rect 50506 16838 50516 16890
rect 50540 16838 50570 16890
rect 50570 16838 50596 16890
rect 50300 16836 50356 16838
rect 50380 16836 50436 16838
rect 50460 16836 50516 16838
rect 50540 16836 50596 16838
rect 50300 15802 50356 15804
rect 50380 15802 50436 15804
rect 50460 15802 50516 15804
rect 50540 15802 50596 15804
rect 50300 15750 50326 15802
rect 50326 15750 50356 15802
rect 50380 15750 50390 15802
rect 50390 15750 50436 15802
rect 50460 15750 50506 15802
rect 50506 15750 50516 15802
rect 50540 15750 50570 15802
rect 50570 15750 50596 15802
rect 50300 15748 50356 15750
rect 50380 15748 50436 15750
rect 50460 15748 50516 15750
rect 50540 15748 50596 15750
rect 50300 14714 50356 14716
rect 50380 14714 50436 14716
rect 50460 14714 50516 14716
rect 50540 14714 50596 14716
rect 50300 14662 50326 14714
rect 50326 14662 50356 14714
rect 50380 14662 50390 14714
rect 50390 14662 50436 14714
rect 50460 14662 50506 14714
rect 50506 14662 50516 14714
rect 50540 14662 50570 14714
rect 50570 14662 50596 14714
rect 50300 14660 50356 14662
rect 50380 14660 50436 14662
rect 50460 14660 50516 14662
rect 50540 14660 50596 14662
rect 50300 13626 50356 13628
rect 50380 13626 50436 13628
rect 50460 13626 50516 13628
rect 50540 13626 50596 13628
rect 50300 13574 50326 13626
rect 50326 13574 50356 13626
rect 50380 13574 50390 13626
rect 50390 13574 50436 13626
rect 50460 13574 50506 13626
rect 50506 13574 50516 13626
rect 50540 13574 50570 13626
rect 50570 13574 50596 13626
rect 50300 13572 50356 13574
rect 50380 13572 50436 13574
rect 50460 13572 50516 13574
rect 50540 13572 50596 13574
rect 50300 12538 50356 12540
rect 50380 12538 50436 12540
rect 50460 12538 50516 12540
rect 50540 12538 50596 12540
rect 50300 12486 50326 12538
rect 50326 12486 50356 12538
rect 50380 12486 50390 12538
rect 50390 12486 50436 12538
rect 50460 12486 50506 12538
rect 50506 12486 50516 12538
rect 50540 12486 50570 12538
rect 50570 12486 50596 12538
rect 50300 12484 50356 12486
rect 50380 12484 50436 12486
rect 50460 12484 50516 12486
rect 50540 12484 50596 12486
rect 50300 11450 50356 11452
rect 50380 11450 50436 11452
rect 50460 11450 50516 11452
rect 50540 11450 50596 11452
rect 50300 11398 50326 11450
rect 50326 11398 50356 11450
rect 50380 11398 50390 11450
rect 50390 11398 50436 11450
rect 50460 11398 50506 11450
rect 50506 11398 50516 11450
rect 50540 11398 50570 11450
rect 50570 11398 50596 11450
rect 50300 11396 50356 11398
rect 50380 11396 50436 11398
rect 50460 11396 50516 11398
rect 50540 11396 50596 11398
rect 50300 10362 50356 10364
rect 50380 10362 50436 10364
rect 50460 10362 50516 10364
rect 50540 10362 50596 10364
rect 50300 10310 50326 10362
rect 50326 10310 50356 10362
rect 50380 10310 50390 10362
rect 50390 10310 50436 10362
rect 50460 10310 50506 10362
rect 50506 10310 50516 10362
rect 50540 10310 50570 10362
rect 50570 10310 50596 10362
rect 50300 10308 50356 10310
rect 50380 10308 50436 10310
rect 50460 10308 50516 10310
rect 50540 10308 50596 10310
rect 50300 9274 50356 9276
rect 50380 9274 50436 9276
rect 50460 9274 50516 9276
rect 50540 9274 50596 9276
rect 50300 9222 50326 9274
rect 50326 9222 50356 9274
rect 50380 9222 50390 9274
rect 50390 9222 50436 9274
rect 50460 9222 50506 9274
rect 50506 9222 50516 9274
rect 50540 9222 50570 9274
rect 50570 9222 50596 9274
rect 50300 9220 50356 9222
rect 50380 9220 50436 9222
rect 50460 9220 50516 9222
rect 50540 9220 50596 9222
rect 51170 18808 51226 18864
rect 51078 14864 51134 14920
rect 50802 8508 50804 8528
rect 50804 8508 50856 8528
rect 50856 8508 50858 8528
rect 50802 8472 50858 8508
rect 51078 8492 51134 8528
rect 51078 8472 51080 8492
rect 51080 8472 51132 8492
rect 51132 8472 51134 8492
rect 50300 8186 50356 8188
rect 50380 8186 50436 8188
rect 50460 8186 50516 8188
rect 50540 8186 50596 8188
rect 50300 8134 50326 8186
rect 50326 8134 50356 8186
rect 50380 8134 50390 8186
rect 50390 8134 50436 8186
rect 50460 8134 50506 8186
rect 50506 8134 50516 8186
rect 50540 8134 50570 8186
rect 50570 8134 50596 8186
rect 50300 8132 50356 8134
rect 50380 8132 50436 8134
rect 50460 8132 50516 8134
rect 50540 8132 50596 8134
rect 50158 7148 50160 7168
rect 50160 7148 50212 7168
rect 50212 7148 50214 7168
rect 50158 7112 50214 7148
rect 50300 7098 50356 7100
rect 50380 7098 50436 7100
rect 50460 7098 50516 7100
rect 50540 7098 50596 7100
rect 50300 7046 50326 7098
rect 50326 7046 50356 7098
rect 50380 7046 50390 7098
rect 50390 7046 50436 7098
rect 50460 7046 50506 7098
rect 50506 7046 50516 7098
rect 50540 7046 50570 7098
rect 50570 7046 50596 7098
rect 50300 7044 50356 7046
rect 50380 7044 50436 7046
rect 50460 7044 50516 7046
rect 50540 7044 50596 7046
rect 50300 6010 50356 6012
rect 50380 6010 50436 6012
rect 50460 6010 50516 6012
rect 50540 6010 50596 6012
rect 50300 5958 50326 6010
rect 50326 5958 50356 6010
rect 50380 5958 50390 6010
rect 50390 5958 50436 6010
rect 50460 5958 50506 6010
rect 50506 5958 50516 6010
rect 50540 5958 50570 6010
rect 50570 5958 50596 6010
rect 50300 5956 50356 5958
rect 50380 5956 50436 5958
rect 50460 5956 50516 5958
rect 50540 5956 50596 5958
rect 50300 4922 50356 4924
rect 50380 4922 50436 4924
rect 50460 4922 50516 4924
rect 50540 4922 50596 4924
rect 50300 4870 50326 4922
rect 50326 4870 50356 4922
rect 50380 4870 50390 4922
rect 50390 4870 50436 4922
rect 50460 4870 50506 4922
rect 50506 4870 50516 4922
rect 50540 4870 50570 4922
rect 50570 4870 50596 4922
rect 50300 4868 50356 4870
rect 50380 4868 50436 4870
rect 50460 4868 50516 4870
rect 50540 4868 50596 4870
rect 50300 3834 50356 3836
rect 50380 3834 50436 3836
rect 50460 3834 50516 3836
rect 50540 3834 50596 3836
rect 50300 3782 50326 3834
rect 50326 3782 50356 3834
rect 50380 3782 50390 3834
rect 50390 3782 50436 3834
rect 50460 3782 50506 3834
rect 50506 3782 50516 3834
rect 50540 3782 50570 3834
rect 50570 3782 50596 3834
rect 50300 3780 50356 3782
rect 50380 3780 50436 3782
rect 50460 3780 50516 3782
rect 50540 3780 50596 3782
rect 50300 2746 50356 2748
rect 50380 2746 50436 2748
rect 50460 2746 50516 2748
rect 50540 2746 50596 2748
rect 50300 2694 50326 2746
rect 50326 2694 50356 2746
rect 50380 2694 50390 2746
rect 50390 2694 50436 2746
rect 50460 2694 50506 2746
rect 50506 2694 50516 2746
rect 50540 2694 50570 2746
rect 50570 2694 50596 2746
rect 50300 2692 50356 2694
rect 50380 2692 50436 2694
rect 50460 2692 50516 2694
rect 50540 2692 50596 2694
rect 51538 24692 51540 24712
rect 51540 24692 51592 24712
rect 51592 24692 51594 24712
rect 51538 24656 51594 24692
rect 51722 18808 51778 18864
rect 51814 9424 51870 9480
rect 51814 8780 51816 8800
rect 51816 8780 51868 8800
rect 51868 8780 51870 8800
rect 51814 8744 51870 8780
rect 52182 35164 52184 35184
rect 52184 35164 52236 35184
rect 52236 35164 52238 35184
rect 52182 35128 52238 35164
rect 52182 31592 52238 31648
rect 52090 25492 52146 25528
rect 52090 25472 52092 25492
rect 52092 25472 52144 25492
rect 52144 25472 52146 25492
rect 52274 30096 52330 30152
rect 52366 29552 52422 29608
rect 52550 26868 52552 26888
rect 52552 26868 52604 26888
rect 52604 26868 52606 26888
rect 52550 26832 52606 26868
rect 52550 26444 52606 26480
rect 52550 26424 52552 26444
rect 52552 26424 52604 26444
rect 52604 26424 52606 26444
rect 52274 18572 52276 18592
rect 52276 18572 52328 18592
rect 52328 18572 52330 18592
rect 52274 18536 52330 18572
rect 52642 19236 52698 19272
rect 52642 19216 52644 19236
rect 52644 19216 52696 19236
rect 52696 19216 52698 19236
rect 52366 6296 52422 6352
rect 52734 6296 52790 6352
rect 53838 30368 53894 30424
rect 53286 27240 53342 27296
rect 53102 19896 53158 19952
rect 53102 13932 53158 13968
rect 53102 13912 53104 13932
rect 53104 13912 53156 13932
rect 53156 13912 53158 13932
rect 53194 6296 53250 6352
rect 53930 27668 53986 27704
rect 53930 27648 53932 27668
rect 53932 27648 53984 27668
rect 53984 27648 53986 27668
rect 53746 27376 53802 27432
rect 53654 27240 53710 27296
rect 53838 26444 53894 26480
rect 53838 26424 53840 26444
rect 53840 26424 53892 26444
rect 53892 26424 53894 26444
rect 53654 25472 53710 25528
rect 54206 31592 54262 31648
rect 54206 30268 54208 30288
rect 54208 30268 54260 30288
rect 54260 30268 54262 30288
rect 54206 30232 54262 30268
rect 54114 28600 54170 28656
rect 54114 27240 54170 27296
rect 53746 20712 53802 20768
rect 54574 34448 54630 34504
rect 54482 33632 54538 33688
rect 53930 15408 53986 15464
rect 54850 36236 54906 36272
rect 54850 36216 54852 36236
rect 54852 36216 54904 36236
rect 54904 36216 54906 36236
rect 54758 35400 54814 35456
rect 54666 29960 54722 30016
rect 54574 25880 54630 25936
rect 54482 20576 54538 20632
rect 55034 34040 55090 34096
rect 55310 35672 55366 35728
rect 55310 35556 55366 35592
rect 55310 35536 55312 35556
rect 55312 35536 55364 35556
rect 55364 35536 55366 35556
rect 55310 34468 55366 34504
rect 55310 34448 55312 34468
rect 55312 34448 55364 34468
rect 55364 34448 55366 34468
rect 55310 33632 55366 33688
rect 55034 30368 55090 30424
rect 55034 27104 55090 27160
rect 55034 23160 55090 23216
rect 54758 20576 54814 20632
rect 55034 21528 55090 21584
rect 55310 29028 55366 29064
rect 55310 29008 55312 29028
rect 55312 29008 55364 29028
rect 55364 29008 55366 29028
rect 55862 36252 55864 36272
rect 55864 36252 55916 36272
rect 55916 36252 55918 36272
rect 55862 36216 55918 36252
rect 55954 35944 56010 36000
rect 55862 35536 55918 35592
rect 55770 35400 55826 35456
rect 55586 26560 55642 26616
rect 55862 20712 55918 20768
rect 55770 18808 55826 18864
rect 55862 15952 55918 16008
rect 55862 15544 55918 15600
rect 55770 15428 55826 15464
rect 55770 15408 55772 15428
rect 55772 15408 55824 15428
rect 55824 15408 55826 15428
rect 56138 32952 56194 33008
rect 56046 27240 56102 27296
rect 56230 26560 56286 26616
rect 56230 25608 56286 25664
rect 56138 20304 56194 20360
rect 57242 35672 57298 35728
rect 56782 35400 56838 35456
rect 56782 31592 56838 31648
rect 56598 30232 56654 30288
rect 57150 29960 57206 30016
rect 56690 29008 56746 29064
rect 56506 8744 56562 8800
rect 56874 25200 56930 25256
rect 57426 35128 57482 35184
rect 56874 13932 56930 13968
rect 56874 13912 56876 13932
rect 56876 13912 56928 13932
rect 56928 13912 56930 13932
rect 57978 32136 58034 32192
rect 57886 32000 57942 32056
rect 57518 31864 57574 31920
rect 58162 31884 58218 31920
rect 58162 31864 58164 31884
rect 58164 31864 58216 31884
rect 58216 31864 58218 31884
rect 57886 31728 57942 31784
rect 57518 26832 57574 26888
rect 57794 14900 57796 14920
rect 57796 14900 57848 14920
rect 57848 14900 57850 14920
rect 57794 14864 57850 14900
rect 58530 29552 58586 29608
rect 58622 20576 58678 20632
rect 58346 14900 58348 14920
rect 58348 14900 58400 14920
rect 58400 14900 58402 14920
rect 58346 14864 58402 14900
rect 58806 32000 58862 32056
rect 59818 36488 59874 36544
rect 59174 26988 59230 27024
rect 59174 26968 59176 26988
rect 59176 26968 59228 26988
rect 59228 26968 59230 26988
rect 59266 26560 59322 26616
rect 59726 31340 59782 31376
rect 59726 31320 59728 31340
rect 59728 31320 59780 31340
rect 59780 31320 59782 31340
rect 59358 19080 59414 19136
rect 59082 5072 59138 5128
rect 59266 8608 59322 8664
rect 61198 34992 61254 35048
rect 60370 33632 60426 33688
rect 60370 33224 60426 33280
rect 60738 33260 60740 33280
rect 60740 33260 60792 33280
rect 60792 33260 60794 33280
rect 60738 33224 60794 33260
rect 60646 31340 60702 31376
rect 60646 31320 60648 31340
rect 60648 31320 60700 31340
rect 60700 31320 60702 31340
rect 60646 26560 60702 26616
rect 60554 26460 60556 26480
rect 60556 26460 60608 26480
rect 60608 26460 60610 26480
rect 60554 26424 60610 26460
rect 60922 26968 60978 27024
rect 62026 35148 62082 35184
rect 62026 35128 62028 35148
rect 62028 35128 62080 35148
rect 62080 35128 62082 35148
rect 62578 34992 62634 35048
rect 61290 33632 61346 33688
rect 61474 33224 61530 33280
rect 63130 35128 63186 35184
rect 62670 33768 62726 33824
rect 61198 26424 61254 26480
rect 61014 22480 61070 22536
rect 60830 21664 60886 21720
rect 61106 21664 61162 21720
rect 60278 14340 60334 14376
rect 60278 14320 60280 14340
rect 60280 14320 60332 14340
rect 60332 14320 60334 14340
rect 60554 20868 60610 20904
rect 60554 20848 60556 20868
rect 60556 20848 60608 20868
rect 60608 20848 60610 20868
rect 60738 19488 60794 19544
rect 60738 19216 60794 19272
rect 60462 18264 60518 18320
rect 60830 19080 60886 19136
rect 60646 18536 60702 18592
rect 61290 21392 61346 21448
rect 61106 19488 61162 19544
rect 61106 19252 61108 19272
rect 61108 19252 61160 19272
rect 61160 19252 61162 19272
rect 61106 19216 61162 19252
rect 61014 14456 61070 14512
rect 60830 8628 60886 8664
rect 60830 8608 60832 8628
rect 60832 8608 60884 8628
rect 60884 8608 60886 8628
rect 60738 8472 60794 8528
rect 61106 14340 61162 14376
rect 61106 14320 61108 14340
rect 61108 14320 61160 14340
rect 61160 14320 61162 14340
rect 61474 23024 61530 23080
rect 61566 21428 61568 21448
rect 61568 21428 61620 21448
rect 61620 21428 61622 21448
rect 61566 21392 61622 21428
rect 61566 21256 61622 21312
rect 62026 25200 62082 25256
rect 62762 30132 62764 30152
rect 62764 30132 62816 30152
rect 62816 30132 62818 30152
rect 62762 30096 62818 30132
rect 62210 22480 62266 22536
rect 62210 18672 62266 18728
rect 61658 8900 61714 8936
rect 61658 8880 61660 8900
rect 61660 8880 61712 8900
rect 61712 8880 61714 8900
rect 61658 8608 61714 8664
rect 61750 4528 61806 4584
rect 62026 4700 62028 4720
rect 62028 4700 62080 4720
rect 62080 4700 62082 4720
rect 62026 4664 62082 4700
rect 62210 8472 62266 8528
rect 62394 14864 62450 14920
rect 62670 15544 62726 15600
rect 62394 9460 62396 9480
rect 62396 9460 62448 9480
rect 62448 9460 62450 9480
rect 62394 9424 62450 9460
rect 62026 4428 62028 4448
rect 62028 4428 62080 4448
rect 62080 4428 62082 4448
rect 62026 4392 62082 4428
rect 55494 720 55550 776
rect 62946 20576 63002 20632
rect 62946 11056 63002 11112
rect 62854 4548 62910 4584
rect 62854 4528 62856 4548
rect 62856 4528 62908 4548
rect 62908 4528 62910 4548
rect 63590 21292 63592 21312
rect 63592 21292 63644 21312
rect 63644 21292 63646 21312
rect 63590 21256 63646 21292
rect 64050 20304 64106 20360
rect 63314 8608 63370 8664
rect 63682 14476 63738 14512
rect 63682 14456 63684 14476
rect 63684 14456 63736 14476
rect 63736 14456 63738 14476
rect 64510 20476 64512 20496
rect 64512 20476 64564 20496
rect 64564 20476 64566 20496
rect 64510 20440 64566 20476
rect 64418 4664 64474 4720
rect 64786 20576 64842 20632
rect 64970 22752 65026 22808
rect 65660 37018 65716 37020
rect 65740 37018 65796 37020
rect 65820 37018 65876 37020
rect 65900 37018 65956 37020
rect 65660 36966 65686 37018
rect 65686 36966 65716 37018
rect 65740 36966 65750 37018
rect 65750 36966 65796 37018
rect 65820 36966 65866 37018
rect 65866 36966 65876 37018
rect 65900 36966 65930 37018
rect 65930 36966 65956 37018
rect 65660 36964 65716 36966
rect 65740 36964 65796 36966
rect 65820 36964 65876 36966
rect 65900 36964 65956 36966
rect 65062 22500 65118 22536
rect 65062 22480 65064 22500
rect 65064 22480 65116 22500
rect 65116 22480 65118 22500
rect 65798 36488 65854 36544
rect 65660 35930 65716 35932
rect 65740 35930 65796 35932
rect 65820 35930 65876 35932
rect 65900 35930 65956 35932
rect 65660 35878 65686 35930
rect 65686 35878 65716 35930
rect 65740 35878 65750 35930
rect 65750 35878 65796 35930
rect 65820 35878 65866 35930
rect 65866 35878 65876 35930
rect 65900 35878 65930 35930
rect 65930 35878 65956 35930
rect 65660 35876 65716 35878
rect 65740 35876 65796 35878
rect 65820 35876 65876 35878
rect 65900 35876 65956 35878
rect 65660 34842 65716 34844
rect 65740 34842 65796 34844
rect 65820 34842 65876 34844
rect 65900 34842 65956 34844
rect 65660 34790 65686 34842
rect 65686 34790 65716 34842
rect 65740 34790 65750 34842
rect 65750 34790 65796 34842
rect 65820 34790 65866 34842
rect 65866 34790 65876 34842
rect 65900 34790 65930 34842
rect 65930 34790 65956 34842
rect 65660 34788 65716 34790
rect 65740 34788 65796 34790
rect 65820 34788 65876 34790
rect 65900 34788 65956 34790
rect 65660 33754 65716 33756
rect 65740 33754 65796 33756
rect 65820 33754 65876 33756
rect 65900 33754 65956 33756
rect 65660 33702 65686 33754
rect 65686 33702 65716 33754
rect 65740 33702 65750 33754
rect 65750 33702 65796 33754
rect 65820 33702 65866 33754
rect 65866 33702 65876 33754
rect 65900 33702 65930 33754
rect 65930 33702 65956 33754
rect 65660 33700 65716 33702
rect 65740 33700 65796 33702
rect 65820 33700 65876 33702
rect 65900 33700 65956 33702
rect 65660 32666 65716 32668
rect 65740 32666 65796 32668
rect 65820 32666 65876 32668
rect 65900 32666 65956 32668
rect 65660 32614 65686 32666
rect 65686 32614 65716 32666
rect 65740 32614 65750 32666
rect 65750 32614 65796 32666
rect 65820 32614 65866 32666
rect 65866 32614 65876 32666
rect 65900 32614 65930 32666
rect 65930 32614 65956 32666
rect 65660 32612 65716 32614
rect 65740 32612 65796 32614
rect 65820 32612 65876 32614
rect 65900 32612 65956 32614
rect 65660 31578 65716 31580
rect 65740 31578 65796 31580
rect 65820 31578 65876 31580
rect 65900 31578 65956 31580
rect 65660 31526 65686 31578
rect 65686 31526 65716 31578
rect 65740 31526 65750 31578
rect 65750 31526 65796 31578
rect 65820 31526 65866 31578
rect 65866 31526 65876 31578
rect 65900 31526 65930 31578
rect 65930 31526 65956 31578
rect 65660 31524 65716 31526
rect 65740 31524 65796 31526
rect 65820 31524 65876 31526
rect 65900 31524 65956 31526
rect 65660 30490 65716 30492
rect 65740 30490 65796 30492
rect 65820 30490 65876 30492
rect 65900 30490 65956 30492
rect 65660 30438 65686 30490
rect 65686 30438 65716 30490
rect 65740 30438 65750 30490
rect 65750 30438 65796 30490
rect 65820 30438 65866 30490
rect 65866 30438 65876 30490
rect 65900 30438 65930 30490
rect 65930 30438 65956 30490
rect 65660 30436 65716 30438
rect 65740 30436 65796 30438
rect 65820 30436 65876 30438
rect 65900 30436 65956 30438
rect 65614 29552 65670 29608
rect 65660 29402 65716 29404
rect 65740 29402 65796 29404
rect 65820 29402 65876 29404
rect 65900 29402 65956 29404
rect 65660 29350 65686 29402
rect 65686 29350 65716 29402
rect 65740 29350 65750 29402
rect 65750 29350 65796 29402
rect 65820 29350 65866 29402
rect 65866 29350 65876 29402
rect 65900 29350 65930 29402
rect 65930 29350 65956 29402
rect 65660 29348 65716 29350
rect 65740 29348 65796 29350
rect 65820 29348 65876 29350
rect 65900 29348 65956 29350
rect 65660 28314 65716 28316
rect 65740 28314 65796 28316
rect 65820 28314 65876 28316
rect 65900 28314 65956 28316
rect 65660 28262 65686 28314
rect 65686 28262 65716 28314
rect 65740 28262 65750 28314
rect 65750 28262 65796 28314
rect 65820 28262 65866 28314
rect 65866 28262 65876 28314
rect 65900 28262 65930 28314
rect 65930 28262 65956 28314
rect 65660 28260 65716 28262
rect 65740 28260 65796 28262
rect 65820 28260 65876 28262
rect 65900 28260 65956 28262
rect 65660 27226 65716 27228
rect 65740 27226 65796 27228
rect 65820 27226 65876 27228
rect 65900 27226 65956 27228
rect 65660 27174 65686 27226
rect 65686 27174 65716 27226
rect 65740 27174 65750 27226
rect 65750 27174 65796 27226
rect 65820 27174 65866 27226
rect 65866 27174 65876 27226
rect 65900 27174 65930 27226
rect 65930 27174 65956 27226
rect 65660 27172 65716 27174
rect 65740 27172 65796 27174
rect 65820 27172 65876 27174
rect 65900 27172 65956 27174
rect 65246 22344 65302 22400
rect 65246 20340 65248 20360
rect 65248 20340 65300 20360
rect 65300 20340 65302 20360
rect 65246 20304 65302 20340
rect 65660 26138 65716 26140
rect 65740 26138 65796 26140
rect 65820 26138 65876 26140
rect 65900 26138 65956 26140
rect 65660 26086 65686 26138
rect 65686 26086 65716 26138
rect 65740 26086 65750 26138
rect 65750 26086 65796 26138
rect 65820 26086 65866 26138
rect 65866 26086 65876 26138
rect 65900 26086 65930 26138
rect 65930 26086 65956 26138
rect 65660 26084 65716 26086
rect 65740 26084 65796 26086
rect 65820 26084 65876 26086
rect 65900 26084 65956 26086
rect 65614 25220 65670 25256
rect 65614 25200 65616 25220
rect 65616 25200 65668 25220
rect 65668 25200 65670 25220
rect 65660 25050 65716 25052
rect 65740 25050 65796 25052
rect 65820 25050 65876 25052
rect 65900 25050 65956 25052
rect 65660 24998 65686 25050
rect 65686 24998 65716 25050
rect 65740 24998 65750 25050
rect 65750 24998 65796 25050
rect 65820 24998 65866 25050
rect 65866 24998 65876 25050
rect 65900 24998 65930 25050
rect 65930 24998 65956 25050
rect 65660 24996 65716 24998
rect 65740 24996 65796 24998
rect 65820 24996 65876 24998
rect 65900 24996 65956 24998
rect 65660 23962 65716 23964
rect 65740 23962 65796 23964
rect 65820 23962 65876 23964
rect 65900 23962 65956 23964
rect 65660 23910 65686 23962
rect 65686 23910 65716 23962
rect 65740 23910 65750 23962
rect 65750 23910 65796 23962
rect 65820 23910 65866 23962
rect 65866 23910 65876 23962
rect 65900 23910 65930 23962
rect 65930 23910 65956 23962
rect 65660 23908 65716 23910
rect 65740 23908 65796 23910
rect 65820 23908 65876 23910
rect 65900 23908 65956 23910
rect 65890 23024 65946 23080
rect 65660 22874 65716 22876
rect 65740 22874 65796 22876
rect 65820 22874 65876 22876
rect 65900 22874 65956 22876
rect 65660 22822 65686 22874
rect 65686 22822 65716 22874
rect 65740 22822 65750 22874
rect 65750 22822 65796 22874
rect 65820 22822 65866 22874
rect 65866 22822 65876 22874
rect 65900 22822 65930 22874
rect 65930 22822 65956 22874
rect 65660 22820 65716 22822
rect 65740 22820 65796 22822
rect 65820 22820 65876 22822
rect 65900 22820 65956 22822
rect 65660 21786 65716 21788
rect 65740 21786 65796 21788
rect 65820 21786 65876 21788
rect 65900 21786 65956 21788
rect 65660 21734 65686 21786
rect 65686 21734 65716 21786
rect 65740 21734 65750 21786
rect 65750 21734 65796 21786
rect 65820 21734 65866 21786
rect 65866 21734 65876 21786
rect 65900 21734 65930 21786
rect 65930 21734 65956 21786
rect 65660 21732 65716 21734
rect 65740 21732 65796 21734
rect 65820 21732 65876 21734
rect 65900 21732 65956 21734
rect 65522 21528 65578 21584
rect 66534 29588 66536 29608
rect 66536 29588 66588 29608
rect 66588 29588 66590 29608
rect 66534 29552 66590 29588
rect 66166 21528 66222 21584
rect 65660 20698 65716 20700
rect 65740 20698 65796 20700
rect 65820 20698 65876 20700
rect 65900 20698 65956 20700
rect 65660 20646 65686 20698
rect 65686 20646 65716 20698
rect 65740 20646 65750 20698
rect 65750 20646 65796 20698
rect 65820 20646 65866 20698
rect 65866 20646 65876 20698
rect 65900 20646 65930 20698
rect 65930 20646 65956 20698
rect 65660 20644 65716 20646
rect 65740 20644 65796 20646
rect 65820 20644 65876 20646
rect 65900 20644 65956 20646
rect 65982 20440 66038 20496
rect 65660 19610 65716 19612
rect 65740 19610 65796 19612
rect 65820 19610 65876 19612
rect 65900 19610 65956 19612
rect 65660 19558 65686 19610
rect 65686 19558 65716 19610
rect 65740 19558 65750 19610
rect 65750 19558 65796 19610
rect 65820 19558 65866 19610
rect 65866 19558 65876 19610
rect 65900 19558 65930 19610
rect 65930 19558 65956 19610
rect 65660 19556 65716 19558
rect 65740 19556 65796 19558
rect 65820 19556 65876 19558
rect 65900 19556 65956 19558
rect 65660 18522 65716 18524
rect 65740 18522 65796 18524
rect 65820 18522 65876 18524
rect 65900 18522 65956 18524
rect 65660 18470 65686 18522
rect 65686 18470 65716 18522
rect 65740 18470 65750 18522
rect 65750 18470 65796 18522
rect 65820 18470 65866 18522
rect 65866 18470 65876 18522
rect 65900 18470 65930 18522
rect 65930 18470 65956 18522
rect 65660 18468 65716 18470
rect 65740 18468 65796 18470
rect 65820 18468 65876 18470
rect 65900 18468 65956 18470
rect 65062 11056 65118 11112
rect 65062 8880 65118 8936
rect 65660 17434 65716 17436
rect 65740 17434 65796 17436
rect 65820 17434 65876 17436
rect 65900 17434 65956 17436
rect 65660 17382 65686 17434
rect 65686 17382 65716 17434
rect 65740 17382 65750 17434
rect 65750 17382 65796 17434
rect 65820 17382 65866 17434
rect 65866 17382 65876 17434
rect 65900 17382 65930 17434
rect 65930 17382 65956 17434
rect 65660 17380 65716 17382
rect 65740 17380 65796 17382
rect 65820 17380 65876 17382
rect 65900 17380 65956 17382
rect 65660 16346 65716 16348
rect 65740 16346 65796 16348
rect 65820 16346 65876 16348
rect 65900 16346 65956 16348
rect 65660 16294 65686 16346
rect 65686 16294 65716 16346
rect 65740 16294 65750 16346
rect 65750 16294 65796 16346
rect 65820 16294 65866 16346
rect 65866 16294 65876 16346
rect 65900 16294 65930 16346
rect 65930 16294 65956 16346
rect 65660 16292 65716 16294
rect 65740 16292 65796 16294
rect 65820 16292 65876 16294
rect 65900 16292 65956 16294
rect 65614 15580 65616 15600
rect 65616 15580 65668 15600
rect 65668 15580 65670 15600
rect 65614 15544 65670 15580
rect 65660 15258 65716 15260
rect 65740 15258 65796 15260
rect 65820 15258 65876 15260
rect 65900 15258 65956 15260
rect 65660 15206 65686 15258
rect 65686 15206 65716 15258
rect 65740 15206 65750 15258
rect 65750 15206 65796 15258
rect 65820 15206 65866 15258
rect 65866 15206 65876 15258
rect 65900 15206 65930 15258
rect 65930 15206 65956 15258
rect 65660 15204 65716 15206
rect 65740 15204 65796 15206
rect 65820 15204 65876 15206
rect 65900 15204 65956 15206
rect 65660 14170 65716 14172
rect 65740 14170 65796 14172
rect 65820 14170 65876 14172
rect 65900 14170 65956 14172
rect 65660 14118 65686 14170
rect 65686 14118 65716 14170
rect 65740 14118 65750 14170
rect 65750 14118 65796 14170
rect 65820 14118 65866 14170
rect 65866 14118 65876 14170
rect 65900 14118 65930 14170
rect 65930 14118 65956 14170
rect 65660 14116 65716 14118
rect 65740 14116 65796 14118
rect 65820 14116 65876 14118
rect 65900 14116 65956 14118
rect 65660 13082 65716 13084
rect 65740 13082 65796 13084
rect 65820 13082 65876 13084
rect 65900 13082 65956 13084
rect 65660 13030 65686 13082
rect 65686 13030 65716 13082
rect 65740 13030 65750 13082
rect 65750 13030 65796 13082
rect 65820 13030 65866 13082
rect 65866 13030 65876 13082
rect 65900 13030 65930 13082
rect 65930 13030 65956 13082
rect 65660 13028 65716 13030
rect 65740 13028 65796 13030
rect 65820 13028 65876 13030
rect 65900 13028 65956 13030
rect 66258 18264 66314 18320
rect 65660 11994 65716 11996
rect 65740 11994 65796 11996
rect 65820 11994 65876 11996
rect 65900 11994 65956 11996
rect 65660 11942 65686 11994
rect 65686 11942 65716 11994
rect 65740 11942 65750 11994
rect 65750 11942 65796 11994
rect 65820 11942 65866 11994
rect 65866 11942 65876 11994
rect 65900 11942 65930 11994
rect 65930 11942 65956 11994
rect 65660 11940 65716 11942
rect 65740 11940 65796 11942
rect 65820 11940 65876 11942
rect 65900 11940 65956 11942
rect 65660 10906 65716 10908
rect 65740 10906 65796 10908
rect 65820 10906 65876 10908
rect 65900 10906 65956 10908
rect 65660 10854 65686 10906
rect 65686 10854 65716 10906
rect 65740 10854 65750 10906
rect 65750 10854 65796 10906
rect 65820 10854 65866 10906
rect 65866 10854 65876 10906
rect 65900 10854 65930 10906
rect 65930 10854 65956 10906
rect 65660 10852 65716 10854
rect 65740 10852 65796 10854
rect 65820 10852 65876 10854
rect 65900 10852 65956 10854
rect 65660 9818 65716 9820
rect 65740 9818 65796 9820
rect 65820 9818 65876 9820
rect 65900 9818 65956 9820
rect 65660 9766 65686 9818
rect 65686 9766 65716 9818
rect 65740 9766 65750 9818
rect 65750 9766 65796 9818
rect 65820 9766 65866 9818
rect 65866 9766 65876 9818
rect 65900 9766 65930 9818
rect 65930 9766 65956 9818
rect 65660 9764 65716 9766
rect 65740 9764 65796 9766
rect 65820 9764 65876 9766
rect 65900 9764 65956 9766
rect 65522 9444 65578 9480
rect 65522 9424 65524 9444
rect 65524 9424 65576 9444
rect 65576 9424 65578 9444
rect 65660 8730 65716 8732
rect 65740 8730 65796 8732
rect 65820 8730 65876 8732
rect 65900 8730 65956 8732
rect 65660 8678 65686 8730
rect 65686 8678 65716 8730
rect 65740 8678 65750 8730
rect 65750 8678 65796 8730
rect 65820 8678 65866 8730
rect 65866 8678 65876 8730
rect 65900 8678 65930 8730
rect 65930 8678 65956 8730
rect 65660 8676 65716 8678
rect 65740 8676 65796 8678
rect 65820 8676 65876 8678
rect 65900 8676 65956 8678
rect 65154 7928 65210 7984
rect 65154 5108 65156 5128
rect 65156 5108 65208 5128
rect 65208 5108 65210 5128
rect 65154 5072 65210 5108
rect 64970 4392 65026 4448
rect 65660 7642 65716 7644
rect 65740 7642 65796 7644
rect 65820 7642 65876 7644
rect 65900 7642 65956 7644
rect 65660 7590 65686 7642
rect 65686 7590 65716 7642
rect 65740 7590 65750 7642
rect 65750 7590 65796 7642
rect 65820 7590 65866 7642
rect 65866 7590 65876 7642
rect 65900 7590 65930 7642
rect 65930 7590 65956 7642
rect 65660 7588 65716 7590
rect 65740 7588 65796 7590
rect 65820 7588 65876 7590
rect 65900 7588 65956 7590
rect 65660 6554 65716 6556
rect 65740 6554 65796 6556
rect 65820 6554 65876 6556
rect 65900 6554 65956 6556
rect 65660 6502 65686 6554
rect 65686 6502 65716 6554
rect 65740 6502 65750 6554
rect 65750 6502 65796 6554
rect 65820 6502 65866 6554
rect 65866 6502 65876 6554
rect 65900 6502 65930 6554
rect 65930 6502 65956 6554
rect 65660 6500 65716 6502
rect 65740 6500 65796 6502
rect 65820 6500 65876 6502
rect 65900 6500 65956 6502
rect 65660 5466 65716 5468
rect 65740 5466 65796 5468
rect 65820 5466 65876 5468
rect 65900 5466 65956 5468
rect 65660 5414 65686 5466
rect 65686 5414 65716 5466
rect 65740 5414 65750 5466
rect 65750 5414 65796 5466
rect 65820 5414 65866 5466
rect 65866 5414 65876 5466
rect 65900 5414 65930 5466
rect 65930 5414 65956 5466
rect 65660 5412 65716 5414
rect 65740 5412 65796 5414
rect 65820 5412 65876 5414
rect 65900 5412 65956 5414
rect 65660 4378 65716 4380
rect 65740 4378 65796 4380
rect 65820 4378 65876 4380
rect 65900 4378 65956 4380
rect 65660 4326 65686 4378
rect 65686 4326 65716 4378
rect 65740 4326 65750 4378
rect 65750 4326 65796 4378
rect 65820 4326 65866 4378
rect 65866 4326 65876 4378
rect 65900 4326 65930 4378
rect 65930 4326 65956 4378
rect 65660 4324 65716 4326
rect 65740 4324 65796 4326
rect 65820 4324 65876 4326
rect 65900 4324 65956 4326
rect 65660 3290 65716 3292
rect 65740 3290 65796 3292
rect 65820 3290 65876 3292
rect 65900 3290 65956 3292
rect 65660 3238 65686 3290
rect 65686 3238 65716 3290
rect 65740 3238 65750 3290
rect 65750 3238 65796 3290
rect 65820 3238 65866 3290
rect 65866 3238 65876 3290
rect 65900 3238 65930 3290
rect 65930 3238 65956 3290
rect 65660 3236 65716 3238
rect 65740 3236 65796 3238
rect 65820 3236 65876 3238
rect 65900 3236 65956 3238
rect 65660 2202 65716 2204
rect 65740 2202 65796 2204
rect 65820 2202 65876 2204
rect 65900 2202 65956 2204
rect 65660 2150 65686 2202
rect 65686 2150 65716 2202
rect 65740 2150 65750 2202
rect 65750 2150 65796 2202
rect 65820 2150 65866 2202
rect 65866 2150 65876 2202
rect 65900 2150 65930 2202
rect 65930 2150 65956 2202
rect 65660 2148 65716 2150
rect 65740 2148 65796 2150
rect 65820 2148 65876 2150
rect 65900 2148 65956 2150
rect 67086 33904 67142 33960
rect 67454 29588 67456 29608
rect 67456 29588 67508 29608
rect 67508 29588 67510 29608
rect 67454 29552 67510 29588
rect 67914 29028 67970 29064
rect 67914 29008 67916 29028
rect 67916 29008 67968 29028
rect 67968 29008 67970 29028
rect 67362 20848 67418 20904
rect 68926 37304 68982 37360
rect 68282 29144 68338 29200
rect 68282 10512 68338 10568
rect 68282 9716 68338 9752
rect 68282 9696 68284 9716
rect 68284 9696 68336 9716
rect 68336 9696 68338 9716
rect 68650 10104 68706 10160
rect 69110 10512 69166 10568
rect 69570 37032 69626 37088
rect 69386 29028 69442 29064
rect 69386 29008 69388 29028
rect 69388 29008 69440 29028
rect 69440 29008 69442 29028
rect 69294 25744 69350 25800
rect 69294 18844 69296 18864
rect 69296 18844 69348 18864
rect 69348 18844 69350 18864
rect 69294 18808 69350 18844
rect 70214 36236 70270 36272
rect 70214 36216 70216 36236
rect 70216 36216 70268 36236
rect 70268 36216 70270 36236
rect 69662 14764 69664 14784
rect 69664 14764 69716 14784
rect 69716 14764 69718 14784
rect 69662 14728 69718 14764
rect 70214 18808 70270 18864
rect 70030 15136 70086 15192
rect 69938 9696 69994 9752
rect 70306 15136 70362 15192
rect 70674 37032 70730 37088
rect 70490 36760 70546 36816
rect 70490 36372 70546 36408
rect 70490 36352 70492 36372
rect 70492 36352 70544 36372
rect 70544 36352 70546 36372
rect 73434 36760 73490 36816
rect 72054 36352 72110 36408
rect 70766 18828 70822 18864
rect 70766 18808 70768 18828
rect 70768 18808 70820 18828
rect 70820 18808 70822 18828
rect 71134 18828 71190 18864
rect 71134 18808 71136 18828
rect 71136 18808 71188 18828
rect 71188 18808 71190 18828
rect 71042 14728 71098 14784
rect 70214 12588 70216 12608
rect 70216 12588 70268 12608
rect 70268 12588 70270 12608
rect 70214 12552 70270 12588
rect 67454 448 67510 504
rect 71870 23724 71926 23760
rect 71870 23704 71872 23724
rect 71872 23704 71924 23724
rect 71924 23704 71926 23724
rect 71962 17720 72018 17776
rect 71686 10104 71742 10160
rect 72514 26324 72516 26344
rect 72516 26324 72568 26344
rect 72568 26324 72570 26344
rect 72514 26288 72570 26324
rect 74078 29144 74134 29200
rect 72422 18672 72478 18728
rect 71962 2488 72018 2544
rect 72330 2488 72386 2544
rect 74354 26324 74356 26344
rect 74356 26324 74408 26344
rect 74408 26324 74410 26344
rect 74354 26288 74410 26324
rect 74170 25336 74226 25392
rect 74170 7384 74226 7440
rect 74722 24132 74778 24168
rect 74722 24112 74724 24132
rect 74724 24112 74776 24132
rect 74776 24112 74778 24132
rect 74538 6704 74594 6760
rect 75274 36216 75330 36272
rect 75090 24384 75146 24440
rect 76102 36896 76158 36952
rect 76838 37340 76840 37360
rect 76840 37340 76892 37360
rect 76892 37340 76894 37360
rect 76838 37304 76894 37340
rect 75734 24268 75790 24304
rect 75734 24248 75736 24268
rect 75736 24248 75788 24268
rect 75788 24248 75790 24268
rect 75642 6160 75698 6216
rect 76378 24384 76434 24440
rect 76286 24248 76342 24304
rect 76286 23704 76342 23760
rect 75918 12588 75920 12608
rect 75920 12588 75972 12608
rect 75972 12588 75974 12608
rect 75918 12552 75974 12588
rect 77022 26696 77078 26752
rect 77390 26868 77392 26888
rect 77392 26868 77444 26888
rect 77444 26868 77446 26888
rect 77390 26832 77446 26868
rect 81020 37562 81076 37564
rect 81100 37562 81156 37564
rect 81180 37562 81236 37564
rect 81260 37562 81316 37564
rect 81020 37510 81046 37562
rect 81046 37510 81076 37562
rect 81100 37510 81110 37562
rect 81110 37510 81156 37562
rect 81180 37510 81226 37562
rect 81226 37510 81236 37562
rect 81260 37510 81290 37562
rect 81290 37510 81316 37562
rect 81020 37508 81076 37510
rect 81100 37508 81156 37510
rect 81180 37508 81236 37510
rect 81260 37508 81316 37510
rect 75550 176 75606 232
rect 78126 26732 78128 26752
rect 78128 26732 78180 26752
rect 78180 26732 78182 26752
rect 78126 26696 78182 26732
rect 78494 26852 78550 26888
rect 78494 26832 78496 26852
rect 78496 26832 78548 26852
rect 78548 26832 78550 26852
rect 78494 24112 78550 24168
rect 77758 856 77814 912
rect 77390 312 77446 368
rect 81020 36474 81076 36476
rect 81100 36474 81156 36476
rect 81180 36474 81236 36476
rect 81260 36474 81316 36476
rect 81020 36422 81046 36474
rect 81046 36422 81076 36474
rect 81100 36422 81110 36474
rect 81110 36422 81156 36474
rect 81180 36422 81226 36474
rect 81226 36422 81236 36474
rect 81260 36422 81290 36474
rect 81290 36422 81316 36474
rect 81020 36420 81076 36422
rect 81100 36420 81156 36422
rect 81180 36420 81236 36422
rect 81260 36420 81316 36422
rect 81020 35386 81076 35388
rect 81100 35386 81156 35388
rect 81180 35386 81236 35388
rect 81260 35386 81316 35388
rect 81020 35334 81046 35386
rect 81046 35334 81076 35386
rect 81100 35334 81110 35386
rect 81110 35334 81156 35386
rect 81180 35334 81226 35386
rect 81226 35334 81236 35386
rect 81260 35334 81290 35386
rect 81290 35334 81316 35386
rect 81020 35332 81076 35334
rect 81100 35332 81156 35334
rect 81180 35332 81236 35334
rect 81260 35332 81316 35334
rect 81020 34298 81076 34300
rect 81100 34298 81156 34300
rect 81180 34298 81236 34300
rect 81260 34298 81316 34300
rect 81020 34246 81046 34298
rect 81046 34246 81076 34298
rect 81100 34246 81110 34298
rect 81110 34246 81156 34298
rect 81180 34246 81226 34298
rect 81226 34246 81236 34298
rect 81260 34246 81290 34298
rect 81290 34246 81316 34298
rect 81020 34244 81076 34246
rect 81100 34244 81156 34246
rect 81180 34244 81236 34246
rect 81260 34244 81316 34246
rect 81020 33210 81076 33212
rect 81100 33210 81156 33212
rect 81180 33210 81236 33212
rect 81260 33210 81316 33212
rect 81020 33158 81046 33210
rect 81046 33158 81076 33210
rect 81100 33158 81110 33210
rect 81110 33158 81156 33210
rect 81180 33158 81226 33210
rect 81226 33158 81236 33210
rect 81260 33158 81290 33210
rect 81290 33158 81316 33210
rect 81020 33156 81076 33158
rect 81100 33156 81156 33158
rect 81180 33156 81236 33158
rect 81260 33156 81316 33158
rect 79506 28464 79562 28520
rect 79046 20324 79102 20360
rect 79046 20304 79048 20324
rect 79048 20304 79100 20324
rect 79100 20304 79102 20324
rect 81020 32122 81076 32124
rect 81100 32122 81156 32124
rect 81180 32122 81236 32124
rect 81260 32122 81316 32124
rect 81020 32070 81046 32122
rect 81046 32070 81076 32122
rect 81100 32070 81110 32122
rect 81110 32070 81156 32122
rect 81180 32070 81226 32122
rect 81226 32070 81236 32122
rect 81260 32070 81290 32122
rect 81290 32070 81316 32122
rect 81020 32068 81076 32070
rect 81100 32068 81156 32070
rect 81180 32068 81236 32070
rect 81260 32068 81316 32070
rect 81020 31034 81076 31036
rect 81100 31034 81156 31036
rect 81180 31034 81236 31036
rect 81260 31034 81316 31036
rect 81020 30982 81046 31034
rect 81046 30982 81076 31034
rect 81100 30982 81110 31034
rect 81110 30982 81156 31034
rect 81180 30982 81226 31034
rect 81226 30982 81236 31034
rect 81260 30982 81290 31034
rect 81290 30982 81316 31034
rect 81020 30980 81076 30982
rect 81100 30980 81156 30982
rect 81180 30980 81236 30982
rect 81260 30980 81316 30982
rect 80058 30640 80114 30696
rect 81020 29946 81076 29948
rect 81100 29946 81156 29948
rect 81180 29946 81236 29948
rect 81260 29946 81316 29948
rect 81020 29894 81046 29946
rect 81046 29894 81076 29946
rect 81100 29894 81110 29946
rect 81110 29894 81156 29946
rect 81180 29894 81226 29946
rect 81226 29894 81236 29946
rect 81260 29894 81290 29946
rect 81290 29894 81316 29946
rect 81020 29892 81076 29894
rect 81100 29892 81156 29894
rect 81180 29892 81236 29894
rect 81260 29892 81316 29894
rect 81020 28858 81076 28860
rect 81100 28858 81156 28860
rect 81180 28858 81236 28860
rect 81260 28858 81316 28860
rect 81020 28806 81046 28858
rect 81046 28806 81076 28858
rect 81100 28806 81110 28858
rect 81110 28806 81156 28858
rect 81180 28806 81226 28858
rect 81226 28806 81236 28858
rect 81260 28806 81290 28858
rect 81290 28806 81316 28858
rect 81020 28804 81076 28806
rect 81100 28804 81156 28806
rect 81180 28804 81236 28806
rect 81260 28804 81316 28806
rect 81020 27770 81076 27772
rect 81100 27770 81156 27772
rect 81180 27770 81236 27772
rect 81260 27770 81316 27772
rect 81020 27718 81046 27770
rect 81046 27718 81076 27770
rect 81100 27718 81110 27770
rect 81110 27718 81156 27770
rect 81180 27718 81226 27770
rect 81226 27718 81236 27770
rect 81260 27718 81290 27770
rect 81290 27718 81316 27770
rect 81020 27716 81076 27718
rect 81100 27716 81156 27718
rect 81180 27716 81236 27718
rect 81260 27716 81316 27718
rect 81020 26682 81076 26684
rect 81100 26682 81156 26684
rect 81180 26682 81236 26684
rect 81260 26682 81316 26684
rect 81020 26630 81046 26682
rect 81046 26630 81076 26682
rect 81100 26630 81110 26682
rect 81110 26630 81156 26682
rect 81180 26630 81226 26682
rect 81226 26630 81236 26682
rect 81260 26630 81290 26682
rect 81290 26630 81316 26682
rect 81020 26628 81076 26630
rect 81100 26628 81156 26630
rect 81180 26628 81236 26630
rect 81260 26628 81316 26630
rect 81020 25594 81076 25596
rect 81100 25594 81156 25596
rect 81180 25594 81236 25596
rect 81260 25594 81316 25596
rect 81020 25542 81046 25594
rect 81046 25542 81076 25594
rect 81100 25542 81110 25594
rect 81110 25542 81156 25594
rect 81180 25542 81226 25594
rect 81226 25542 81236 25594
rect 81260 25542 81290 25594
rect 81290 25542 81316 25594
rect 81020 25540 81076 25542
rect 81100 25540 81156 25542
rect 81180 25540 81236 25542
rect 81260 25540 81316 25542
rect 81020 24506 81076 24508
rect 81100 24506 81156 24508
rect 81180 24506 81236 24508
rect 81260 24506 81316 24508
rect 81020 24454 81046 24506
rect 81046 24454 81076 24506
rect 81100 24454 81110 24506
rect 81110 24454 81156 24506
rect 81180 24454 81226 24506
rect 81226 24454 81236 24506
rect 81260 24454 81290 24506
rect 81290 24454 81316 24506
rect 81020 24452 81076 24454
rect 81100 24452 81156 24454
rect 81180 24452 81236 24454
rect 81260 24452 81316 24454
rect 81020 23418 81076 23420
rect 81100 23418 81156 23420
rect 81180 23418 81236 23420
rect 81260 23418 81316 23420
rect 81020 23366 81046 23418
rect 81046 23366 81076 23418
rect 81100 23366 81110 23418
rect 81110 23366 81156 23418
rect 81180 23366 81226 23418
rect 81226 23366 81236 23418
rect 81260 23366 81290 23418
rect 81290 23366 81316 23418
rect 81020 23364 81076 23366
rect 81100 23364 81156 23366
rect 81180 23364 81236 23366
rect 81260 23364 81316 23366
rect 81020 22330 81076 22332
rect 81100 22330 81156 22332
rect 81180 22330 81236 22332
rect 81260 22330 81316 22332
rect 81020 22278 81046 22330
rect 81046 22278 81076 22330
rect 81100 22278 81110 22330
rect 81110 22278 81156 22330
rect 81180 22278 81226 22330
rect 81226 22278 81236 22330
rect 81260 22278 81290 22330
rect 81290 22278 81316 22330
rect 81020 22276 81076 22278
rect 81100 22276 81156 22278
rect 81180 22276 81236 22278
rect 81260 22276 81316 22278
rect 81020 21242 81076 21244
rect 81100 21242 81156 21244
rect 81180 21242 81236 21244
rect 81260 21242 81316 21244
rect 81020 21190 81046 21242
rect 81046 21190 81076 21242
rect 81100 21190 81110 21242
rect 81110 21190 81156 21242
rect 81180 21190 81226 21242
rect 81226 21190 81236 21242
rect 81260 21190 81290 21242
rect 81290 21190 81316 21242
rect 81020 21188 81076 21190
rect 81100 21188 81156 21190
rect 81180 21188 81236 21190
rect 81260 21188 81316 21190
rect 80978 20460 81034 20496
rect 80978 20440 80980 20460
rect 80980 20440 81032 20460
rect 81032 20440 81034 20460
rect 81020 20154 81076 20156
rect 81100 20154 81156 20156
rect 81180 20154 81236 20156
rect 81260 20154 81316 20156
rect 81020 20102 81046 20154
rect 81046 20102 81076 20154
rect 81100 20102 81110 20154
rect 81110 20102 81156 20154
rect 81180 20102 81226 20154
rect 81226 20102 81236 20154
rect 81260 20102 81290 20154
rect 81290 20102 81316 20154
rect 81020 20100 81076 20102
rect 81100 20100 81156 20102
rect 81180 20100 81236 20102
rect 81260 20100 81316 20102
rect 81020 19066 81076 19068
rect 81100 19066 81156 19068
rect 81180 19066 81236 19068
rect 81260 19066 81316 19068
rect 81020 19014 81046 19066
rect 81046 19014 81076 19066
rect 81100 19014 81110 19066
rect 81110 19014 81156 19066
rect 81180 19014 81226 19066
rect 81226 19014 81236 19066
rect 81260 19014 81290 19066
rect 81290 19014 81316 19066
rect 81020 19012 81076 19014
rect 81100 19012 81156 19014
rect 81180 19012 81236 19014
rect 81260 19012 81316 19014
rect 81020 17978 81076 17980
rect 81100 17978 81156 17980
rect 81180 17978 81236 17980
rect 81260 17978 81316 17980
rect 81020 17926 81046 17978
rect 81046 17926 81076 17978
rect 81100 17926 81110 17978
rect 81110 17926 81156 17978
rect 81180 17926 81226 17978
rect 81226 17926 81236 17978
rect 81260 17926 81290 17978
rect 81290 17926 81316 17978
rect 81020 17924 81076 17926
rect 81100 17924 81156 17926
rect 81180 17924 81236 17926
rect 81260 17924 81316 17926
rect 81020 16890 81076 16892
rect 81100 16890 81156 16892
rect 81180 16890 81236 16892
rect 81260 16890 81316 16892
rect 81020 16838 81046 16890
rect 81046 16838 81076 16890
rect 81100 16838 81110 16890
rect 81110 16838 81156 16890
rect 81180 16838 81226 16890
rect 81226 16838 81236 16890
rect 81260 16838 81290 16890
rect 81290 16838 81316 16890
rect 81020 16836 81076 16838
rect 81100 16836 81156 16838
rect 81180 16836 81236 16838
rect 81260 16836 81316 16838
rect 81020 15802 81076 15804
rect 81100 15802 81156 15804
rect 81180 15802 81236 15804
rect 81260 15802 81316 15804
rect 81020 15750 81046 15802
rect 81046 15750 81076 15802
rect 81100 15750 81110 15802
rect 81110 15750 81156 15802
rect 81180 15750 81226 15802
rect 81226 15750 81236 15802
rect 81260 15750 81290 15802
rect 81290 15750 81316 15802
rect 81020 15748 81076 15750
rect 81100 15748 81156 15750
rect 81180 15748 81236 15750
rect 81260 15748 81316 15750
rect 81020 14714 81076 14716
rect 81100 14714 81156 14716
rect 81180 14714 81236 14716
rect 81260 14714 81316 14716
rect 81020 14662 81046 14714
rect 81046 14662 81076 14714
rect 81100 14662 81110 14714
rect 81110 14662 81156 14714
rect 81180 14662 81226 14714
rect 81226 14662 81236 14714
rect 81260 14662 81290 14714
rect 81290 14662 81316 14714
rect 81020 14660 81076 14662
rect 81100 14660 81156 14662
rect 81180 14660 81236 14662
rect 81260 14660 81316 14662
rect 81020 13626 81076 13628
rect 81100 13626 81156 13628
rect 81180 13626 81236 13628
rect 81260 13626 81316 13628
rect 81020 13574 81046 13626
rect 81046 13574 81076 13626
rect 81100 13574 81110 13626
rect 81110 13574 81156 13626
rect 81180 13574 81226 13626
rect 81226 13574 81236 13626
rect 81260 13574 81290 13626
rect 81290 13574 81316 13626
rect 81020 13572 81076 13574
rect 81100 13572 81156 13574
rect 81180 13572 81236 13574
rect 81260 13572 81316 13574
rect 81020 12538 81076 12540
rect 81100 12538 81156 12540
rect 81180 12538 81236 12540
rect 81260 12538 81316 12540
rect 81020 12486 81046 12538
rect 81046 12486 81076 12538
rect 81100 12486 81110 12538
rect 81110 12486 81156 12538
rect 81180 12486 81226 12538
rect 81226 12486 81236 12538
rect 81260 12486 81290 12538
rect 81290 12486 81316 12538
rect 81020 12484 81076 12486
rect 81100 12484 81156 12486
rect 81180 12484 81236 12486
rect 81260 12484 81316 12486
rect 81020 11450 81076 11452
rect 81100 11450 81156 11452
rect 81180 11450 81236 11452
rect 81260 11450 81316 11452
rect 81020 11398 81046 11450
rect 81046 11398 81076 11450
rect 81100 11398 81110 11450
rect 81110 11398 81156 11450
rect 81180 11398 81226 11450
rect 81226 11398 81236 11450
rect 81260 11398 81290 11450
rect 81290 11398 81316 11450
rect 81020 11396 81076 11398
rect 81100 11396 81156 11398
rect 81180 11396 81236 11398
rect 81260 11396 81316 11398
rect 81020 10362 81076 10364
rect 81100 10362 81156 10364
rect 81180 10362 81236 10364
rect 81260 10362 81316 10364
rect 81020 10310 81046 10362
rect 81046 10310 81076 10362
rect 81100 10310 81110 10362
rect 81110 10310 81156 10362
rect 81180 10310 81226 10362
rect 81226 10310 81236 10362
rect 81260 10310 81290 10362
rect 81290 10310 81316 10362
rect 81020 10308 81076 10310
rect 81100 10308 81156 10310
rect 81180 10308 81236 10310
rect 81260 10308 81316 10310
rect 81020 9274 81076 9276
rect 81100 9274 81156 9276
rect 81180 9274 81236 9276
rect 81260 9274 81316 9276
rect 81020 9222 81046 9274
rect 81046 9222 81076 9274
rect 81100 9222 81110 9274
rect 81110 9222 81156 9274
rect 81180 9222 81226 9274
rect 81226 9222 81236 9274
rect 81260 9222 81290 9274
rect 81290 9222 81316 9274
rect 81020 9220 81076 9222
rect 81100 9220 81156 9222
rect 81180 9220 81236 9222
rect 81260 9220 81316 9222
rect 81020 8186 81076 8188
rect 81100 8186 81156 8188
rect 81180 8186 81236 8188
rect 81260 8186 81316 8188
rect 81020 8134 81046 8186
rect 81046 8134 81076 8186
rect 81100 8134 81110 8186
rect 81110 8134 81156 8186
rect 81180 8134 81226 8186
rect 81226 8134 81236 8186
rect 81260 8134 81290 8186
rect 81290 8134 81316 8186
rect 81020 8132 81076 8134
rect 81100 8132 81156 8134
rect 81180 8132 81236 8134
rect 81260 8132 81316 8134
rect 81020 7098 81076 7100
rect 81100 7098 81156 7100
rect 81180 7098 81236 7100
rect 81260 7098 81316 7100
rect 81020 7046 81046 7098
rect 81046 7046 81076 7098
rect 81100 7046 81110 7098
rect 81110 7046 81156 7098
rect 81180 7046 81226 7098
rect 81226 7046 81236 7098
rect 81260 7046 81290 7098
rect 81290 7046 81316 7098
rect 81020 7044 81076 7046
rect 81100 7044 81156 7046
rect 81180 7044 81236 7046
rect 81260 7044 81316 7046
rect 83738 34584 83794 34640
rect 82266 20460 82322 20496
rect 82266 20440 82268 20460
rect 82268 20440 82320 20460
rect 82320 20440 82322 20460
rect 82174 20340 82176 20360
rect 82176 20340 82228 20360
rect 82228 20340 82230 20360
rect 82174 20304 82230 20340
rect 81020 6010 81076 6012
rect 81100 6010 81156 6012
rect 81180 6010 81236 6012
rect 81260 6010 81316 6012
rect 81020 5958 81046 6010
rect 81046 5958 81076 6010
rect 81100 5958 81110 6010
rect 81110 5958 81156 6010
rect 81180 5958 81226 6010
rect 81226 5958 81236 6010
rect 81260 5958 81290 6010
rect 81290 5958 81316 6010
rect 81020 5956 81076 5958
rect 81100 5956 81156 5958
rect 81180 5956 81236 5958
rect 81260 5956 81316 5958
rect 81020 4922 81076 4924
rect 81100 4922 81156 4924
rect 81180 4922 81236 4924
rect 81260 4922 81316 4924
rect 81020 4870 81046 4922
rect 81046 4870 81076 4922
rect 81100 4870 81110 4922
rect 81110 4870 81156 4922
rect 81180 4870 81226 4922
rect 81226 4870 81236 4922
rect 81260 4870 81290 4922
rect 81290 4870 81316 4922
rect 81020 4868 81076 4870
rect 81100 4868 81156 4870
rect 81180 4868 81236 4870
rect 81260 4868 81316 4870
rect 81020 3834 81076 3836
rect 81100 3834 81156 3836
rect 81180 3834 81236 3836
rect 81260 3834 81316 3836
rect 81020 3782 81046 3834
rect 81046 3782 81076 3834
rect 81100 3782 81110 3834
rect 81110 3782 81156 3834
rect 81180 3782 81226 3834
rect 81226 3782 81236 3834
rect 81260 3782 81290 3834
rect 81290 3782 81316 3834
rect 81020 3780 81076 3782
rect 81100 3780 81156 3782
rect 81180 3780 81236 3782
rect 81260 3780 81316 3782
rect 81020 2746 81076 2748
rect 81100 2746 81156 2748
rect 81180 2746 81236 2748
rect 81260 2746 81316 2748
rect 81020 2694 81046 2746
rect 81046 2694 81076 2746
rect 81100 2694 81110 2746
rect 81110 2694 81156 2746
rect 81180 2694 81226 2746
rect 81226 2694 81236 2746
rect 81260 2694 81290 2746
rect 81290 2694 81316 2746
rect 81020 2692 81076 2694
rect 81100 2692 81156 2694
rect 81180 2692 81236 2694
rect 81260 2692 81316 2694
rect 84658 36080 84714 36136
rect 85302 21972 85304 21992
rect 85304 21972 85356 21992
rect 85356 21972 85358 21992
rect 85302 21936 85358 21972
rect 85578 12860 85580 12880
rect 85580 12860 85632 12880
rect 85632 12860 85634 12880
rect 85578 12824 85634 12860
rect 85578 7248 85634 7304
rect 85118 992 85174 1048
rect 86130 26324 86132 26344
rect 86132 26324 86184 26344
rect 86184 26324 86186 26344
rect 86130 26288 86186 26324
rect 86038 12824 86094 12880
rect 88246 26324 88248 26344
rect 88248 26324 88300 26344
rect 88300 26324 88302 26344
rect 88246 26288 88302 26324
rect 90362 33496 90418 33552
rect 89902 33360 89958 33416
rect 82082 584 82138 640
rect 87970 1264 88026 1320
rect 88430 1128 88486 1184
rect 89258 11192 89314 11248
rect 90454 5208 90510 5264
rect 90822 5208 90878 5264
rect 91466 27920 91522 27976
rect 96380 37018 96436 37020
rect 96460 37018 96516 37020
rect 96540 37018 96596 37020
rect 96620 37018 96676 37020
rect 96380 36966 96406 37018
rect 96406 36966 96436 37018
rect 96460 36966 96470 37018
rect 96470 36966 96516 37018
rect 96540 36966 96586 37018
rect 96586 36966 96596 37018
rect 96620 36966 96650 37018
rect 96650 36966 96676 37018
rect 96380 36964 96436 36966
rect 96460 36964 96516 36966
rect 96540 36964 96596 36966
rect 96620 36964 96676 36966
rect 97630 36644 97686 36680
rect 97630 36624 97632 36644
rect 97632 36624 97684 36644
rect 97684 36624 97686 36644
rect 96380 35930 96436 35932
rect 96460 35930 96516 35932
rect 96540 35930 96596 35932
rect 96620 35930 96676 35932
rect 96380 35878 96406 35930
rect 96406 35878 96436 35930
rect 96460 35878 96470 35930
rect 96470 35878 96516 35930
rect 96540 35878 96586 35930
rect 96586 35878 96596 35930
rect 96620 35878 96650 35930
rect 96650 35878 96676 35930
rect 96380 35876 96436 35878
rect 96460 35876 96516 35878
rect 96540 35876 96596 35878
rect 96620 35876 96676 35878
rect 94134 16088 94190 16144
rect 96380 34842 96436 34844
rect 96460 34842 96516 34844
rect 96540 34842 96596 34844
rect 96620 34842 96676 34844
rect 96380 34790 96406 34842
rect 96406 34790 96436 34842
rect 96460 34790 96470 34842
rect 96470 34790 96516 34842
rect 96540 34790 96586 34842
rect 96586 34790 96596 34842
rect 96620 34790 96650 34842
rect 96650 34790 96676 34842
rect 96380 34788 96436 34790
rect 96460 34788 96516 34790
rect 96540 34788 96596 34790
rect 96620 34788 96676 34790
rect 96380 33754 96436 33756
rect 96460 33754 96516 33756
rect 96540 33754 96596 33756
rect 96620 33754 96676 33756
rect 96380 33702 96406 33754
rect 96406 33702 96436 33754
rect 96460 33702 96470 33754
rect 96470 33702 96516 33754
rect 96540 33702 96586 33754
rect 96586 33702 96596 33754
rect 96620 33702 96650 33754
rect 96650 33702 96676 33754
rect 96380 33700 96436 33702
rect 96460 33700 96516 33702
rect 96540 33700 96596 33702
rect 96620 33700 96676 33702
rect 96380 32666 96436 32668
rect 96460 32666 96516 32668
rect 96540 32666 96596 32668
rect 96620 32666 96676 32668
rect 96380 32614 96406 32666
rect 96406 32614 96436 32666
rect 96460 32614 96470 32666
rect 96470 32614 96516 32666
rect 96540 32614 96586 32666
rect 96586 32614 96596 32666
rect 96620 32614 96650 32666
rect 96650 32614 96676 32666
rect 96380 32612 96436 32614
rect 96460 32612 96516 32614
rect 96540 32612 96596 32614
rect 96620 32612 96676 32614
rect 96380 31578 96436 31580
rect 96460 31578 96516 31580
rect 96540 31578 96596 31580
rect 96620 31578 96676 31580
rect 96380 31526 96406 31578
rect 96406 31526 96436 31578
rect 96460 31526 96470 31578
rect 96470 31526 96516 31578
rect 96540 31526 96586 31578
rect 96586 31526 96596 31578
rect 96620 31526 96650 31578
rect 96650 31526 96676 31578
rect 96380 31524 96436 31526
rect 96460 31524 96516 31526
rect 96540 31524 96596 31526
rect 96620 31524 96676 31526
rect 96380 30490 96436 30492
rect 96460 30490 96516 30492
rect 96540 30490 96596 30492
rect 96620 30490 96676 30492
rect 96380 30438 96406 30490
rect 96406 30438 96436 30490
rect 96460 30438 96470 30490
rect 96470 30438 96516 30490
rect 96540 30438 96586 30490
rect 96586 30438 96596 30490
rect 96620 30438 96650 30490
rect 96650 30438 96676 30490
rect 96380 30436 96436 30438
rect 96460 30436 96516 30438
rect 96540 30436 96596 30438
rect 96620 30436 96676 30438
rect 96380 29402 96436 29404
rect 96460 29402 96516 29404
rect 96540 29402 96596 29404
rect 96620 29402 96676 29404
rect 96380 29350 96406 29402
rect 96406 29350 96436 29402
rect 96460 29350 96470 29402
rect 96470 29350 96516 29402
rect 96540 29350 96586 29402
rect 96586 29350 96596 29402
rect 96620 29350 96650 29402
rect 96650 29350 96676 29402
rect 96380 29348 96436 29350
rect 96460 29348 96516 29350
rect 96540 29348 96596 29350
rect 96620 29348 96676 29350
rect 96380 28314 96436 28316
rect 96460 28314 96516 28316
rect 96540 28314 96596 28316
rect 96620 28314 96676 28316
rect 96380 28262 96406 28314
rect 96406 28262 96436 28314
rect 96460 28262 96470 28314
rect 96470 28262 96516 28314
rect 96540 28262 96586 28314
rect 96586 28262 96596 28314
rect 96620 28262 96650 28314
rect 96650 28262 96676 28314
rect 96380 28260 96436 28262
rect 96460 28260 96516 28262
rect 96540 28260 96596 28262
rect 96620 28260 96676 28262
rect 96380 27226 96436 27228
rect 96460 27226 96516 27228
rect 96540 27226 96596 27228
rect 96620 27226 96676 27228
rect 96380 27174 96406 27226
rect 96406 27174 96436 27226
rect 96460 27174 96470 27226
rect 96470 27174 96516 27226
rect 96540 27174 96586 27226
rect 96586 27174 96596 27226
rect 96620 27174 96650 27226
rect 96650 27174 96676 27226
rect 96380 27172 96436 27174
rect 96460 27172 96516 27174
rect 96540 27172 96596 27174
rect 96620 27172 96676 27174
rect 96380 26138 96436 26140
rect 96460 26138 96516 26140
rect 96540 26138 96596 26140
rect 96620 26138 96676 26140
rect 96380 26086 96406 26138
rect 96406 26086 96436 26138
rect 96460 26086 96470 26138
rect 96470 26086 96516 26138
rect 96540 26086 96586 26138
rect 96586 26086 96596 26138
rect 96620 26086 96650 26138
rect 96650 26086 96676 26138
rect 96380 26084 96436 26086
rect 96460 26084 96516 26086
rect 96540 26084 96596 26086
rect 96620 26084 96676 26086
rect 96380 25050 96436 25052
rect 96460 25050 96516 25052
rect 96540 25050 96596 25052
rect 96620 25050 96676 25052
rect 96380 24998 96406 25050
rect 96406 24998 96436 25050
rect 96460 24998 96470 25050
rect 96470 24998 96516 25050
rect 96540 24998 96586 25050
rect 96586 24998 96596 25050
rect 96620 24998 96650 25050
rect 96650 24998 96676 25050
rect 96380 24996 96436 24998
rect 96460 24996 96516 24998
rect 96540 24996 96596 24998
rect 96620 24996 96676 24998
rect 96380 23962 96436 23964
rect 96460 23962 96516 23964
rect 96540 23962 96596 23964
rect 96620 23962 96676 23964
rect 96380 23910 96406 23962
rect 96406 23910 96436 23962
rect 96460 23910 96470 23962
rect 96470 23910 96516 23962
rect 96540 23910 96586 23962
rect 96586 23910 96596 23962
rect 96620 23910 96650 23962
rect 96650 23910 96676 23962
rect 96380 23908 96436 23910
rect 96460 23908 96516 23910
rect 96540 23908 96596 23910
rect 96620 23908 96676 23910
rect 96380 22874 96436 22876
rect 96460 22874 96516 22876
rect 96540 22874 96596 22876
rect 96620 22874 96676 22876
rect 96380 22822 96406 22874
rect 96406 22822 96436 22874
rect 96460 22822 96470 22874
rect 96470 22822 96516 22874
rect 96540 22822 96586 22874
rect 96586 22822 96596 22874
rect 96620 22822 96650 22874
rect 96650 22822 96676 22874
rect 96380 22820 96436 22822
rect 96460 22820 96516 22822
rect 96540 22820 96596 22822
rect 96620 22820 96676 22822
rect 96380 21786 96436 21788
rect 96460 21786 96516 21788
rect 96540 21786 96596 21788
rect 96620 21786 96676 21788
rect 96380 21734 96406 21786
rect 96406 21734 96436 21786
rect 96460 21734 96470 21786
rect 96470 21734 96516 21786
rect 96540 21734 96586 21786
rect 96586 21734 96596 21786
rect 96620 21734 96650 21786
rect 96650 21734 96676 21786
rect 96380 21732 96436 21734
rect 96460 21732 96516 21734
rect 96540 21732 96596 21734
rect 96620 21732 96676 21734
rect 96380 20698 96436 20700
rect 96460 20698 96516 20700
rect 96540 20698 96596 20700
rect 96620 20698 96676 20700
rect 96380 20646 96406 20698
rect 96406 20646 96436 20698
rect 96460 20646 96470 20698
rect 96470 20646 96516 20698
rect 96540 20646 96586 20698
rect 96586 20646 96596 20698
rect 96620 20646 96650 20698
rect 96650 20646 96676 20698
rect 96380 20644 96436 20646
rect 96460 20644 96516 20646
rect 96540 20644 96596 20646
rect 96620 20644 96676 20646
rect 96380 19610 96436 19612
rect 96460 19610 96516 19612
rect 96540 19610 96596 19612
rect 96620 19610 96676 19612
rect 96380 19558 96406 19610
rect 96406 19558 96436 19610
rect 96460 19558 96470 19610
rect 96470 19558 96516 19610
rect 96540 19558 96586 19610
rect 96586 19558 96596 19610
rect 96620 19558 96650 19610
rect 96650 19558 96676 19610
rect 96380 19556 96436 19558
rect 96460 19556 96516 19558
rect 96540 19556 96596 19558
rect 96620 19556 96676 19558
rect 96380 18522 96436 18524
rect 96460 18522 96516 18524
rect 96540 18522 96596 18524
rect 96620 18522 96676 18524
rect 96380 18470 96406 18522
rect 96406 18470 96436 18522
rect 96460 18470 96470 18522
rect 96470 18470 96516 18522
rect 96540 18470 96586 18522
rect 96586 18470 96596 18522
rect 96620 18470 96650 18522
rect 96650 18470 96676 18522
rect 96380 18468 96436 18470
rect 96460 18468 96516 18470
rect 96540 18468 96596 18470
rect 96620 18468 96676 18470
rect 96380 17434 96436 17436
rect 96460 17434 96516 17436
rect 96540 17434 96596 17436
rect 96620 17434 96676 17436
rect 96380 17382 96406 17434
rect 96406 17382 96436 17434
rect 96460 17382 96470 17434
rect 96470 17382 96516 17434
rect 96540 17382 96586 17434
rect 96586 17382 96596 17434
rect 96620 17382 96650 17434
rect 96650 17382 96676 17434
rect 96380 17380 96436 17382
rect 96460 17380 96516 17382
rect 96540 17380 96596 17382
rect 96620 17380 96676 17382
rect 97538 31184 97594 31240
rect 97630 20052 97686 20088
rect 97630 20032 97632 20052
rect 97632 20032 97684 20052
rect 97684 20032 97686 20052
rect 96986 18128 97042 18184
rect 96380 16346 96436 16348
rect 96460 16346 96516 16348
rect 96540 16346 96596 16348
rect 96620 16346 96676 16348
rect 96380 16294 96406 16346
rect 96406 16294 96436 16346
rect 96460 16294 96470 16346
rect 96470 16294 96516 16346
rect 96540 16294 96586 16346
rect 96586 16294 96596 16346
rect 96620 16294 96650 16346
rect 96650 16294 96676 16346
rect 96380 16292 96436 16294
rect 96460 16292 96516 16294
rect 96540 16292 96596 16294
rect 96620 16292 96676 16294
rect 96380 15258 96436 15260
rect 96460 15258 96516 15260
rect 96540 15258 96596 15260
rect 96620 15258 96676 15260
rect 96380 15206 96406 15258
rect 96406 15206 96436 15258
rect 96460 15206 96470 15258
rect 96470 15206 96516 15258
rect 96540 15206 96586 15258
rect 96586 15206 96596 15258
rect 96620 15206 96650 15258
rect 96650 15206 96676 15258
rect 96380 15204 96436 15206
rect 96460 15204 96516 15206
rect 96540 15204 96596 15206
rect 96620 15204 96676 15206
rect 96380 14170 96436 14172
rect 96460 14170 96516 14172
rect 96540 14170 96596 14172
rect 96620 14170 96676 14172
rect 96380 14118 96406 14170
rect 96406 14118 96436 14170
rect 96460 14118 96470 14170
rect 96470 14118 96516 14170
rect 96540 14118 96586 14170
rect 96586 14118 96596 14170
rect 96620 14118 96650 14170
rect 96650 14118 96676 14170
rect 96380 14116 96436 14118
rect 96460 14116 96516 14118
rect 96540 14116 96596 14118
rect 96620 14116 96676 14118
rect 96380 13082 96436 13084
rect 96460 13082 96516 13084
rect 96540 13082 96596 13084
rect 96620 13082 96676 13084
rect 96380 13030 96406 13082
rect 96406 13030 96436 13082
rect 96460 13030 96470 13082
rect 96470 13030 96516 13082
rect 96540 13030 96586 13082
rect 96586 13030 96596 13082
rect 96620 13030 96650 13082
rect 96650 13030 96676 13082
rect 96380 13028 96436 13030
rect 96460 13028 96516 13030
rect 96540 13028 96596 13030
rect 96620 13028 96676 13030
rect 96380 11994 96436 11996
rect 96460 11994 96516 11996
rect 96540 11994 96596 11996
rect 96620 11994 96676 11996
rect 96380 11942 96406 11994
rect 96406 11942 96436 11994
rect 96460 11942 96470 11994
rect 96470 11942 96516 11994
rect 96540 11942 96586 11994
rect 96586 11942 96596 11994
rect 96620 11942 96650 11994
rect 96650 11942 96676 11994
rect 96380 11940 96436 11942
rect 96460 11940 96516 11942
rect 96540 11940 96596 11942
rect 96620 11940 96676 11942
rect 96380 10906 96436 10908
rect 96460 10906 96516 10908
rect 96540 10906 96596 10908
rect 96620 10906 96676 10908
rect 96380 10854 96406 10906
rect 96406 10854 96436 10906
rect 96460 10854 96470 10906
rect 96470 10854 96516 10906
rect 96540 10854 96586 10906
rect 96586 10854 96596 10906
rect 96620 10854 96650 10906
rect 96650 10854 96676 10906
rect 96380 10852 96436 10854
rect 96460 10852 96516 10854
rect 96540 10852 96596 10854
rect 96620 10852 96676 10854
rect 95974 9016 96030 9072
rect 96380 9818 96436 9820
rect 96460 9818 96516 9820
rect 96540 9818 96596 9820
rect 96620 9818 96676 9820
rect 96380 9766 96406 9818
rect 96406 9766 96436 9818
rect 96460 9766 96470 9818
rect 96470 9766 96516 9818
rect 96540 9766 96586 9818
rect 96586 9766 96596 9818
rect 96620 9766 96650 9818
rect 96650 9766 96676 9818
rect 96380 9764 96436 9766
rect 96460 9764 96516 9766
rect 96540 9764 96596 9766
rect 96620 9764 96676 9766
rect 96380 8730 96436 8732
rect 96460 8730 96516 8732
rect 96540 8730 96596 8732
rect 96620 8730 96676 8732
rect 96380 8678 96406 8730
rect 96406 8678 96436 8730
rect 96460 8678 96470 8730
rect 96470 8678 96516 8730
rect 96540 8678 96586 8730
rect 96586 8678 96596 8730
rect 96620 8678 96650 8730
rect 96650 8678 96676 8730
rect 96380 8676 96436 8678
rect 96460 8676 96516 8678
rect 96540 8676 96596 8678
rect 96620 8676 96676 8678
rect 96380 7642 96436 7644
rect 96460 7642 96516 7644
rect 96540 7642 96596 7644
rect 96620 7642 96676 7644
rect 96380 7590 96406 7642
rect 96406 7590 96436 7642
rect 96460 7590 96470 7642
rect 96470 7590 96516 7642
rect 96540 7590 96586 7642
rect 96586 7590 96596 7642
rect 96620 7590 96650 7642
rect 96650 7590 96676 7642
rect 96380 7588 96436 7590
rect 96460 7588 96516 7590
rect 96540 7588 96596 7590
rect 96620 7588 96676 7590
rect 96380 6554 96436 6556
rect 96460 6554 96516 6556
rect 96540 6554 96596 6556
rect 96620 6554 96676 6556
rect 96380 6502 96406 6554
rect 96406 6502 96436 6554
rect 96460 6502 96470 6554
rect 96470 6502 96516 6554
rect 96540 6502 96586 6554
rect 96586 6502 96596 6554
rect 96620 6502 96650 6554
rect 96650 6502 96676 6554
rect 96380 6500 96436 6502
rect 96460 6500 96516 6502
rect 96540 6500 96596 6502
rect 96620 6500 96676 6502
rect 96380 5466 96436 5468
rect 96460 5466 96516 5468
rect 96540 5466 96596 5468
rect 96620 5466 96676 5468
rect 96380 5414 96406 5466
rect 96406 5414 96436 5466
rect 96460 5414 96470 5466
rect 96470 5414 96516 5466
rect 96540 5414 96586 5466
rect 96586 5414 96596 5466
rect 96620 5414 96650 5466
rect 96650 5414 96676 5466
rect 96380 5412 96436 5414
rect 96460 5412 96516 5414
rect 96540 5412 96596 5414
rect 96620 5412 96676 5414
rect 96380 4378 96436 4380
rect 96460 4378 96516 4380
rect 96540 4378 96596 4380
rect 96620 4378 96676 4380
rect 96380 4326 96406 4378
rect 96406 4326 96436 4378
rect 96460 4326 96470 4378
rect 96470 4326 96516 4378
rect 96540 4326 96586 4378
rect 96586 4326 96596 4378
rect 96620 4326 96650 4378
rect 96650 4326 96676 4378
rect 96380 4324 96436 4326
rect 96460 4324 96516 4326
rect 96540 4324 96596 4326
rect 96620 4324 96676 4326
rect 96380 3290 96436 3292
rect 96460 3290 96516 3292
rect 96540 3290 96596 3292
rect 96620 3290 96676 3292
rect 96380 3238 96406 3290
rect 96406 3238 96436 3290
rect 96460 3238 96470 3290
rect 96470 3238 96516 3290
rect 96540 3238 96586 3290
rect 96586 3238 96596 3290
rect 96620 3238 96650 3290
rect 96650 3238 96676 3290
rect 96380 3236 96436 3238
rect 96460 3236 96516 3238
rect 96540 3236 96596 3238
rect 96620 3236 96676 3238
rect 96380 2202 96436 2204
rect 96460 2202 96516 2204
rect 96540 2202 96596 2204
rect 96620 2202 96676 2204
rect 96380 2150 96406 2202
rect 96406 2150 96436 2202
rect 96460 2150 96470 2202
rect 96470 2150 96516 2202
rect 96540 2150 96586 2202
rect 96586 2150 96596 2202
rect 96620 2150 96650 2202
rect 96650 2150 96676 2202
rect 96380 2148 96436 2150
rect 96460 2148 96516 2150
rect 96540 2148 96596 2150
rect 96620 2148 96676 2150
rect 98090 15000 98146 15056
<< metal3 >>
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 50288 37568 50608 37569
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 37503 50608 37504
rect 81008 37568 81328 37569
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 37503 81328 37504
rect 68921 37362 68987 37365
rect 76833 37362 76899 37365
rect 68921 37360 76899 37362
rect 68921 37304 68926 37360
rect 68982 37304 76838 37360
rect 76894 37304 76899 37360
rect 68921 37302 76899 37304
rect 68921 37299 68987 37302
rect 76833 37299 76899 37302
rect 69565 37090 69631 37093
rect 70669 37090 70735 37093
rect 69565 37088 70735 37090
rect 69565 37032 69570 37088
rect 69626 37032 70674 37088
rect 70730 37032 70735 37088
rect 69565 37030 70735 37032
rect 69565 37027 69631 37030
rect 70669 37027 70735 37030
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 65648 37024 65968 37025
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 36959 65968 36960
rect 96368 37024 96688 37025
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 36959 96688 36960
rect 42149 36954 42215 36957
rect 48497 36954 48563 36957
rect 76097 36954 76163 36957
rect 42149 36952 48563 36954
rect 42149 36896 42154 36952
rect 42210 36896 48502 36952
rect 48558 36896 48563 36952
rect 42149 36894 48563 36896
rect 42149 36891 42215 36894
rect 48497 36891 48563 36894
rect 70350 36952 76163 36954
rect 70350 36896 76102 36952
rect 76158 36896 76163 36952
rect 70350 36894 76163 36896
rect 3233 36818 3299 36821
rect 70350 36818 70410 36894
rect 76097 36891 76163 36894
rect 3233 36816 70410 36818
rect 3233 36760 3238 36816
rect 3294 36760 70410 36816
rect 3233 36758 70410 36760
rect 70485 36818 70551 36821
rect 73429 36818 73495 36821
rect 70485 36816 73495 36818
rect 70485 36760 70490 36816
rect 70546 36760 73434 36816
rect 73490 36760 73495 36816
rect 70485 36758 73495 36760
rect 3233 36755 3299 36758
rect 70485 36755 70551 36758
rect 73429 36755 73495 36758
rect 49693 36682 49759 36685
rect 97625 36682 97691 36685
rect 49693 36680 97691 36682
rect 49693 36624 49698 36680
rect 49754 36624 97630 36680
rect 97686 36624 97691 36680
rect 49693 36622 97691 36624
rect 49693 36619 49759 36622
rect 97625 36619 97691 36622
rect 39941 36546 40007 36549
rect 41505 36546 41571 36549
rect 39941 36544 41571 36546
rect 39941 36488 39946 36544
rect 40002 36488 41510 36544
rect 41566 36488 41571 36544
rect 39941 36486 41571 36488
rect 39941 36483 40007 36486
rect 41505 36483 41571 36486
rect 43345 36546 43411 36549
rect 47761 36546 47827 36549
rect 43345 36544 47827 36546
rect 43345 36488 43350 36544
rect 43406 36488 47766 36544
rect 47822 36488 47827 36544
rect 43345 36486 47827 36488
rect 43345 36483 43411 36486
rect 47761 36483 47827 36486
rect 59813 36546 59879 36549
rect 65793 36546 65859 36549
rect 59813 36544 65859 36546
rect 59813 36488 59818 36544
rect 59874 36488 65798 36544
rect 65854 36488 65859 36544
rect 59813 36486 65859 36488
rect 59813 36483 59879 36486
rect 65793 36483 65859 36486
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 50288 36480 50608 36481
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 36415 50608 36416
rect 81008 36480 81328 36481
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 36415 81328 36416
rect 43437 36410 43503 36413
rect 47393 36410 47459 36413
rect 43437 36408 47459 36410
rect 43437 36352 43442 36408
rect 43498 36352 47398 36408
rect 47454 36352 47459 36408
rect 43437 36350 47459 36352
rect 43437 36347 43503 36350
rect 47393 36347 47459 36350
rect 70485 36410 70551 36413
rect 72049 36410 72115 36413
rect 70485 36408 72115 36410
rect 70485 36352 70490 36408
rect 70546 36352 72054 36408
rect 72110 36352 72115 36408
rect 70485 36350 72115 36352
rect 70485 36347 70551 36350
rect 72049 36347 72115 36350
rect 41413 36274 41479 36277
rect 48405 36274 48471 36277
rect 41413 36272 48471 36274
rect 41413 36216 41418 36272
rect 41474 36216 48410 36272
rect 48466 36216 48471 36272
rect 41413 36214 48471 36216
rect 41413 36211 41479 36214
rect 48405 36211 48471 36214
rect 54845 36274 54911 36277
rect 55857 36274 55923 36277
rect 54845 36272 55923 36274
rect 54845 36216 54850 36272
rect 54906 36216 55862 36272
rect 55918 36216 55923 36272
rect 54845 36214 55923 36216
rect 54845 36211 54911 36214
rect 55857 36211 55923 36214
rect 70209 36274 70275 36277
rect 75269 36274 75335 36277
rect 70209 36272 75335 36274
rect 70209 36216 70214 36272
rect 70270 36216 75274 36272
rect 75330 36216 75335 36272
rect 70209 36214 75335 36216
rect 70209 36211 70275 36214
rect 75269 36211 75335 36214
rect 28717 36138 28783 36141
rect 84653 36138 84719 36141
rect 28717 36136 84719 36138
rect 28717 36080 28722 36136
rect 28778 36080 84658 36136
rect 84714 36080 84719 36136
rect 28717 36078 84719 36080
rect 28717 36075 28783 36078
rect 84653 36075 84719 36078
rect 48589 36002 48655 36005
rect 55949 36002 56015 36005
rect 48589 36000 56015 36002
rect 48589 35944 48594 36000
rect 48650 35944 55954 36000
rect 56010 35944 56015 36000
rect 48589 35942 56015 35944
rect 48589 35939 48655 35942
rect 55949 35939 56015 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 65648 35936 65968 35937
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 35871 65968 35872
rect 96368 35936 96688 35937
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 35871 96688 35872
rect 39665 35730 39731 35733
rect 46749 35730 46815 35733
rect 39665 35728 46815 35730
rect 39665 35672 39670 35728
rect 39726 35672 46754 35728
rect 46810 35672 46815 35728
rect 39665 35670 46815 35672
rect 39665 35667 39731 35670
rect 46749 35667 46815 35670
rect 55305 35730 55371 35733
rect 57237 35730 57303 35733
rect 55305 35728 57303 35730
rect 55305 35672 55310 35728
rect 55366 35672 57242 35728
rect 57298 35672 57303 35728
rect 55305 35670 57303 35672
rect 55305 35667 55371 35670
rect 57237 35667 57303 35670
rect 39297 35594 39363 35597
rect 41413 35594 41479 35597
rect 39297 35592 41479 35594
rect 39297 35536 39302 35592
rect 39358 35536 41418 35592
rect 41474 35536 41479 35592
rect 39297 35534 41479 35536
rect 39297 35531 39363 35534
rect 41413 35531 41479 35534
rect 55305 35594 55371 35597
rect 55857 35594 55923 35597
rect 55305 35592 55923 35594
rect 55305 35536 55310 35592
rect 55366 35536 55862 35592
rect 55918 35536 55923 35592
rect 55305 35534 55923 35536
rect 55305 35531 55371 35534
rect 55857 35531 55923 35534
rect 35985 35458 36051 35461
rect 37273 35458 37339 35461
rect 35985 35456 37339 35458
rect 35985 35400 35990 35456
rect 36046 35400 37278 35456
rect 37334 35400 37339 35456
rect 35985 35398 37339 35400
rect 35985 35395 36051 35398
rect 37273 35395 37339 35398
rect 54753 35458 54819 35461
rect 55765 35458 55831 35461
rect 56777 35458 56843 35461
rect 54753 35456 56843 35458
rect 54753 35400 54758 35456
rect 54814 35400 55770 35456
rect 55826 35400 56782 35456
rect 56838 35400 56843 35456
rect 54753 35398 56843 35400
rect 54753 35395 54819 35398
rect 55765 35395 55831 35398
rect 56777 35395 56843 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 50288 35392 50608 35393
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 35327 50608 35328
rect 81008 35392 81328 35393
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 35327 81328 35328
rect 41321 35322 41387 35325
rect 47301 35322 47367 35325
rect 41321 35320 47367 35322
rect 41321 35264 41326 35320
rect 41382 35264 47306 35320
rect 47362 35264 47367 35320
rect 41321 35262 47367 35264
rect 41321 35259 41387 35262
rect 47301 35259 47367 35262
rect 39481 35186 39547 35189
rect 43621 35186 43687 35189
rect 39481 35184 43687 35186
rect 39481 35128 39486 35184
rect 39542 35128 43626 35184
rect 43682 35128 43687 35184
rect 39481 35126 43687 35128
rect 39481 35123 39547 35126
rect 43621 35123 43687 35126
rect 52177 35186 52243 35189
rect 57421 35186 57487 35189
rect 52177 35184 57487 35186
rect 52177 35128 52182 35184
rect 52238 35128 57426 35184
rect 57482 35128 57487 35184
rect 52177 35126 57487 35128
rect 52177 35123 52243 35126
rect 57421 35123 57487 35126
rect 62021 35186 62087 35189
rect 63125 35186 63191 35189
rect 62021 35184 63191 35186
rect 62021 35128 62026 35184
rect 62082 35128 63130 35184
rect 63186 35128 63191 35184
rect 62021 35126 63191 35128
rect 62021 35123 62087 35126
rect 63125 35123 63191 35126
rect 41321 35050 41387 35053
rect 44265 35050 44331 35053
rect 49877 35050 49943 35053
rect 41321 35048 44331 35050
rect 41321 34992 41326 35048
rect 41382 34992 44270 35048
rect 44326 34992 44331 35048
rect 41321 34990 44331 34992
rect 41321 34987 41387 34990
rect 44265 34987 44331 34990
rect 48270 35048 49943 35050
rect 48270 34992 49882 35048
rect 49938 34992 49943 35048
rect 48270 34990 49943 34992
rect 43345 34914 43411 34917
rect 48270 34914 48330 34990
rect 49877 34987 49943 34990
rect 61193 35050 61259 35053
rect 62573 35050 62639 35053
rect 61193 35048 62639 35050
rect 61193 34992 61198 35048
rect 61254 34992 62578 35048
rect 62634 34992 62639 35048
rect 61193 34990 62639 34992
rect 61193 34987 61259 34990
rect 62573 34987 62639 34990
rect 43345 34912 48330 34914
rect 43345 34856 43350 34912
rect 43406 34856 48330 34912
rect 43345 34854 48330 34856
rect 43345 34851 43411 34854
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 65648 34848 65968 34849
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 34783 65968 34784
rect 96368 34848 96688 34849
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 34783 96688 34784
rect 13261 34642 13327 34645
rect 83733 34642 83799 34645
rect 13261 34640 83799 34642
rect 13261 34584 13266 34640
rect 13322 34584 83738 34640
rect 83794 34584 83799 34640
rect 13261 34582 83799 34584
rect 13261 34579 13327 34582
rect 83733 34579 83799 34582
rect 33869 34506 33935 34509
rect 38653 34506 38719 34509
rect 33869 34504 38719 34506
rect 33869 34448 33874 34504
rect 33930 34448 38658 34504
rect 38714 34448 38719 34504
rect 33869 34446 38719 34448
rect 33869 34443 33935 34446
rect 38653 34443 38719 34446
rect 50981 34506 51047 34509
rect 51165 34506 51231 34509
rect 50981 34504 51231 34506
rect 50981 34448 50986 34504
rect 51042 34448 51170 34504
rect 51226 34448 51231 34504
rect 50981 34446 51231 34448
rect 50981 34443 51047 34446
rect 51165 34443 51231 34446
rect 54569 34506 54635 34509
rect 55305 34506 55371 34509
rect 54569 34504 55371 34506
rect 54569 34448 54574 34504
rect 54630 34448 55310 34504
rect 55366 34448 55371 34504
rect 54569 34446 55371 34448
rect 54569 34443 54635 34446
rect 55305 34443 55371 34446
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 50288 34304 50608 34305
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 34239 50608 34240
rect 81008 34304 81328 34305
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 34239 81328 34240
rect 38193 34234 38259 34237
rect 41505 34234 41571 34237
rect 38193 34232 41571 34234
rect 38193 34176 38198 34232
rect 38254 34176 41510 34232
rect 41566 34176 41571 34232
rect 38193 34174 41571 34176
rect 38193 34171 38259 34174
rect 41505 34171 41571 34174
rect 45461 34098 45527 34101
rect 47301 34098 47367 34101
rect 45461 34096 47367 34098
rect 45461 34040 45466 34096
rect 45522 34040 47306 34096
rect 47362 34040 47367 34096
rect 45461 34038 47367 34040
rect 45461 34035 45527 34038
rect 47301 34035 47367 34038
rect 50889 34098 50955 34101
rect 55029 34098 55095 34101
rect 50889 34096 55095 34098
rect 50889 34040 50894 34096
rect 50950 34040 55034 34096
rect 55090 34040 55095 34096
rect 50889 34038 55095 34040
rect 50889 34035 50955 34038
rect 55029 34035 55095 34038
rect 15009 33962 15075 33965
rect 67081 33962 67147 33965
rect 15009 33960 67147 33962
rect 15009 33904 15014 33960
rect 15070 33904 67086 33960
rect 67142 33904 67147 33960
rect 15009 33902 67147 33904
rect 15009 33899 15075 33902
rect 67081 33899 67147 33902
rect 40861 33826 40927 33829
rect 46473 33826 46539 33829
rect 62665 33826 62731 33829
rect 40861 33824 62731 33826
rect 40861 33768 40866 33824
rect 40922 33768 46478 33824
rect 46534 33768 62670 33824
rect 62726 33768 62731 33824
rect 40861 33766 62731 33768
rect 40861 33763 40927 33766
rect 46473 33763 46539 33766
rect 62665 33763 62731 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 65648 33760 65968 33761
rect 65648 33696 65656 33760
rect 65720 33696 65736 33760
rect 65800 33696 65816 33760
rect 65880 33696 65896 33760
rect 65960 33696 65968 33760
rect 65648 33695 65968 33696
rect 96368 33760 96688 33761
rect 96368 33696 96376 33760
rect 96440 33696 96456 33760
rect 96520 33696 96536 33760
rect 96600 33696 96616 33760
rect 96680 33696 96688 33760
rect 96368 33695 96688 33696
rect 30189 33690 30255 33693
rect 34237 33690 34303 33693
rect 30189 33688 34303 33690
rect 30189 33632 30194 33688
rect 30250 33632 34242 33688
rect 34298 33632 34303 33688
rect 30189 33630 34303 33632
rect 30189 33627 30255 33630
rect 34237 33627 34303 33630
rect 39941 33690 40007 33693
rect 41321 33690 41387 33693
rect 39941 33688 41387 33690
rect 39941 33632 39946 33688
rect 40002 33632 41326 33688
rect 41382 33632 41387 33688
rect 39941 33630 41387 33632
rect 39941 33627 40007 33630
rect 41321 33627 41387 33630
rect 54477 33690 54543 33693
rect 55305 33690 55371 33693
rect 54477 33688 55371 33690
rect 54477 33632 54482 33688
rect 54538 33632 55310 33688
rect 55366 33632 55371 33688
rect 54477 33630 55371 33632
rect 54477 33627 54543 33630
rect 55305 33627 55371 33630
rect 60365 33690 60431 33693
rect 61285 33690 61351 33693
rect 60365 33688 61351 33690
rect 60365 33632 60370 33688
rect 60426 33632 61290 33688
rect 61346 33632 61351 33688
rect 60365 33630 61351 33632
rect 60365 33627 60431 33630
rect 61285 33627 61351 33630
rect 17585 33554 17651 33557
rect 90357 33554 90423 33557
rect 17585 33552 90423 33554
rect 17585 33496 17590 33552
rect 17646 33496 90362 33552
rect 90418 33496 90423 33552
rect 17585 33494 90423 33496
rect 17585 33491 17651 33494
rect 90357 33491 90423 33494
rect 30005 33418 30071 33421
rect 30925 33418 30991 33421
rect 30005 33416 30991 33418
rect 30005 33360 30010 33416
rect 30066 33360 30930 33416
rect 30986 33360 30991 33416
rect 30005 33358 30991 33360
rect 30005 33355 30071 33358
rect 30925 33355 30991 33358
rect 40125 33418 40191 33421
rect 43713 33418 43779 33421
rect 40125 33416 43779 33418
rect 40125 33360 40130 33416
rect 40186 33360 43718 33416
rect 43774 33360 43779 33416
rect 40125 33358 43779 33360
rect 40125 33355 40191 33358
rect 43713 33355 43779 33358
rect 43989 33418 44055 33421
rect 89897 33418 89963 33421
rect 43989 33416 89963 33418
rect 43989 33360 43994 33416
rect 44050 33360 89902 33416
rect 89958 33360 89963 33416
rect 43989 33358 89963 33360
rect 43989 33355 44055 33358
rect 89897 33355 89963 33358
rect 30465 33282 30531 33285
rect 38009 33282 38075 33285
rect 30465 33280 38075 33282
rect 30465 33224 30470 33280
rect 30526 33224 38014 33280
rect 38070 33224 38075 33280
rect 30465 33222 38075 33224
rect 30465 33219 30531 33222
rect 38009 33219 38075 33222
rect 51073 33282 51139 33285
rect 60365 33282 60431 33285
rect 51073 33280 60431 33282
rect 51073 33224 51078 33280
rect 51134 33224 60370 33280
rect 60426 33224 60431 33280
rect 51073 33222 60431 33224
rect 51073 33219 51139 33222
rect 60365 33219 60431 33222
rect 60733 33282 60799 33285
rect 61469 33282 61535 33285
rect 60733 33280 61535 33282
rect 60733 33224 60738 33280
rect 60794 33224 61474 33280
rect 61530 33224 61535 33280
rect 60733 33222 61535 33224
rect 60733 33219 60799 33222
rect 61469 33219 61535 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 50288 33216 50608 33217
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 33151 50608 33152
rect 81008 33216 81328 33217
rect 81008 33152 81016 33216
rect 81080 33152 81096 33216
rect 81160 33152 81176 33216
rect 81240 33152 81256 33216
rect 81320 33152 81328 33216
rect 81008 33151 81328 33152
rect 38929 33146 38995 33149
rect 41229 33146 41295 33149
rect 38929 33144 41295 33146
rect 38929 33088 38934 33144
rect 38990 33088 41234 33144
rect 41290 33088 41295 33144
rect 38929 33086 41295 33088
rect 38929 33083 38995 33086
rect 41229 33083 41295 33086
rect 42149 33146 42215 33149
rect 47301 33146 47367 33149
rect 42149 33144 47367 33146
rect 42149 33088 42154 33144
rect 42210 33088 47306 33144
rect 47362 33088 47367 33144
rect 42149 33086 47367 33088
rect 42149 33083 42215 33086
rect 47301 33083 47367 33086
rect 22001 33010 22067 33013
rect 22185 33010 22251 33013
rect 22001 33008 22251 33010
rect 22001 32952 22006 33008
rect 22062 32952 22190 33008
rect 22246 32952 22251 33008
rect 22001 32950 22251 32952
rect 22001 32947 22067 32950
rect 22185 32947 22251 32950
rect 39573 33010 39639 33013
rect 45461 33010 45527 33013
rect 47209 33010 47275 33013
rect 39573 33008 47275 33010
rect 39573 32952 39578 33008
rect 39634 32952 45466 33008
rect 45522 32952 47214 33008
rect 47270 32952 47275 33008
rect 39573 32950 47275 32952
rect 39573 32947 39639 32950
rect 45461 32947 45527 32950
rect 47209 32947 47275 32950
rect 49049 33010 49115 33013
rect 56133 33010 56199 33013
rect 49049 33008 56199 33010
rect 49049 32952 49054 33008
rect 49110 32952 56138 33008
rect 56194 32952 56199 33008
rect 49049 32950 56199 32952
rect 49049 32947 49115 32950
rect 56133 32947 56199 32950
rect 39389 32874 39455 32877
rect 46565 32874 46631 32877
rect 39389 32872 46631 32874
rect 39389 32816 39394 32872
rect 39450 32816 46570 32872
rect 46626 32816 46631 32872
rect 39389 32814 46631 32816
rect 39389 32811 39455 32814
rect 46565 32811 46631 32814
rect 38653 32738 38719 32741
rect 40677 32738 40743 32741
rect 38653 32736 40743 32738
rect 38653 32680 38658 32736
rect 38714 32680 40682 32736
rect 40738 32680 40743 32736
rect 38653 32678 40743 32680
rect 38653 32675 38719 32678
rect 40677 32675 40743 32678
rect 50613 32738 50679 32741
rect 51073 32738 51139 32741
rect 50613 32736 51139 32738
rect 50613 32680 50618 32736
rect 50674 32680 51078 32736
rect 51134 32680 51139 32736
rect 50613 32678 51139 32680
rect 50613 32675 50679 32678
rect 51073 32675 51139 32678
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 65648 32672 65968 32673
rect 65648 32608 65656 32672
rect 65720 32608 65736 32672
rect 65800 32608 65816 32672
rect 65880 32608 65896 32672
rect 65960 32608 65968 32672
rect 65648 32607 65968 32608
rect 96368 32672 96688 32673
rect 96368 32608 96376 32672
rect 96440 32608 96456 32672
rect 96520 32608 96536 32672
rect 96600 32608 96616 32672
rect 96680 32608 96688 32672
rect 96368 32607 96688 32608
rect 41965 32602 42031 32605
rect 42701 32602 42767 32605
rect 41965 32600 42767 32602
rect 41965 32544 41970 32600
rect 42026 32544 42706 32600
rect 42762 32544 42767 32600
rect 41965 32542 42767 32544
rect 41965 32539 42031 32542
rect 42701 32539 42767 32542
rect 22369 32330 22435 32333
rect 26969 32330 27035 32333
rect 22369 32328 27035 32330
rect 22369 32272 22374 32328
rect 22430 32272 26974 32328
rect 27030 32272 27035 32328
rect 22369 32270 27035 32272
rect 22369 32267 22435 32270
rect 26969 32267 27035 32270
rect 39941 32330 40007 32333
rect 44173 32330 44239 32333
rect 39941 32328 44239 32330
rect 39941 32272 39946 32328
rect 40002 32272 44178 32328
rect 44234 32272 44239 32328
rect 39941 32270 44239 32272
rect 39941 32267 40007 32270
rect 44173 32267 44239 32270
rect 50981 32194 51047 32197
rect 57973 32194 58039 32197
rect 50981 32192 58039 32194
rect 50981 32136 50986 32192
rect 51042 32136 57978 32192
rect 58034 32136 58039 32192
rect 50981 32134 58039 32136
rect 50981 32131 51047 32134
rect 57973 32131 58039 32134
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 50288 32128 50608 32129
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 32063 50608 32064
rect 81008 32128 81328 32129
rect 81008 32064 81016 32128
rect 81080 32064 81096 32128
rect 81160 32064 81176 32128
rect 81240 32064 81256 32128
rect 81320 32064 81328 32128
rect 81008 32063 81328 32064
rect 57881 32058 57947 32061
rect 58801 32058 58867 32061
rect 57881 32056 58867 32058
rect 57881 32000 57886 32056
rect 57942 32000 58806 32056
rect 58862 32000 58867 32056
rect 57881 31998 58867 32000
rect 57881 31995 57947 31998
rect 58801 31995 58867 31998
rect 57513 31922 57579 31925
rect 58157 31922 58223 31925
rect 57513 31920 58223 31922
rect 57513 31864 57518 31920
rect 57574 31864 58162 31920
rect 58218 31864 58223 31920
rect 57513 31862 58223 31864
rect 57513 31859 57579 31862
rect 58157 31859 58223 31862
rect 48405 31786 48471 31789
rect 57881 31786 57947 31789
rect 48405 31784 57947 31786
rect 48405 31728 48410 31784
rect 48466 31728 57886 31784
rect 57942 31728 57947 31784
rect 48405 31726 57947 31728
rect 48405 31723 48471 31726
rect 57881 31723 57947 31726
rect 24025 31650 24091 31653
rect 27521 31650 27587 31653
rect 24025 31648 27587 31650
rect 24025 31592 24030 31648
rect 24086 31592 27526 31648
rect 27582 31592 27587 31648
rect 24025 31590 27587 31592
rect 24025 31587 24091 31590
rect 27521 31587 27587 31590
rect 52177 31650 52243 31653
rect 54201 31650 54267 31653
rect 56777 31650 56843 31653
rect 52177 31648 56843 31650
rect 52177 31592 52182 31648
rect 52238 31592 54206 31648
rect 54262 31592 56782 31648
rect 56838 31592 56843 31648
rect 52177 31590 56843 31592
rect 52177 31587 52243 31590
rect 54201 31587 54267 31590
rect 56777 31587 56843 31590
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 65648 31584 65968 31585
rect 65648 31520 65656 31584
rect 65720 31520 65736 31584
rect 65800 31520 65816 31584
rect 65880 31520 65896 31584
rect 65960 31520 65968 31584
rect 65648 31519 65968 31520
rect 96368 31584 96688 31585
rect 96368 31520 96376 31584
rect 96440 31520 96456 31584
rect 96520 31520 96536 31584
rect 96600 31520 96616 31584
rect 96680 31520 96688 31584
rect 96368 31519 96688 31520
rect 18965 31378 19031 31381
rect 19609 31378 19675 31381
rect 18965 31376 19675 31378
rect 18965 31320 18970 31376
rect 19026 31320 19614 31376
rect 19670 31320 19675 31376
rect 18965 31318 19675 31320
rect 18965 31315 19031 31318
rect 19609 31315 19675 31318
rect 27521 31378 27587 31381
rect 28349 31378 28415 31381
rect 27521 31376 28415 31378
rect 27521 31320 27526 31376
rect 27582 31320 28354 31376
rect 28410 31320 28415 31376
rect 27521 31318 28415 31320
rect 27521 31315 27587 31318
rect 28349 31315 28415 31318
rect 59721 31378 59787 31381
rect 60641 31378 60707 31381
rect 59721 31376 60707 31378
rect 59721 31320 59726 31376
rect 59782 31320 60646 31376
rect 60702 31320 60707 31376
rect 59721 31318 60707 31320
rect 59721 31315 59787 31318
rect 60641 31315 60707 31318
rect 28073 31242 28139 31245
rect 97533 31242 97599 31245
rect 28073 31240 97599 31242
rect 28073 31184 28078 31240
rect 28134 31184 97538 31240
rect 97594 31184 97599 31240
rect 28073 31182 97599 31184
rect 28073 31179 28139 31182
rect 97533 31179 97599 31182
rect 20069 31106 20135 31109
rect 28165 31106 28231 31109
rect 20069 31104 28231 31106
rect 20069 31048 20074 31104
rect 20130 31048 28170 31104
rect 28226 31048 28231 31104
rect 20069 31046 28231 31048
rect 20069 31043 20135 31046
rect 28165 31043 28231 31046
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 50288 31040 50608 31041
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 30975 50608 30976
rect 81008 31040 81328 31041
rect 81008 30976 81016 31040
rect 81080 30976 81096 31040
rect 81160 30976 81176 31040
rect 81240 30976 81256 31040
rect 81320 30976 81328 31040
rect 81008 30975 81328 30976
rect 26877 30834 26943 30837
rect 28349 30834 28415 30837
rect 26877 30832 28415 30834
rect 26877 30776 26882 30832
rect 26938 30776 28354 30832
rect 28410 30776 28415 30832
rect 26877 30774 28415 30776
rect 26877 30771 26943 30774
rect 28349 30771 28415 30774
rect 33869 30834 33935 30837
rect 36261 30834 36327 30837
rect 33869 30832 36327 30834
rect 33869 30776 33874 30832
rect 33930 30776 36266 30832
rect 36322 30776 36327 30832
rect 33869 30774 36327 30776
rect 33869 30771 33935 30774
rect 36261 30771 36327 30774
rect 46289 30834 46355 30837
rect 47209 30834 47275 30837
rect 46289 30832 47275 30834
rect 46289 30776 46294 30832
rect 46350 30776 47214 30832
rect 47270 30776 47275 30832
rect 46289 30774 47275 30776
rect 46289 30771 46355 30774
rect 47209 30771 47275 30774
rect 31293 30698 31359 30701
rect 80053 30698 80119 30701
rect 31293 30696 80119 30698
rect 31293 30640 31298 30696
rect 31354 30640 80058 30696
rect 80114 30640 80119 30696
rect 31293 30638 80119 30640
rect 31293 30635 31359 30638
rect 80053 30635 80119 30638
rect 43529 30562 43595 30565
rect 46657 30562 46723 30565
rect 43529 30560 46723 30562
rect 43529 30504 43534 30560
rect 43590 30504 46662 30560
rect 46718 30504 46723 30560
rect 43529 30502 46723 30504
rect 43529 30499 43595 30502
rect 46657 30499 46723 30502
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 65648 30496 65968 30497
rect 65648 30432 65656 30496
rect 65720 30432 65736 30496
rect 65800 30432 65816 30496
rect 65880 30432 65896 30496
rect 65960 30432 65968 30496
rect 65648 30431 65968 30432
rect 96368 30496 96688 30497
rect 96368 30432 96376 30496
rect 96440 30432 96456 30496
rect 96520 30432 96536 30496
rect 96600 30432 96616 30496
rect 96680 30432 96688 30496
rect 96368 30431 96688 30432
rect 53833 30426 53899 30429
rect 55029 30426 55095 30429
rect 53833 30424 55095 30426
rect 53833 30368 53838 30424
rect 53894 30368 55034 30424
rect 55090 30368 55095 30424
rect 53833 30366 55095 30368
rect 53833 30363 53899 30366
rect 55029 30363 55095 30366
rect 54201 30290 54267 30293
rect 56593 30290 56659 30293
rect 54201 30288 56659 30290
rect 54201 30232 54206 30288
rect 54262 30232 56598 30288
rect 56654 30232 56659 30288
rect 54201 30230 56659 30232
rect 54201 30227 54267 30230
rect 56593 30227 56659 30230
rect 46105 30154 46171 30157
rect 46657 30154 46723 30157
rect 46105 30152 46723 30154
rect 46105 30096 46110 30152
rect 46166 30096 46662 30152
rect 46718 30096 46723 30152
rect 46105 30094 46723 30096
rect 46105 30091 46171 30094
rect 46657 30091 46723 30094
rect 52269 30154 52335 30157
rect 62757 30154 62823 30157
rect 52269 30152 62823 30154
rect 52269 30096 52274 30152
rect 52330 30096 62762 30152
rect 62818 30096 62823 30152
rect 52269 30094 62823 30096
rect 52269 30091 52335 30094
rect 62757 30091 62823 30094
rect 43345 30018 43411 30021
rect 46933 30018 46999 30021
rect 43345 30016 46999 30018
rect 43345 29960 43350 30016
rect 43406 29960 46938 30016
rect 46994 29960 46999 30016
rect 43345 29958 46999 29960
rect 43345 29955 43411 29958
rect 46933 29955 46999 29958
rect 54661 30018 54727 30021
rect 57145 30018 57211 30021
rect 54661 30016 57211 30018
rect 54661 29960 54666 30016
rect 54722 29960 57150 30016
rect 57206 29960 57211 30016
rect 54661 29958 57211 29960
rect 54661 29955 54727 29958
rect 57145 29955 57211 29958
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 50288 29952 50608 29953
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 29887 50608 29888
rect 81008 29952 81328 29953
rect 81008 29888 81016 29952
rect 81080 29888 81096 29952
rect 81160 29888 81176 29952
rect 81240 29888 81256 29952
rect 81320 29888 81328 29952
rect 81008 29887 81328 29888
rect 45921 29882 45987 29885
rect 47577 29882 47643 29885
rect 45921 29880 47643 29882
rect 45921 29824 45926 29880
rect 45982 29824 47582 29880
rect 47638 29824 47643 29880
rect 45921 29822 47643 29824
rect 45921 29819 45987 29822
rect 47577 29819 47643 29822
rect 45829 29746 45895 29749
rect 47301 29746 47367 29749
rect 45829 29744 47367 29746
rect 45829 29688 45834 29744
rect 45890 29688 47306 29744
rect 47362 29688 47367 29744
rect 45829 29686 47367 29688
rect 45829 29683 45895 29686
rect 47301 29683 47367 29686
rect 2497 29610 2563 29613
rect 52361 29610 52427 29613
rect 2497 29608 52427 29610
rect 2497 29552 2502 29608
rect 2558 29552 52366 29608
rect 52422 29552 52427 29608
rect 2497 29550 52427 29552
rect 2497 29547 2563 29550
rect 52361 29547 52427 29550
rect 58525 29610 58591 29613
rect 65609 29610 65675 29613
rect 58525 29608 65675 29610
rect 58525 29552 58530 29608
rect 58586 29552 65614 29608
rect 65670 29552 65675 29608
rect 58525 29550 65675 29552
rect 58525 29547 58591 29550
rect 65609 29547 65675 29550
rect 66529 29610 66595 29613
rect 67449 29610 67515 29613
rect 66529 29608 67515 29610
rect 66529 29552 66534 29608
rect 66590 29552 67454 29608
rect 67510 29552 67515 29608
rect 66529 29550 67515 29552
rect 66529 29547 66595 29550
rect 67449 29547 67515 29550
rect 35709 29474 35775 29477
rect 38561 29474 38627 29477
rect 35709 29472 38627 29474
rect 35709 29416 35714 29472
rect 35770 29416 38566 29472
rect 38622 29416 38627 29472
rect 35709 29414 38627 29416
rect 35709 29411 35775 29414
rect 38561 29411 38627 29414
rect 43345 29474 43411 29477
rect 47209 29474 47275 29477
rect 43345 29472 47275 29474
rect 43345 29416 43350 29472
rect 43406 29416 47214 29472
rect 47270 29416 47275 29472
rect 43345 29414 47275 29416
rect 43345 29411 43411 29414
rect 47209 29411 47275 29414
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 65648 29408 65968 29409
rect 65648 29344 65656 29408
rect 65720 29344 65736 29408
rect 65800 29344 65816 29408
rect 65880 29344 65896 29408
rect 65960 29344 65968 29408
rect 65648 29343 65968 29344
rect 96368 29408 96688 29409
rect 96368 29344 96376 29408
rect 96440 29344 96456 29408
rect 96520 29344 96536 29408
rect 96600 29344 96616 29408
rect 96680 29344 96688 29408
rect 96368 29343 96688 29344
rect 68277 29202 68343 29205
rect 74073 29202 74139 29205
rect 68277 29200 74139 29202
rect 68277 29144 68282 29200
rect 68338 29144 74078 29200
rect 74134 29144 74139 29200
rect 68277 29142 74139 29144
rect 68277 29139 68343 29142
rect 74073 29139 74139 29142
rect 55305 29066 55371 29069
rect 56685 29066 56751 29069
rect 55305 29064 56751 29066
rect 55305 29008 55310 29064
rect 55366 29008 56690 29064
rect 56746 29008 56751 29064
rect 55305 29006 56751 29008
rect 55305 29003 55371 29006
rect 56685 29003 56751 29006
rect 67909 29066 67975 29069
rect 69381 29066 69447 29069
rect 67909 29064 69447 29066
rect 67909 29008 67914 29064
rect 67970 29008 69386 29064
rect 69442 29008 69447 29064
rect 67909 29006 69447 29008
rect 67909 29003 67975 29006
rect 69381 29003 69447 29006
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 50288 28864 50608 28865
rect 50288 28800 50296 28864
rect 50360 28800 50376 28864
rect 50440 28800 50456 28864
rect 50520 28800 50536 28864
rect 50600 28800 50608 28864
rect 50288 28799 50608 28800
rect 81008 28864 81328 28865
rect 81008 28800 81016 28864
rect 81080 28800 81096 28864
rect 81160 28800 81176 28864
rect 81240 28800 81256 28864
rect 81320 28800 81328 28864
rect 81008 28799 81328 28800
rect 15653 28794 15719 28797
rect 16021 28794 16087 28797
rect 15653 28792 16087 28794
rect 15653 28736 15658 28792
rect 15714 28736 16026 28792
rect 16082 28736 16087 28792
rect 15653 28734 16087 28736
rect 15653 28731 15719 28734
rect 16021 28731 16087 28734
rect 30005 28658 30071 28661
rect 37549 28658 37615 28661
rect 43529 28658 43595 28661
rect 30005 28656 43595 28658
rect 30005 28600 30010 28656
rect 30066 28600 37554 28656
rect 37610 28600 43534 28656
rect 43590 28600 43595 28656
rect 30005 28598 43595 28600
rect 30005 28595 30071 28598
rect 37549 28595 37615 28598
rect 43529 28595 43595 28598
rect 49417 28658 49483 28661
rect 50889 28658 50955 28661
rect 54109 28658 54175 28661
rect 49417 28656 54175 28658
rect 49417 28600 49422 28656
rect 49478 28600 50894 28656
rect 50950 28600 54114 28656
rect 54170 28600 54175 28656
rect 49417 28598 54175 28600
rect 49417 28595 49483 28598
rect 50889 28595 50955 28598
rect 54109 28595 54175 28598
rect 36997 28522 37063 28525
rect 37733 28522 37799 28525
rect 36997 28520 37799 28522
rect 36997 28464 37002 28520
rect 37058 28464 37738 28520
rect 37794 28464 37799 28520
rect 36997 28462 37799 28464
rect 36997 28459 37063 28462
rect 37733 28459 37799 28462
rect 42057 28522 42123 28525
rect 79501 28522 79567 28525
rect 42057 28520 79567 28522
rect 42057 28464 42062 28520
rect 42118 28464 79506 28520
rect 79562 28464 79567 28520
rect 42057 28462 79567 28464
rect 42057 28459 42123 28462
rect 79501 28459 79567 28462
rect 42425 28386 42491 28389
rect 50981 28386 51047 28389
rect 51165 28386 51231 28389
rect 42425 28384 51231 28386
rect 42425 28328 42430 28384
rect 42486 28328 50986 28384
rect 51042 28328 51170 28384
rect 51226 28328 51231 28384
rect 42425 28326 51231 28328
rect 42425 28323 42491 28326
rect 50981 28323 51047 28326
rect 51165 28323 51231 28326
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 65648 28320 65968 28321
rect 65648 28256 65656 28320
rect 65720 28256 65736 28320
rect 65800 28256 65816 28320
rect 65880 28256 65896 28320
rect 65960 28256 65968 28320
rect 65648 28255 65968 28256
rect 96368 28320 96688 28321
rect 96368 28256 96376 28320
rect 96440 28256 96456 28320
rect 96520 28256 96536 28320
rect 96600 28256 96616 28320
rect 96680 28256 96688 28320
rect 96368 28255 96688 28256
rect 20345 28250 20411 28253
rect 27889 28250 27955 28253
rect 20345 28248 27955 28250
rect 20345 28192 20350 28248
rect 20406 28192 27894 28248
rect 27950 28192 27955 28248
rect 20345 28190 27955 28192
rect 20345 28187 20411 28190
rect 27889 28187 27955 28190
rect 36169 28250 36235 28253
rect 41505 28250 41571 28253
rect 36169 28248 41571 28250
rect 36169 28192 36174 28248
rect 36230 28192 41510 28248
rect 41566 28192 41571 28248
rect 36169 28190 41571 28192
rect 36169 28187 36235 28190
rect 41505 28187 41571 28190
rect 18873 28114 18939 28117
rect 19057 28114 19123 28117
rect 18873 28112 19123 28114
rect 18873 28056 18878 28112
rect 18934 28056 19062 28112
rect 19118 28056 19123 28112
rect 18873 28054 19123 28056
rect 18873 28051 18939 28054
rect 19057 28051 19123 28054
rect 31753 28114 31819 28117
rect 40585 28114 40651 28117
rect 31753 28112 40651 28114
rect 31753 28056 31758 28112
rect 31814 28056 40590 28112
rect 40646 28056 40651 28112
rect 31753 28054 40651 28056
rect 31753 28051 31819 28054
rect 40585 28051 40651 28054
rect 46841 28114 46907 28117
rect 49969 28114 50035 28117
rect 46841 28112 50035 28114
rect 46841 28056 46846 28112
rect 46902 28056 49974 28112
rect 50030 28056 50035 28112
rect 46841 28054 50035 28056
rect 46841 28051 46907 28054
rect 49969 28051 50035 28054
rect 17125 27978 17191 27981
rect 18597 27978 18663 27981
rect 19149 27978 19215 27981
rect 91461 27978 91527 27981
rect 17125 27976 91527 27978
rect 17125 27920 17130 27976
rect 17186 27920 18602 27976
rect 18658 27920 19154 27976
rect 19210 27920 91466 27976
rect 91522 27920 91527 27976
rect 17125 27918 91527 27920
rect 17125 27915 17191 27918
rect 18597 27915 18663 27918
rect 19149 27915 19215 27918
rect 91461 27915 91527 27918
rect 21173 27842 21239 27845
rect 33593 27842 33659 27845
rect 40033 27842 40099 27845
rect 21173 27840 40099 27842
rect 21173 27784 21178 27840
rect 21234 27784 33598 27840
rect 33654 27784 40038 27840
rect 40094 27784 40099 27840
rect 21173 27782 40099 27784
rect 21173 27779 21239 27782
rect 33593 27779 33659 27782
rect 40033 27779 40099 27782
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 50288 27776 50608 27777
rect 50288 27712 50296 27776
rect 50360 27712 50376 27776
rect 50440 27712 50456 27776
rect 50520 27712 50536 27776
rect 50600 27712 50608 27776
rect 50288 27711 50608 27712
rect 81008 27776 81328 27777
rect 81008 27712 81016 27776
rect 81080 27712 81096 27776
rect 81160 27712 81176 27776
rect 81240 27712 81256 27776
rect 81320 27712 81328 27776
rect 81008 27711 81328 27712
rect 39297 27706 39363 27709
rect 46013 27706 46079 27709
rect 39297 27704 46079 27706
rect 39297 27648 39302 27704
rect 39358 27648 46018 27704
rect 46074 27648 46079 27704
rect 39297 27646 46079 27648
rect 39297 27643 39363 27646
rect 46013 27643 46079 27646
rect 51073 27706 51139 27709
rect 53925 27706 53991 27709
rect 51073 27704 53991 27706
rect 51073 27648 51078 27704
rect 51134 27648 53930 27704
rect 53986 27648 53991 27704
rect 51073 27646 53991 27648
rect 51073 27643 51139 27646
rect 53925 27643 53991 27646
rect 35893 27570 35959 27573
rect 39573 27570 39639 27573
rect 35893 27568 39639 27570
rect 35893 27512 35898 27568
rect 35954 27512 39578 27568
rect 39634 27512 39639 27568
rect 35893 27510 39639 27512
rect 35893 27507 35959 27510
rect 39573 27507 39639 27510
rect 41505 27570 41571 27573
rect 42609 27570 42675 27573
rect 50705 27570 50771 27573
rect 41505 27568 50771 27570
rect 41505 27512 41510 27568
rect 41566 27512 42614 27568
rect 42670 27512 50710 27568
rect 50766 27512 50771 27568
rect 41505 27510 50771 27512
rect 41505 27507 41571 27510
rect 42609 27507 42675 27510
rect 50705 27507 50771 27510
rect 27153 27434 27219 27437
rect 30465 27434 30531 27437
rect 27153 27432 30531 27434
rect 27153 27376 27158 27432
rect 27214 27376 30470 27432
rect 30526 27376 30531 27432
rect 27153 27374 30531 27376
rect 27153 27371 27219 27374
rect 30465 27371 30531 27374
rect 48681 27434 48747 27437
rect 53741 27434 53807 27437
rect 48681 27432 53807 27434
rect 48681 27376 48686 27432
rect 48742 27376 53746 27432
rect 53802 27376 53807 27432
rect 48681 27374 53807 27376
rect 48681 27371 48747 27374
rect 53741 27371 53807 27374
rect 40493 27298 40559 27301
rect 42517 27298 42583 27301
rect 40493 27296 42583 27298
rect 40493 27240 40498 27296
rect 40554 27240 42522 27296
rect 42578 27240 42583 27296
rect 40493 27238 42583 27240
rect 40493 27235 40559 27238
rect 42517 27235 42583 27238
rect 49233 27298 49299 27301
rect 53281 27298 53347 27301
rect 53649 27298 53715 27301
rect 49233 27296 53715 27298
rect 49233 27240 49238 27296
rect 49294 27240 53286 27296
rect 53342 27240 53654 27296
rect 53710 27240 53715 27296
rect 49233 27238 53715 27240
rect 49233 27235 49299 27238
rect 53281 27235 53347 27238
rect 53649 27235 53715 27238
rect 54109 27298 54175 27301
rect 56041 27298 56107 27301
rect 54109 27296 56107 27298
rect 54109 27240 54114 27296
rect 54170 27240 56046 27296
rect 56102 27240 56107 27296
rect 54109 27238 56107 27240
rect 54109 27235 54175 27238
rect 56041 27235 56107 27238
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 65648 27232 65968 27233
rect 65648 27168 65656 27232
rect 65720 27168 65736 27232
rect 65800 27168 65816 27232
rect 65880 27168 65896 27232
rect 65960 27168 65968 27232
rect 65648 27167 65968 27168
rect 96368 27232 96688 27233
rect 96368 27168 96376 27232
rect 96440 27168 96456 27232
rect 96520 27168 96536 27232
rect 96600 27168 96616 27232
rect 96680 27168 96688 27232
rect 96368 27167 96688 27168
rect 44081 27162 44147 27165
rect 46289 27162 46355 27165
rect 44081 27160 46355 27162
rect 44081 27104 44086 27160
rect 44142 27104 46294 27160
rect 46350 27104 46355 27160
rect 44081 27102 46355 27104
rect 44081 27099 44147 27102
rect 46289 27099 46355 27102
rect 50705 27162 50771 27165
rect 51441 27162 51507 27165
rect 55029 27162 55095 27165
rect 50705 27160 55095 27162
rect 50705 27104 50710 27160
rect 50766 27104 51446 27160
rect 51502 27104 55034 27160
rect 55090 27104 55095 27160
rect 50705 27102 55095 27104
rect 50705 27099 50771 27102
rect 51441 27099 51507 27102
rect 55029 27099 55095 27102
rect 21541 27026 21607 27029
rect 22277 27026 22343 27029
rect 21541 27024 22343 27026
rect 21541 26968 21546 27024
rect 21602 26968 22282 27024
rect 22338 26968 22343 27024
rect 21541 26966 22343 26968
rect 21541 26963 21607 26966
rect 22277 26963 22343 26966
rect 30465 27026 30531 27029
rect 36353 27026 36419 27029
rect 30465 27024 36419 27026
rect 30465 26968 30470 27024
rect 30526 26968 36358 27024
rect 36414 26968 36419 27024
rect 30465 26966 36419 26968
rect 30465 26963 30531 26966
rect 36353 26963 36419 26966
rect 59169 27026 59235 27029
rect 60917 27026 60983 27029
rect 59169 27024 60983 27026
rect 59169 26968 59174 27024
rect 59230 26968 60922 27024
rect 60978 26968 60983 27024
rect 59169 26966 60983 26968
rect 59169 26963 59235 26966
rect 60917 26963 60983 26966
rect 27797 26890 27863 26893
rect 36077 26890 36143 26893
rect 27797 26888 36143 26890
rect 27797 26832 27802 26888
rect 27858 26832 36082 26888
rect 36138 26832 36143 26888
rect 27797 26830 36143 26832
rect 27797 26827 27863 26830
rect 36077 26827 36143 26830
rect 52545 26890 52611 26893
rect 57513 26890 57579 26893
rect 52545 26888 57579 26890
rect 52545 26832 52550 26888
rect 52606 26832 57518 26888
rect 57574 26832 57579 26888
rect 52545 26830 57579 26832
rect 52545 26827 52611 26830
rect 57513 26827 57579 26830
rect 77385 26890 77451 26893
rect 78489 26890 78555 26893
rect 77385 26888 78555 26890
rect 77385 26832 77390 26888
rect 77446 26832 78494 26888
rect 78550 26832 78555 26888
rect 77385 26830 78555 26832
rect 77385 26827 77451 26830
rect 78489 26827 78555 26830
rect 33317 26754 33383 26757
rect 38929 26754 38995 26757
rect 41505 26754 41571 26757
rect 33317 26752 41571 26754
rect 33317 26696 33322 26752
rect 33378 26696 38934 26752
rect 38990 26696 41510 26752
rect 41566 26696 41571 26752
rect 33317 26694 41571 26696
rect 33317 26691 33383 26694
rect 38929 26691 38995 26694
rect 41505 26691 41571 26694
rect 77017 26754 77083 26757
rect 78121 26754 78187 26757
rect 77017 26752 78187 26754
rect 77017 26696 77022 26752
rect 77078 26696 78126 26752
rect 78182 26696 78187 26752
rect 77017 26694 78187 26696
rect 77017 26691 77083 26694
rect 78121 26691 78187 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 50288 26688 50608 26689
rect 50288 26624 50296 26688
rect 50360 26624 50376 26688
rect 50440 26624 50456 26688
rect 50520 26624 50536 26688
rect 50600 26624 50608 26688
rect 50288 26623 50608 26624
rect 81008 26688 81328 26689
rect 81008 26624 81016 26688
rect 81080 26624 81096 26688
rect 81160 26624 81176 26688
rect 81240 26624 81256 26688
rect 81320 26624 81328 26688
rect 81008 26623 81328 26624
rect 30373 26618 30439 26621
rect 36445 26618 36511 26621
rect 30373 26616 36511 26618
rect 30373 26560 30378 26616
rect 30434 26560 36450 26616
rect 36506 26560 36511 26616
rect 30373 26558 36511 26560
rect 30373 26555 30439 26558
rect 36445 26555 36511 26558
rect 37825 26618 37891 26621
rect 38510 26618 38516 26620
rect 37825 26616 38516 26618
rect 37825 26560 37830 26616
rect 37886 26560 38516 26616
rect 37825 26558 38516 26560
rect 37825 26555 37891 26558
rect 38510 26556 38516 26558
rect 38580 26618 38586 26620
rect 43345 26618 43411 26621
rect 38580 26616 43411 26618
rect 38580 26560 43350 26616
rect 43406 26560 43411 26616
rect 38580 26558 43411 26560
rect 38580 26556 38586 26558
rect 43345 26555 43411 26558
rect 55581 26618 55647 26621
rect 56225 26618 56291 26621
rect 55581 26616 56291 26618
rect 55581 26560 55586 26616
rect 55642 26560 56230 26616
rect 56286 26560 56291 26616
rect 55581 26558 56291 26560
rect 55581 26555 55647 26558
rect 56225 26555 56291 26558
rect 59261 26618 59327 26621
rect 60641 26618 60707 26621
rect 59261 26616 60707 26618
rect 59261 26560 59266 26616
rect 59322 26560 60646 26616
rect 60702 26560 60707 26616
rect 59261 26558 60707 26560
rect 59261 26555 59327 26558
rect 60641 26555 60707 26558
rect 20713 26482 20779 26485
rect 21541 26482 21607 26485
rect 20713 26480 21607 26482
rect 20713 26424 20718 26480
rect 20774 26424 21546 26480
rect 21602 26424 21607 26480
rect 20713 26422 21607 26424
rect 20713 26419 20779 26422
rect 21541 26419 21607 26422
rect 33685 26482 33751 26485
rect 36721 26482 36787 26485
rect 33685 26480 36787 26482
rect 33685 26424 33690 26480
rect 33746 26424 36726 26480
rect 36782 26424 36787 26480
rect 33685 26422 36787 26424
rect 33685 26419 33751 26422
rect 36721 26419 36787 26422
rect 40493 26482 40559 26485
rect 48313 26482 48379 26485
rect 40493 26480 48379 26482
rect 40493 26424 40498 26480
rect 40554 26424 48318 26480
rect 48374 26424 48379 26480
rect 40493 26422 48379 26424
rect 40493 26419 40559 26422
rect 48313 26419 48379 26422
rect 52545 26482 52611 26485
rect 53833 26482 53899 26485
rect 52545 26480 53899 26482
rect 52545 26424 52550 26480
rect 52606 26424 53838 26480
rect 53894 26424 53899 26480
rect 52545 26422 53899 26424
rect 52545 26419 52611 26422
rect 53833 26419 53899 26422
rect 60549 26482 60615 26485
rect 61193 26482 61259 26485
rect 60549 26480 61259 26482
rect 60549 26424 60554 26480
rect 60610 26424 61198 26480
rect 61254 26424 61259 26480
rect 60549 26422 61259 26424
rect 60549 26419 60615 26422
rect 61193 26419 61259 26422
rect 33685 26346 33751 26349
rect 36721 26346 36787 26349
rect 33685 26344 36787 26346
rect 33685 26288 33690 26344
rect 33746 26288 36726 26344
rect 36782 26288 36787 26344
rect 33685 26286 36787 26288
rect 33685 26283 33751 26286
rect 36721 26283 36787 26286
rect 41045 26346 41111 26349
rect 42333 26346 42399 26349
rect 41045 26344 42399 26346
rect 41045 26288 41050 26344
rect 41106 26288 42338 26344
rect 42394 26288 42399 26344
rect 41045 26286 42399 26288
rect 41045 26283 41111 26286
rect 42333 26283 42399 26286
rect 42885 26346 42951 26349
rect 46657 26346 46723 26349
rect 42885 26344 46723 26346
rect 42885 26288 42890 26344
rect 42946 26288 46662 26344
rect 46718 26288 46723 26344
rect 42885 26286 46723 26288
rect 42885 26283 42951 26286
rect 46657 26283 46723 26286
rect 72509 26346 72575 26349
rect 74349 26346 74415 26349
rect 72509 26344 74415 26346
rect 72509 26288 72514 26344
rect 72570 26288 74354 26344
rect 74410 26288 74415 26344
rect 72509 26286 74415 26288
rect 72509 26283 72575 26286
rect 74349 26283 74415 26286
rect 86125 26346 86191 26349
rect 88241 26346 88307 26349
rect 86125 26344 88307 26346
rect 86125 26288 86130 26344
rect 86186 26288 88246 26344
rect 88302 26288 88307 26344
rect 86125 26286 88307 26288
rect 86125 26283 86191 26286
rect 88241 26283 88307 26286
rect 40953 26210 41019 26213
rect 48037 26210 48103 26213
rect 40953 26208 48103 26210
rect 40953 26152 40958 26208
rect 41014 26152 48042 26208
rect 48098 26152 48103 26208
rect 40953 26150 48103 26152
rect 40953 26147 41019 26150
rect 48037 26147 48103 26150
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 65648 26144 65968 26145
rect 65648 26080 65656 26144
rect 65720 26080 65736 26144
rect 65800 26080 65816 26144
rect 65880 26080 65896 26144
rect 65960 26080 65968 26144
rect 65648 26079 65968 26080
rect 96368 26144 96688 26145
rect 96368 26080 96376 26144
rect 96440 26080 96456 26144
rect 96520 26080 96536 26144
rect 96600 26080 96616 26144
rect 96680 26080 96688 26144
rect 96368 26079 96688 26080
rect 39849 25938 39915 25941
rect 54569 25938 54635 25941
rect 39849 25936 54635 25938
rect 39849 25880 39854 25936
rect 39910 25880 54574 25936
rect 54630 25880 54635 25936
rect 39849 25878 54635 25880
rect 39849 25875 39915 25878
rect 54569 25875 54635 25878
rect 35801 25802 35867 25805
rect 69289 25802 69355 25805
rect 35801 25800 69355 25802
rect 35801 25744 35806 25800
rect 35862 25744 69294 25800
rect 69350 25744 69355 25800
rect 35801 25742 69355 25744
rect 35801 25739 35867 25742
rect 69289 25739 69355 25742
rect 43253 25666 43319 25669
rect 43713 25666 43779 25669
rect 43253 25664 43779 25666
rect 43253 25608 43258 25664
rect 43314 25608 43718 25664
rect 43774 25608 43779 25664
rect 43253 25606 43779 25608
rect 43253 25603 43319 25606
rect 43713 25603 43779 25606
rect 50981 25666 51047 25669
rect 56225 25666 56291 25669
rect 50981 25664 56291 25666
rect 50981 25608 50986 25664
rect 51042 25608 56230 25664
rect 56286 25608 56291 25664
rect 50981 25606 56291 25608
rect 50981 25603 51047 25606
rect 56225 25603 56291 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 50288 25600 50608 25601
rect 50288 25536 50296 25600
rect 50360 25536 50376 25600
rect 50440 25536 50456 25600
rect 50520 25536 50536 25600
rect 50600 25536 50608 25600
rect 50288 25535 50608 25536
rect 81008 25600 81328 25601
rect 81008 25536 81016 25600
rect 81080 25536 81096 25600
rect 81160 25536 81176 25600
rect 81240 25536 81256 25600
rect 81320 25536 81328 25600
rect 81008 25535 81328 25536
rect 40493 25530 40559 25533
rect 41505 25530 41571 25533
rect 40493 25528 41571 25530
rect 40493 25472 40498 25528
rect 40554 25472 41510 25528
rect 41566 25472 41571 25528
rect 40493 25470 41571 25472
rect 40493 25467 40559 25470
rect 41505 25467 41571 25470
rect 52085 25530 52151 25533
rect 53649 25530 53715 25533
rect 52085 25528 53715 25530
rect 52085 25472 52090 25528
rect 52146 25472 53654 25528
rect 53710 25472 53715 25528
rect 52085 25470 53715 25472
rect 52085 25467 52151 25470
rect 53649 25467 53715 25470
rect 43621 25394 43687 25397
rect 74165 25394 74231 25397
rect 22050 25392 74231 25394
rect 22050 25336 43626 25392
rect 43682 25336 74170 25392
rect 74226 25336 74231 25392
rect 22050 25334 74231 25336
rect 13813 25258 13879 25261
rect 14273 25258 14339 25261
rect 22050 25258 22110 25334
rect 43621 25331 43687 25334
rect 74165 25331 74231 25334
rect 13813 25256 22110 25258
rect 13813 25200 13818 25256
rect 13874 25200 14278 25256
rect 14334 25200 22110 25256
rect 13813 25198 22110 25200
rect 41413 25258 41479 25261
rect 43713 25258 43779 25261
rect 41413 25256 43779 25258
rect 41413 25200 41418 25256
rect 41474 25200 43718 25256
rect 43774 25200 43779 25256
rect 41413 25198 43779 25200
rect 13813 25195 13879 25198
rect 14273 25195 14339 25198
rect 41413 25195 41479 25198
rect 43713 25195 43779 25198
rect 51257 25258 51323 25261
rect 56869 25258 56935 25261
rect 51257 25256 56935 25258
rect 51257 25200 51262 25256
rect 51318 25200 56874 25256
rect 56930 25200 56935 25256
rect 51257 25198 56935 25200
rect 51257 25195 51323 25198
rect 56869 25195 56935 25198
rect 62021 25258 62087 25261
rect 65609 25258 65675 25261
rect 62021 25256 65675 25258
rect 62021 25200 62026 25256
rect 62082 25200 65614 25256
rect 65670 25200 65675 25256
rect 62021 25198 65675 25200
rect 62021 25195 62087 25198
rect 65609 25195 65675 25198
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 65648 25056 65968 25057
rect 65648 24992 65656 25056
rect 65720 24992 65736 25056
rect 65800 24992 65816 25056
rect 65880 24992 65896 25056
rect 65960 24992 65968 25056
rect 65648 24991 65968 24992
rect 96368 25056 96688 25057
rect 96368 24992 96376 25056
rect 96440 24992 96456 25056
rect 96520 24992 96536 25056
rect 96600 24992 96616 25056
rect 96680 24992 96688 25056
rect 96368 24991 96688 24992
rect 43437 24850 43503 24853
rect 44633 24850 44699 24853
rect 43437 24848 44699 24850
rect 43437 24792 43442 24848
rect 43498 24792 44638 24848
rect 44694 24792 44699 24848
rect 43437 24790 44699 24792
rect 43437 24787 43503 24790
rect 44633 24787 44699 24790
rect 50521 24850 50587 24853
rect 51349 24850 51415 24853
rect 50521 24848 51415 24850
rect 50521 24792 50526 24848
rect 50582 24792 51354 24848
rect 51410 24792 51415 24848
rect 50521 24790 51415 24792
rect 50521 24787 50587 24790
rect 51349 24787 51415 24790
rect 40493 24714 40559 24717
rect 47025 24714 47091 24717
rect 40493 24712 47091 24714
rect 40493 24656 40498 24712
rect 40554 24656 47030 24712
rect 47086 24656 47091 24712
rect 40493 24654 47091 24656
rect 40493 24651 40559 24654
rect 47025 24651 47091 24654
rect 50521 24714 50587 24717
rect 51533 24714 51599 24717
rect 50521 24712 51599 24714
rect 50521 24656 50526 24712
rect 50582 24656 51538 24712
rect 51594 24656 51599 24712
rect 50521 24654 51599 24656
rect 50521 24651 50587 24654
rect 51533 24651 51599 24654
rect 30373 24578 30439 24581
rect 36997 24578 37063 24581
rect 30373 24576 37063 24578
rect 30373 24520 30378 24576
rect 30434 24520 37002 24576
rect 37058 24520 37063 24576
rect 30373 24518 37063 24520
rect 30373 24515 30439 24518
rect 36997 24515 37063 24518
rect 43529 24578 43595 24581
rect 46933 24578 46999 24581
rect 43529 24576 46999 24578
rect 43529 24520 43534 24576
rect 43590 24520 46938 24576
rect 46994 24520 46999 24576
rect 43529 24518 46999 24520
rect 43529 24515 43595 24518
rect 46933 24515 46999 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 50288 24512 50608 24513
rect 50288 24448 50296 24512
rect 50360 24448 50376 24512
rect 50440 24448 50456 24512
rect 50520 24448 50536 24512
rect 50600 24448 50608 24512
rect 50288 24447 50608 24448
rect 81008 24512 81328 24513
rect 81008 24448 81016 24512
rect 81080 24448 81096 24512
rect 81160 24448 81176 24512
rect 81240 24448 81256 24512
rect 81320 24448 81328 24512
rect 81008 24447 81328 24448
rect 41781 24442 41847 24445
rect 46657 24442 46723 24445
rect 46841 24442 46907 24445
rect 41781 24440 46723 24442
rect 41781 24384 41786 24440
rect 41842 24384 46662 24440
rect 46718 24384 46723 24440
rect 41781 24382 46723 24384
rect 41781 24379 41847 24382
rect 46657 24379 46723 24382
rect 46798 24440 46907 24442
rect 46798 24384 46846 24440
rect 46902 24384 46907 24440
rect 46798 24379 46907 24384
rect 75085 24442 75151 24445
rect 76373 24442 76439 24445
rect 75085 24440 76439 24442
rect 75085 24384 75090 24440
rect 75146 24384 76378 24440
rect 76434 24384 76439 24440
rect 75085 24382 76439 24384
rect 75085 24379 75151 24382
rect 76373 24379 76439 24382
rect 46657 24170 46723 24173
rect 46798 24170 46858 24379
rect 75729 24306 75795 24309
rect 76281 24306 76347 24309
rect 75729 24304 76347 24306
rect 75729 24248 75734 24304
rect 75790 24248 76286 24304
rect 76342 24248 76347 24304
rect 75729 24246 76347 24248
rect 75729 24243 75795 24246
rect 76281 24243 76347 24246
rect 46657 24168 46858 24170
rect 46657 24112 46662 24168
rect 46718 24112 46858 24168
rect 46657 24110 46858 24112
rect 74717 24170 74783 24173
rect 78489 24170 78555 24173
rect 74717 24168 78555 24170
rect 74717 24112 74722 24168
rect 74778 24112 78494 24168
rect 78550 24112 78555 24168
rect 74717 24110 78555 24112
rect 46657 24107 46723 24110
rect 74717 24107 74783 24110
rect 78489 24107 78555 24110
rect 40953 24034 41019 24037
rect 46933 24034 46999 24037
rect 40953 24032 46999 24034
rect 40953 23976 40958 24032
rect 41014 23976 46938 24032
rect 46994 23976 46999 24032
rect 40953 23974 46999 23976
rect 40953 23971 41019 23974
rect 46933 23971 46999 23974
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 65648 23968 65968 23969
rect 65648 23904 65656 23968
rect 65720 23904 65736 23968
rect 65800 23904 65816 23968
rect 65880 23904 65896 23968
rect 65960 23904 65968 23968
rect 65648 23903 65968 23904
rect 96368 23968 96688 23969
rect 96368 23904 96376 23968
rect 96440 23904 96456 23968
rect 96520 23904 96536 23968
rect 96600 23904 96616 23968
rect 96680 23904 96688 23968
rect 96368 23903 96688 23904
rect 42977 23762 43043 23765
rect 45369 23762 45435 23765
rect 42977 23760 45435 23762
rect 42977 23704 42982 23760
rect 43038 23704 45374 23760
rect 45430 23704 45435 23760
rect 42977 23702 45435 23704
rect 42977 23699 43043 23702
rect 45369 23699 45435 23702
rect 71865 23762 71931 23765
rect 76281 23762 76347 23765
rect 71865 23760 76347 23762
rect 71865 23704 71870 23760
rect 71926 23704 76286 23760
rect 76342 23704 76347 23760
rect 71865 23702 76347 23704
rect 71865 23699 71931 23702
rect 76281 23699 76347 23702
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 50288 23424 50608 23425
rect 50288 23360 50296 23424
rect 50360 23360 50376 23424
rect 50440 23360 50456 23424
rect 50520 23360 50536 23424
rect 50600 23360 50608 23424
rect 50288 23359 50608 23360
rect 81008 23424 81328 23425
rect 81008 23360 81016 23424
rect 81080 23360 81096 23424
rect 81160 23360 81176 23424
rect 81240 23360 81256 23424
rect 81320 23360 81328 23424
rect 81008 23359 81328 23360
rect 26509 23354 26575 23357
rect 26374 23352 26575 23354
rect 26374 23296 26514 23352
rect 26570 23296 26575 23352
rect 26374 23294 26575 23296
rect 26374 23085 26434 23294
rect 26509 23291 26575 23294
rect 51165 23218 51231 23221
rect 55029 23218 55095 23221
rect 51165 23216 55095 23218
rect 51165 23160 51170 23216
rect 51226 23160 55034 23216
rect 55090 23160 55095 23216
rect 51165 23158 55095 23160
rect 51165 23155 51231 23158
rect 55029 23155 55095 23158
rect 26325 23080 26434 23085
rect 26877 23082 26943 23085
rect 26325 23024 26330 23080
rect 26386 23024 26434 23080
rect 26325 23022 26434 23024
rect 26558 23080 26943 23082
rect 26558 23024 26882 23080
rect 26938 23024 26943 23080
rect 26558 23022 26943 23024
rect 26325 23019 26391 23022
rect 25313 22946 25379 22949
rect 26558 22946 26618 23022
rect 26877 23019 26943 23022
rect 47301 23082 47367 23085
rect 48037 23082 48103 23085
rect 47301 23080 48103 23082
rect 47301 23024 47306 23080
rect 47362 23024 48042 23080
rect 48098 23024 48103 23080
rect 47301 23022 48103 23024
rect 47301 23019 47367 23022
rect 48037 23019 48103 23022
rect 61469 23082 61535 23085
rect 65885 23082 65951 23085
rect 61469 23080 65951 23082
rect 61469 23024 61474 23080
rect 61530 23024 65890 23080
rect 65946 23024 65951 23080
rect 61469 23022 65951 23024
rect 61469 23019 61535 23022
rect 65885 23019 65951 23022
rect 25313 22944 26618 22946
rect 25313 22888 25318 22944
rect 25374 22888 26618 22944
rect 25313 22886 26618 22888
rect 25313 22883 25379 22886
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 65648 22880 65968 22881
rect 65648 22816 65656 22880
rect 65720 22816 65736 22880
rect 65800 22816 65816 22880
rect 65880 22816 65896 22880
rect 65960 22816 65968 22880
rect 65648 22815 65968 22816
rect 96368 22880 96688 22881
rect 96368 22816 96376 22880
rect 96440 22816 96456 22880
rect 96520 22816 96536 22880
rect 96600 22816 96616 22880
rect 96680 22816 96688 22880
rect 96368 22815 96688 22816
rect 64965 22810 65031 22813
rect 64965 22808 65258 22810
rect 64965 22752 64970 22808
rect 65026 22752 65258 22808
rect 64965 22750 65258 22752
rect 64965 22747 65031 22750
rect 33593 22674 33659 22677
rect 33869 22674 33935 22677
rect 33593 22672 33935 22674
rect 33593 22616 33598 22672
rect 33654 22616 33874 22672
rect 33930 22616 33935 22672
rect 33593 22614 33935 22616
rect 33593 22611 33659 22614
rect 33869 22611 33935 22614
rect 61009 22538 61075 22541
rect 62205 22538 62271 22541
rect 65057 22538 65123 22541
rect 61009 22536 65123 22538
rect 61009 22480 61014 22536
rect 61070 22480 62210 22536
rect 62266 22480 65062 22536
rect 65118 22480 65123 22536
rect 61009 22478 65123 22480
rect 61009 22475 61075 22478
rect 62205 22475 62271 22478
rect 65057 22475 65123 22478
rect 65198 22405 65258 22750
rect 33961 22402 34027 22405
rect 38561 22402 38627 22405
rect 33961 22400 38627 22402
rect 33961 22344 33966 22400
rect 34022 22344 38566 22400
rect 38622 22344 38627 22400
rect 33961 22342 38627 22344
rect 65198 22400 65307 22405
rect 65198 22344 65246 22400
rect 65302 22344 65307 22400
rect 65198 22342 65307 22344
rect 33961 22339 34027 22342
rect 38561 22339 38627 22342
rect 65241 22339 65307 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 50288 22336 50608 22337
rect 50288 22272 50296 22336
rect 50360 22272 50376 22336
rect 50440 22272 50456 22336
rect 50520 22272 50536 22336
rect 50600 22272 50608 22336
rect 50288 22271 50608 22272
rect 81008 22336 81328 22337
rect 81008 22272 81016 22336
rect 81080 22272 81096 22336
rect 81160 22272 81176 22336
rect 81240 22272 81256 22336
rect 81320 22272 81328 22336
rect 81008 22271 81328 22272
rect 32489 22266 32555 22269
rect 38469 22266 38535 22269
rect 32489 22264 38535 22266
rect 32489 22208 32494 22264
rect 32550 22208 38474 22264
rect 38530 22208 38535 22264
rect 32489 22206 38535 22208
rect 32489 22203 32555 22206
rect 38469 22203 38535 22206
rect 33041 22130 33107 22133
rect 37641 22130 37707 22133
rect 33041 22128 37707 22130
rect 33041 22072 33046 22128
rect 33102 22072 37646 22128
rect 37702 22072 37707 22128
rect 33041 22070 37707 22072
rect 33041 22067 33107 22070
rect 37641 22067 37707 22070
rect 9949 21994 10015 21997
rect 85297 21994 85363 21997
rect 9949 21992 85363 21994
rect 9949 21936 9954 21992
rect 10010 21936 85302 21992
rect 85358 21936 85363 21992
rect 9949 21934 85363 21936
rect 9949 21931 10015 21934
rect 85297 21931 85363 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 65648 21792 65968 21793
rect 65648 21728 65656 21792
rect 65720 21728 65736 21792
rect 65800 21728 65816 21792
rect 65880 21728 65896 21792
rect 65960 21728 65968 21792
rect 65648 21727 65968 21728
rect 96368 21792 96688 21793
rect 96368 21728 96376 21792
rect 96440 21728 96456 21792
rect 96520 21728 96536 21792
rect 96600 21728 96616 21792
rect 96680 21728 96688 21792
rect 96368 21727 96688 21728
rect 60825 21722 60891 21725
rect 61101 21722 61167 21725
rect 60825 21720 61167 21722
rect 60825 21664 60830 21720
rect 60886 21664 61106 21720
rect 61162 21664 61167 21720
rect 60825 21662 61167 21664
rect 60825 21659 60891 21662
rect 61101 21659 61167 21662
rect 37825 21586 37891 21589
rect 38561 21588 38627 21589
rect 38510 21586 38516 21588
rect 37825 21584 38516 21586
rect 38580 21584 38627 21588
rect 37825 21528 37830 21584
rect 37886 21528 38516 21584
rect 38622 21528 38627 21584
rect 37825 21526 38516 21528
rect 37825 21523 37891 21526
rect 38510 21524 38516 21526
rect 38580 21524 38627 21528
rect 38561 21523 38627 21524
rect 50889 21586 50955 21589
rect 55029 21586 55095 21589
rect 50889 21584 55095 21586
rect 50889 21528 50894 21584
rect 50950 21528 55034 21584
rect 55090 21528 55095 21584
rect 50889 21526 55095 21528
rect 50889 21523 50955 21526
rect 55029 21523 55095 21526
rect 65517 21586 65583 21589
rect 66161 21586 66227 21589
rect 65517 21584 66227 21586
rect 65517 21528 65522 21584
rect 65578 21528 66166 21584
rect 66222 21528 66227 21584
rect 65517 21526 66227 21528
rect 65517 21523 65583 21526
rect 66161 21523 66227 21526
rect 41505 21450 41571 21453
rect 44541 21450 44607 21453
rect 41505 21448 44607 21450
rect 41505 21392 41510 21448
rect 41566 21392 44546 21448
rect 44602 21392 44607 21448
rect 41505 21390 44607 21392
rect 41505 21387 41571 21390
rect 44541 21387 44607 21390
rect 61285 21450 61351 21453
rect 61561 21450 61627 21453
rect 61285 21448 61627 21450
rect 61285 21392 61290 21448
rect 61346 21392 61566 21448
rect 61622 21392 61627 21448
rect 61285 21390 61627 21392
rect 61285 21387 61351 21390
rect 61561 21387 61627 21390
rect 61561 21314 61627 21317
rect 63585 21314 63651 21317
rect 61561 21312 63651 21314
rect 61561 21256 61566 21312
rect 61622 21256 63590 21312
rect 63646 21256 63651 21312
rect 61561 21254 63651 21256
rect 61561 21251 61627 21254
rect 63585 21251 63651 21254
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 50288 21248 50608 21249
rect 50288 21184 50296 21248
rect 50360 21184 50376 21248
rect 50440 21184 50456 21248
rect 50520 21184 50536 21248
rect 50600 21184 50608 21248
rect 50288 21183 50608 21184
rect 81008 21248 81328 21249
rect 81008 21184 81016 21248
rect 81080 21184 81096 21248
rect 81160 21184 81176 21248
rect 81240 21184 81256 21248
rect 81320 21184 81328 21248
rect 81008 21183 81328 21184
rect 50889 20906 50955 20909
rect 51165 20906 51231 20909
rect 50889 20904 51231 20906
rect 50889 20848 50894 20904
rect 50950 20848 51170 20904
rect 51226 20848 51231 20904
rect 50889 20846 51231 20848
rect 50889 20843 50955 20846
rect 51165 20843 51231 20846
rect 60549 20906 60615 20909
rect 67357 20906 67423 20909
rect 60549 20904 67423 20906
rect 60549 20848 60554 20904
rect 60610 20848 67362 20904
rect 67418 20848 67423 20904
rect 60549 20846 67423 20848
rect 60549 20843 60615 20846
rect 67357 20843 67423 20846
rect 53741 20770 53807 20773
rect 55857 20770 55923 20773
rect 53741 20768 55923 20770
rect 53741 20712 53746 20768
rect 53802 20712 55862 20768
rect 55918 20712 55923 20768
rect 53741 20710 55923 20712
rect 53741 20707 53807 20710
rect 55857 20707 55923 20710
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 65648 20704 65968 20705
rect 65648 20640 65656 20704
rect 65720 20640 65736 20704
rect 65800 20640 65816 20704
rect 65880 20640 65896 20704
rect 65960 20640 65968 20704
rect 65648 20639 65968 20640
rect 96368 20704 96688 20705
rect 96368 20640 96376 20704
rect 96440 20640 96456 20704
rect 96520 20640 96536 20704
rect 96600 20640 96616 20704
rect 96680 20640 96688 20704
rect 96368 20639 96688 20640
rect 22461 20634 22527 20637
rect 23013 20634 23079 20637
rect 22461 20632 23079 20634
rect 22461 20576 22466 20632
rect 22522 20576 23018 20632
rect 23074 20576 23079 20632
rect 22461 20574 23079 20576
rect 22461 20571 22527 20574
rect 23013 20571 23079 20574
rect 54477 20634 54543 20637
rect 54753 20634 54819 20637
rect 58617 20634 58683 20637
rect 54477 20632 58683 20634
rect 54477 20576 54482 20632
rect 54538 20576 54758 20632
rect 54814 20576 58622 20632
rect 58678 20576 58683 20632
rect 54477 20574 58683 20576
rect 54477 20571 54543 20574
rect 54753 20571 54819 20574
rect 58617 20571 58683 20574
rect 62941 20634 63007 20637
rect 64781 20634 64847 20637
rect 62941 20632 64847 20634
rect 62941 20576 62946 20632
rect 63002 20576 64786 20632
rect 64842 20576 64847 20632
rect 62941 20574 64847 20576
rect 62941 20571 63007 20574
rect 64781 20571 64847 20574
rect 22461 20498 22527 20501
rect 23013 20498 23079 20501
rect 22461 20496 23079 20498
rect 22461 20440 22466 20496
rect 22522 20440 23018 20496
rect 23074 20440 23079 20496
rect 22461 20438 23079 20440
rect 22461 20435 22527 20438
rect 23013 20435 23079 20438
rect 64505 20498 64571 20501
rect 65977 20498 66043 20501
rect 64505 20496 66043 20498
rect 64505 20440 64510 20496
rect 64566 20440 65982 20496
rect 66038 20440 66043 20496
rect 64505 20438 66043 20440
rect 64505 20435 64571 20438
rect 65977 20435 66043 20438
rect 80973 20498 81039 20501
rect 82261 20498 82327 20501
rect 80973 20496 82327 20498
rect 80973 20440 80978 20496
rect 81034 20440 82266 20496
rect 82322 20440 82327 20496
rect 80973 20438 82327 20440
rect 80973 20435 81039 20438
rect 82261 20435 82327 20438
rect 33685 20362 33751 20365
rect 34697 20362 34763 20365
rect 33685 20360 34763 20362
rect 33685 20304 33690 20360
rect 33746 20304 34702 20360
rect 34758 20304 34763 20360
rect 33685 20302 34763 20304
rect 33685 20299 33751 20302
rect 34697 20299 34763 20302
rect 48313 20362 48379 20365
rect 56133 20362 56199 20365
rect 48313 20360 56199 20362
rect 48313 20304 48318 20360
rect 48374 20304 56138 20360
rect 56194 20304 56199 20360
rect 48313 20302 56199 20304
rect 48313 20299 48379 20302
rect 56133 20299 56199 20302
rect 64045 20362 64111 20365
rect 65241 20362 65307 20365
rect 64045 20360 65307 20362
rect 64045 20304 64050 20360
rect 64106 20304 65246 20360
rect 65302 20304 65307 20360
rect 64045 20302 65307 20304
rect 64045 20299 64111 20302
rect 65241 20299 65307 20302
rect 79041 20362 79107 20365
rect 82169 20362 82235 20365
rect 79041 20360 82235 20362
rect 79041 20304 79046 20360
rect 79102 20304 82174 20360
rect 82230 20304 82235 20360
rect 79041 20302 82235 20304
rect 79041 20299 79107 20302
rect 82169 20299 82235 20302
rect 19568 20160 19888 20161
rect 0 20090 800 20120
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 50288 20160 50608 20161
rect 50288 20096 50296 20160
rect 50360 20096 50376 20160
rect 50440 20096 50456 20160
rect 50520 20096 50536 20160
rect 50600 20096 50608 20160
rect 50288 20095 50608 20096
rect 81008 20160 81328 20161
rect 81008 20096 81016 20160
rect 81080 20096 81096 20160
rect 81160 20096 81176 20160
rect 81240 20096 81256 20160
rect 81320 20096 81328 20160
rect 81008 20095 81328 20096
rect 1393 20090 1459 20093
rect 0 20088 1459 20090
rect 0 20032 1398 20088
rect 1454 20032 1459 20088
rect 0 20030 1459 20032
rect 0 20000 800 20030
rect 1393 20027 1459 20030
rect 33685 20090 33751 20093
rect 38561 20090 38627 20093
rect 33685 20088 38627 20090
rect 33685 20032 33690 20088
rect 33746 20032 38566 20088
rect 38622 20032 38627 20088
rect 33685 20030 38627 20032
rect 33685 20027 33751 20030
rect 38561 20027 38627 20030
rect 97625 20090 97691 20093
rect 99200 20090 100000 20120
rect 97625 20088 100000 20090
rect 97625 20032 97630 20088
rect 97686 20032 100000 20088
rect 97625 20030 100000 20032
rect 97625 20027 97691 20030
rect 99200 20000 100000 20030
rect 34053 19954 34119 19957
rect 37733 19954 37799 19957
rect 34053 19952 37799 19954
rect 34053 19896 34058 19952
rect 34114 19896 37738 19952
rect 37794 19896 37799 19952
rect 34053 19894 37799 19896
rect 34053 19891 34119 19894
rect 37733 19891 37799 19894
rect 48313 19954 48379 19957
rect 53097 19954 53163 19957
rect 48313 19952 53163 19954
rect 48313 19896 48318 19952
rect 48374 19896 53102 19952
rect 53158 19896 53163 19952
rect 48313 19894 53163 19896
rect 48313 19891 48379 19894
rect 53097 19891 53163 19894
rect 38653 19818 38719 19821
rect 39113 19818 39179 19821
rect 43989 19818 44055 19821
rect 38653 19816 44055 19818
rect 38653 19760 38658 19816
rect 38714 19760 39118 19816
rect 39174 19760 43994 19816
rect 44050 19760 44055 19816
rect 38653 19758 44055 19760
rect 38653 19755 38719 19758
rect 39113 19755 39179 19758
rect 43989 19755 44055 19758
rect 38745 19682 38811 19685
rect 43437 19682 43503 19685
rect 38745 19680 43503 19682
rect 38745 19624 38750 19680
rect 38806 19624 43442 19680
rect 43498 19624 43503 19680
rect 38745 19622 43503 19624
rect 38745 19619 38811 19622
rect 43437 19619 43503 19622
rect 43897 19682 43963 19685
rect 45921 19682 45987 19685
rect 43897 19680 45987 19682
rect 43897 19624 43902 19680
rect 43958 19624 45926 19680
rect 45982 19624 45987 19680
rect 43897 19622 45987 19624
rect 43897 19619 43963 19622
rect 45921 19619 45987 19622
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 65648 19616 65968 19617
rect 65648 19552 65656 19616
rect 65720 19552 65736 19616
rect 65800 19552 65816 19616
rect 65880 19552 65896 19616
rect 65960 19552 65968 19616
rect 65648 19551 65968 19552
rect 96368 19616 96688 19617
rect 96368 19552 96376 19616
rect 96440 19552 96456 19616
rect 96520 19552 96536 19616
rect 96600 19552 96616 19616
rect 96680 19552 96688 19616
rect 96368 19551 96688 19552
rect 44081 19546 44147 19549
rect 44817 19546 44883 19549
rect 46933 19546 46999 19549
rect 44081 19544 46999 19546
rect 44081 19488 44086 19544
rect 44142 19488 44822 19544
rect 44878 19488 46938 19544
rect 46994 19488 46999 19544
rect 44081 19486 46999 19488
rect 44081 19483 44147 19486
rect 44817 19483 44883 19486
rect 46933 19483 46999 19486
rect 60733 19546 60799 19549
rect 61101 19546 61167 19549
rect 60733 19544 61167 19546
rect 60733 19488 60738 19544
rect 60794 19488 61106 19544
rect 61162 19488 61167 19544
rect 60733 19486 61167 19488
rect 60733 19483 60799 19486
rect 61101 19483 61167 19486
rect 33685 19410 33751 19413
rect 36629 19410 36695 19413
rect 33685 19408 36695 19410
rect 33685 19352 33690 19408
rect 33746 19352 36634 19408
rect 36690 19352 36695 19408
rect 33685 19350 36695 19352
rect 33685 19347 33751 19350
rect 36629 19347 36695 19350
rect 45093 19410 45159 19413
rect 46105 19410 46171 19413
rect 45093 19408 46171 19410
rect 45093 19352 45098 19408
rect 45154 19352 46110 19408
rect 46166 19352 46171 19408
rect 45093 19350 46171 19352
rect 45093 19347 45159 19350
rect 46105 19347 46171 19350
rect 21633 19274 21699 19277
rect 22737 19274 22803 19277
rect 21633 19272 22803 19274
rect 21633 19216 21638 19272
rect 21694 19216 22742 19272
rect 22798 19216 22803 19272
rect 21633 19214 22803 19216
rect 21633 19211 21699 19214
rect 22737 19211 22803 19214
rect 36077 19274 36143 19277
rect 36721 19274 36787 19277
rect 52637 19274 52703 19277
rect 36077 19272 36787 19274
rect 36077 19216 36082 19272
rect 36138 19216 36726 19272
rect 36782 19216 36787 19272
rect 36077 19214 36787 19216
rect 36077 19211 36143 19214
rect 36721 19211 36787 19214
rect 41370 19272 52703 19274
rect 41370 19216 52642 19272
rect 52698 19216 52703 19272
rect 41370 19214 52703 19216
rect 22461 19138 22527 19141
rect 23013 19138 23079 19141
rect 22461 19136 23079 19138
rect 22461 19080 22466 19136
rect 22522 19080 23018 19136
rect 23074 19080 23079 19136
rect 22461 19078 23079 19080
rect 22461 19075 22527 19078
rect 23013 19075 23079 19078
rect 25037 19138 25103 19141
rect 34421 19138 34487 19141
rect 25037 19136 34487 19138
rect 25037 19080 25042 19136
rect 25098 19080 34426 19136
rect 34482 19080 34487 19136
rect 25037 19078 34487 19080
rect 25037 19075 25103 19078
rect 34421 19075 34487 19078
rect 34697 19138 34763 19141
rect 36721 19138 36787 19141
rect 34697 19136 36787 19138
rect 34697 19080 34702 19136
rect 34758 19080 36726 19136
rect 36782 19080 36787 19136
rect 34697 19078 36787 19080
rect 34697 19075 34763 19078
rect 36721 19075 36787 19078
rect 38193 19138 38259 19141
rect 41370 19138 41430 19214
rect 52637 19211 52703 19214
rect 60733 19274 60799 19277
rect 61101 19274 61167 19277
rect 60733 19272 61167 19274
rect 60733 19216 60738 19272
rect 60794 19216 61106 19272
rect 61162 19216 61167 19272
rect 60733 19214 61167 19216
rect 60733 19211 60799 19214
rect 61101 19211 61167 19214
rect 38193 19136 41430 19138
rect 38193 19080 38198 19136
rect 38254 19080 41430 19136
rect 38193 19078 41430 19080
rect 43437 19138 43503 19141
rect 47117 19138 47183 19141
rect 43437 19136 47183 19138
rect 43437 19080 43442 19136
rect 43498 19080 47122 19136
rect 47178 19080 47183 19136
rect 43437 19078 47183 19080
rect 38193 19075 38259 19078
rect 43437 19075 43503 19078
rect 47117 19075 47183 19078
rect 59353 19138 59419 19141
rect 60825 19138 60891 19141
rect 59353 19136 60891 19138
rect 59353 19080 59358 19136
rect 59414 19080 60830 19136
rect 60886 19080 60891 19136
rect 59353 19078 60891 19080
rect 59353 19075 59419 19078
rect 60825 19075 60891 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 50288 19072 50608 19073
rect 50288 19008 50296 19072
rect 50360 19008 50376 19072
rect 50440 19008 50456 19072
rect 50520 19008 50536 19072
rect 50600 19008 50608 19072
rect 50288 19007 50608 19008
rect 81008 19072 81328 19073
rect 81008 19008 81016 19072
rect 81080 19008 81096 19072
rect 81160 19008 81176 19072
rect 81240 19008 81256 19072
rect 81320 19008 81328 19072
rect 81008 19007 81328 19008
rect 34237 19002 34303 19005
rect 39849 19002 39915 19005
rect 34237 19000 39915 19002
rect 34237 18944 34242 19000
rect 34298 18944 39854 19000
rect 39910 18944 39915 19000
rect 34237 18942 39915 18944
rect 34237 18939 34303 18942
rect 39849 18939 39915 18942
rect 40033 19002 40099 19005
rect 43161 19002 43227 19005
rect 40033 19000 43227 19002
rect 40033 18944 40038 19000
rect 40094 18944 43166 19000
rect 43222 18944 43227 19000
rect 40033 18942 43227 18944
rect 40033 18939 40099 18942
rect 43161 18939 43227 18942
rect 44633 19002 44699 19005
rect 46289 19002 46355 19005
rect 44633 19000 46355 19002
rect 44633 18944 44638 19000
rect 44694 18944 46294 19000
rect 46350 18944 46355 19000
rect 44633 18942 46355 18944
rect 44633 18939 44699 18942
rect 46289 18939 46355 18942
rect 33593 18866 33659 18869
rect 38510 18866 38516 18868
rect 33593 18864 38516 18866
rect 33593 18808 33598 18864
rect 33654 18808 38516 18864
rect 33593 18806 38516 18808
rect 33593 18803 33659 18806
rect 38510 18804 38516 18806
rect 38580 18866 38586 18868
rect 46105 18866 46171 18869
rect 38580 18864 46171 18866
rect 38580 18808 46110 18864
rect 46166 18808 46171 18864
rect 38580 18806 46171 18808
rect 38580 18804 38586 18806
rect 46105 18803 46171 18806
rect 50705 18866 50771 18869
rect 51165 18866 51231 18869
rect 50705 18864 51231 18866
rect 50705 18808 50710 18864
rect 50766 18808 51170 18864
rect 51226 18808 51231 18864
rect 50705 18806 51231 18808
rect 50705 18803 50771 18806
rect 51165 18803 51231 18806
rect 51717 18866 51783 18869
rect 55765 18866 55831 18869
rect 51717 18864 55831 18866
rect 51717 18808 51722 18864
rect 51778 18808 55770 18864
rect 55826 18808 55831 18864
rect 51717 18806 55831 18808
rect 51717 18803 51783 18806
rect 55765 18803 55831 18806
rect 69289 18866 69355 18869
rect 70209 18866 70275 18869
rect 69289 18864 70275 18866
rect 69289 18808 69294 18864
rect 69350 18808 70214 18864
rect 70270 18808 70275 18864
rect 69289 18806 70275 18808
rect 69289 18803 69355 18806
rect 70209 18803 70275 18806
rect 70761 18866 70827 18869
rect 71129 18866 71195 18869
rect 70761 18864 71195 18866
rect 70761 18808 70766 18864
rect 70822 18808 71134 18864
rect 71190 18808 71195 18864
rect 70761 18806 71195 18808
rect 70761 18803 70827 18806
rect 71129 18803 71195 18806
rect 33409 18730 33475 18733
rect 36629 18730 36695 18733
rect 33409 18728 36695 18730
rect 33409 18672 33414 18728
rect 33470 18672 36634 18728
rect 36690 18672 36695 18728
rect 33409 18670 36695 18672
rect 33409 18667 33475 18670
rect 36629 18667 36695 18670
rect 40953 18730 41019 18733
rect 42793 18730 42859 18733
rect 40953 18728 42859 18730
rect 40953 18672 40958 18728
rect 41014 18672 42798 18728
rect 42854 18672 42859 18728
rect 40953 18670 42859 18672
rect 40953 18667 41019 18670
rect 42793 18667 42859 18670
rect 44725 18730 44791 18733
rect 50797 18730 50863 18733
rect 62205 18730 62271 18733
rect 72417 18730 72483 18733
rect 44725 18728 50863 18730
rect 44725 18672 44730 18728
rect 44786 18672 50802 18728
rect 50858 18672 50863 18728
rect 44725 18670 50863 18672
rect 44725 18667 44791 18670
rect 50797 18667 50863 18670
rect 60690 18728 72483 18730
rect 60690 18672 62210 18728
rect 62266 18672 72422 18728
rect 72478 18672 72483 18728
rect 60690 18670 72483 18672
rect 60690 18597 60750 18670
rect 62205 18667 62271 18670
rect 72417 18667 72483 18670
rect 20713 18594 20779 18597
rect 23013 18594 23079 18597
rect 20713 18592 23079 18594
rect 20713 18536 20718 18592
rect 20774 18536 23018 18592
rect 23074 18536 23079 18592
rect 20713 18534 23079 18536
rect 20713 18531 20779 18534
rect 23013 18531 23079 18534
rect 39757 18594 39823 18597
rect 44541 18594 44607 18597
rect 39757 18592 44607 18594
rect 39757 18536 39762 18592
rect 39818 18536 44546 18592
rect 44602 18536 44607 18592
rect 39757 18534 44607 18536
rect 39757 18531 39823 18534
rect 44541 18531 44607 18534
rect 48681 18594 48747 18597
rect 52269 18594 52335 18597
rect 48681 18592 52335 18594
rect 48681 18536 48686 18592
rect 48742 18536 52274 18592
rect 52330 18536 52335 18592
rect 48681 18534 52335 18536
rect 48681 18531 48747 18534
rect 52269 18531 52335 18534
rect 60641 18592 60750 18597
rect 60641 18536 60646 18592
rect 60702 18536 60750 18592
rect 60641 18534 60750 18536
rect 60641 18531 60707 18534
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 65648 18528 65968 18529
rect 65648 18464 65656 18528
rect 65720 18464 65736 18528
rect 65800 18464 65816 18528
rect 65880 18464 65896 18528
rect 65960 18464 65968 18528
rect 65648 18463 65968 18464
rect 96368 18528 96688 18529
rect 96368 18464 96376 18528
rect 96440 18464 96456 18528
rect 96520 18464 96536 18528
rect 96600 18464 96616 18528
rect 96680 18464 96688 18528
rect 96368 18463 96688 18464
rect 33501 18458 33567 18461
rect 34145 18458 34211 18461
rect 33501 18456 34211 18458
rect 33501 18400 33506 18456
rect 33562 18400 34150 18456
rect 34206 18400 34211 18456
rect 33501 18398 34211 18400
rect 33501 18395 33567 18398
rect 34145 18395 34211 18398
rect 41413 18458 41479 18461
rect 46933 18458 46999 18461
rect 41413 18456 46999 18458
rect 41413 18400 41418 18456
rect 41474 18400 46938 18456
rect 46994 18400 46999 18456
rect 41413 18398 46999 18400
rect 41413 18395 41479 18398
rect 46933 18395 46999 18398
rect 25221 18322 25287 18325
rect 33041 18322 33107 18325
rect 25221 18320 33107 18322
rect 25221 18264 25226 18320
rect 25282 18264 33046 18320
rect 33102 18264 33107 18320
rect 25221 18262 33107 18264
rect 25221 18259 25287 18262
rect 33041 18259 33107 18262
rect 33593 18322 33659 18325
rect 35157 18322 35223 18325
rect 33593 18320 35223 18322
rect 33593 18264 33598 18320
rect 33654 18264 35162 18320
rect 35218 18264 35223 18320
rect 33593 18262 35223 18264
rect 33593 18259 33659 18262
rect 35157 18259 35223 18262
rect 35341 18322 35407 18325
rect 43437 18322 43503 18325
rect 35341 18320 43503 18322
rect 35341 18264 35346 18320
rect 35402 18264 43442 18320
rect 43498 18264 43503 18320
rect 35341 18262 43503 18264
rect 35341 18259 35407 18262
rect 43437 18259 43503 18262
rect 60457 18322 60523 18325
rect 66253 18322 66319 18325
rect 60457 18320 66319 18322
rect 60457 18264 60462 18320
rect 60518 18264 66258 18320
rect 66314 18264 66319 18320
rect 60457 18262 66319 18264
rect 60457 18259 60523 18262
rect 66253 18259 66319 18262
rect 10869 18186 10935 18189
rect 96981 18186 97047 18189
rect 10869 18184 97047 18186
rect 10869 18128 10874 18184
rect 10930 18128 96986 18184
rect 97042 18128 97047 18184
rect 10869 18126 97047 18128
rect 10869 18123 10935 18126
rect 96981 18123 97047 18126
rect 29085 18050 29151 18053
rect 36721 18050 36787 18053
rect 29085 18048 36787 18050
rect 29085 17992 29090 18048
rect 29146 17992 36726 18048
rect 36782 17992 36787 18048
rect 29085 17990 36787 17992
rect 29085 17987 29151 17990
rect 36721 17987 36787 17990
rect 39297 18050 39363 18053
rect 41781 18050 41847 18053
rect 39297 18048 41847 18050
rect 39297 17992 39302 18048
rect 39358 17992 41786 18048
rect 41842 17992 41847 18048
rect 39297 17990 41847 17992
rect 39297 17987 39363 17990
rect 41781 17987 41847 17990
rect 46105 18050 46171 18053
rect 46381 18050 46447 18053
rect 46105 18048 46447 18050
rect 46105 17992 46110 18048
rect 46166 17992 46386 18048
rect 46442 17992 46447 18048
rect 46105 17990 46447 17992
rect 46105 17987 46171 17990
rect 46381 17987 46447 17990
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 50288 17984 50608 17985
rect 50288 17920 50296 17984
rect 50360 17920 50376 17984
rect 50440 17920 50456 17984
rect 50520 17920 50536 17984
rect 50600 17920 50608 17984
rect 50288 17919 50608 17920
rect 81008 17984 81328 17985
rect 81008 17920 81016 17984
rect 81080 17920 81096 17984
rect 81160 17920 81176 17984
rect 81240 17920 81256 17984
rect 81320 17920 81328 17984
rect 81008 17919 81328 17920
rect 21817 17914 21883 17917
rect 24669 17914 24735 17917
rect 29085 17914 29151 17917
rect 21817 17912 29151 17914
rect 21817 17856 21822 17912
rect 21878 17856 24674 17912
rect 24730 17856 29090 17912
rect 29146 17856 29151 17912
rect 21817 17854 29151 17856
rect 21817 17851 21883 17854
rect 24669 17851 24735 17854
rect 29085 17851 29151 17854
rect 38561 17914 38627 17917
rect 41413 17914 41479 17917
rect 38561 17912 41479 17914
rect 38561 17856 38566 17912
rect 38622 17856 41418 17912
rect 41474 17856 41479 17912
rect 38561 17854 41479 17856
rect 38561 17851 38627 17854
rect 41413 17851 41479 17854
rect 45461 17914 45527 17917
rect 46381 17914 46447 17917
rect 45461 17912 46447 17914
rect 45461 17856 45466 17912
rect 45522 17856 46386 17912
rect 46442 17856 46447 17912
rect 45461 17854 46447 17856
rect 45461 17851 45527 17854
rect 46381 17851 46447 17854
rect 2129 17778 2195 17781
rect 71957 17778 72023 17781
rect 2129 17776 72023 17778
rect 2129 17720 2134 17776
rect 2190 17720 71962 17776
rect 72018 17720 72023 17776
rect 2129 17718 72023 17720
rect 2129 17715 2195 17718
rect 71957 17715 72023 17718
rect 26877 17642 26943 17645
rect 28625 17642 28691 17645
rect 26877 17640 28691 17642
rect 26877 17584 26882 17640
rect 26938 17584 28630 17640
rect 28686 17584 28691 17640
rect 26877 17582 28691 17584
rect 26877 17579 26943 17582
rect 28625 17579 28691 17582
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 65648 17440 65968 17441
rect 65648 17376 65656 17440
rect 65720 17376 65736 17440
rect 65800 17376 65816 17440
rect 65880 17376 65896 17440
rect 65960 17376 65968 17440
rect 65648 17375 65968 17376
rect 96368 17440 96688 17441
rect 96368 17376 96376 17440
rect 96440 17376 96456 17440
rect 96520 17376 96536 17440
rect 96600 17376 96616 17440
rect 96680 17376 96688 17440
rect 96368 17375 96688 17376
rect 25589 17370 25655 17373
rect 25589 17368 29010 17370
rect 25589 17312 25594 17368
rect 25650 17312 29010 17368
rect 25589 17310 29010 17312
rect 25589 17307 25655 17310
rect 28950 17234 29010 17310
rect 33501 17234 33567 17237
rect 35157 17234 35223 17237
rect 28950 17232 35223 17234
rect 28950 17176 33506 17232
rect 33562 17176 35162 17232
rect 35218 17176 35223 17232
rect 28950 17174 35223 17176
rect 33501 17171 33567 17174
rect 35157 17171 35223 17174
rect 34421 17098 34487 17101
rect 35893 17098 35959 17101
rect 34421 17096 35959 17098
rect 34421 17040 34426 17096
rect 34482 17040 35898 17096
rect 35954 17040 35959 17096
rect 34421 17038 35959 17040
rect 34421 17035 34487 17038
rect 35893 17035 35959 17038
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 50288 16896 50608 16897
rect 50288 16832 50296 16896
rect 50360 16832 50376 16896
rect 50440 16832 50456 16896
rect 50520 16832 50536 16896
rect 50600 16832 50608 16896
rect 50288 16831 50608 16832
rect 81008 16896 81328 16897
rect 81008 16832 81016 16896
rect 81080 16832 81096 16896
rect 81160 16832 81176 16896
rect 81240 16832 81256 16896
rect 81320 16832 81328 16896
rect 81008 16831 81328 16832
rect 40033 16690 40099 16693
rect 46933 16690 46999 16693
rect 40033 16688 46999 16690
rect 40033 16632 40038 16688
rect 40094 16632 46938 16688
rect 46994 16632 46999 16688
rect 40033 16630 46999 16632
rect 40033 16627 40099 16630
rect 46933 16627 46999 16630
rect 24117 16554 24183 16557
rect 26509 16554 26575 16557
rect 24117 16552 26575 16554
rect 24117 16496 24122 16552
rect 24178 16496 26514 16552
rect 26570 16496 26575 16552
rect 24117 16494 26575 16496
rect 24117 16491 24183 16494
rect 26509 16491 26575 16494
rect 31753 16418 31819 16421
rect 34697 16418 34763 16421
rect 31753 16416 34763 16418
rect 31753 16360 31758 16416
rect 31814 16360 34702 16416
rect 34758 16360 34763 16416
rect 31753 16358 34763 16360
rect 31753 16355 31819 16358
rect 34697 16355 34763 16358
rect 46565 16418 46631 16421
rect 46841 16418 46907 16421
rect 46565 16416 46907 16418
rect 46565 16360 46570 16416
rect 46626 16360 46846 16416
rect 46902 16360 46907 16416
rect 46565 16358 46907 16360
rect 46565 16355 46631 16358
rect 46841 16355 46907 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 65648 16352 65968 16353
rect 65648 16288 65656 16352
rect 65720 16288 65736 16352
rect 65800 16288 65816 16352
rect 65880 16288 65896 16352
rect 65960 16288 65968 16352
rect 65648 16287 65968 16288
rect 96368 16352 96688 16353
rect 96368 16288 96376 16352
rect 96440 16288 96456 16352
rect 96520 16288 96536 16352
rect 96600 16288 96616 16352
rect 96680 16288 96688 16352
rect 96368 16287 96688 16288
rect 31385 16282 31451 16285
rect 31753 16282 31819 16285
rect 31385 16280 31819 16282
rect 31385 16224 31390 16280
rect 31446 16224 31758 16280
rect 31814 16224 31819 16280
rect 31385 16222 31819 16224
rect 31385 16219 31451 16222
rect 31753 16219 31819 16222
rect 31385 16146 31451 16149
rect 32029 16146 32095 16149
rect 31385 16144 32095 16146
rect 31385 16088 31390 16144
rect 31446 16088 32034 16144
rect 32090 16088 32095 16144
rect 31385 16086 32095 16088
rect 31385 16083 31451 16086
rect 32029 16083 32095 16086
rect 34053 16146 34119 16149
rect 94129 16146 94195 16149
rect 34053 16144 94195 16146
rect 34053 16088 34058 16144
rect 34114 16088 94134 16144
rect 94190 16088 94195 16144
rect 34053 16086 94195 16088
rect 34053 16083 34119 16086
rect 94129 16083 94195 16086
rect 31017 16010 31083 16013
rect 31753 16010 31819 16013
rect 31017 16008 31819 16010
rect 31017 15952 31022 16008
rect 31078 15952 31758 16008
rect 31814 15952 31819 16008
rect 31017 15950 31819 15952
rect 31017 15947 31083 15950
rect 31753 15947 31819 15950
rect 49509 16010 49575 16013
rect 55857 16010 55923 16013
rect 49509 16008 55923 16010
rect 49509 15952 49514 16008
rect 49570 15952 55862 16008
rect 55918 15952 55923 16008
rect 49509 15950 55923 15952
rect 49509 15947 49575 15950
rect 55857 15947 55923 15950
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 50288 15808 50608 15809
rect 50288 15744 50296 15808
rect 50360 15744 50376 15808
rect 50440 15744 50456 15808
rect 50520 15744 50536 15808
rect 50600 15744 50608 15808
rect 50288 15743 50608 15744
rect 81008 15808 81328 15809
rect 81008 15744 81016 15808
rect 81080 15744 81096 15808
rect 81160 15744 81176 15808
rect 81240 15744 81256 15808
rect 81320 15744 81328 15808
rect 81008 15743 81328 15744
rect 31201 15738 31267 15741
rect 32029 15738 32095 15741
rect 31201 15736 32095 15738
rect 31201 15680 31206 15736
rect 31262 15680 32034 15736
rect 32090 15680 32095 15736
rect 31201 15678 32095 15680
rect 31201 15675 31267 15678
rect 32029 15675 32095 15678
rect 41045 15738 41111 15741
rect 41781 15738 41847 15741
rect 41045 15736 41847 15738
rect 41045 15680 41050 15736
rect 41106 15680 41786 15736
rect 41842 15680 41847 15736
rect 41045 15678 41847 15680
rect 41045 15675 41111 15678
rect 41781 15675 41847 15678
rect 40309 15602 40375 15605
rect 41505 15602 41571 15605
rect 40309 15600 41571 15602
rect 40309 15544 40314 15600
rect 40370 15544 41510 15600
rect 41566 15544 41571 15600
rect 40309 15542 41571 15544
rect 40309 15539 40375 15542
rect 41505 15539 41571 15542
rect 48773 15602 48839 15605
rect 55857 15602 55923 15605
rect 48773 15600 55923 15602
rect 48773 15544 48778 15600
rect 48834 15544 55862 15600
rect 55918 15544 55923 15600
rect 48773 15542 55923 15544
rect 48773 15539 48839 15542
rect 55857 15539 55923 15542
rect 62665 15602 62731 15605
rect 65609 15602 65675 15605
rect 62665 15600 65675 15602
rect 62665 15544 62670 15600
rect 62726 15544 65614 15600
rect 65670 15544 65675 15600
rect 62665 15542 65675 15544
rect 62665 15539 62731 15542
rect 65609 15539 65675 15542
rect 31477 15466 31543 15469
rect 32029 15466 32095 15469
rect 31477 15464 32095 15466
rect 31477 15408 31482 15464
rect 31538 15408 32034 15464
rect 32090 15408 32095 15464
rect 31477 15406 32095 15408
rect 31477 15403 31543 15406
rect 32029 15403 32095 15406
rect 53925 15466 53991 15469
rect 55765 15466 55831 15469
rect 53925 15464 55831 15466
rect 53925 15408 53930 15464
rect 53986 15408 55770 15464
rect 55826 15408 55831 15464
rect 53925 15406 55831 15408
rect 53925 15403 53991 15406
rect 55765 15403 55831 15406
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 65648 15264 65968 15265
rect 65648 15200 65656 15264
rect 65720 15200 65736 15264
rect 65800 15200 65816 15264
rect 65880 15200 65896 15264
rect 65960 15200 65968 15264
rect 65648 15199 65968 15200
rect 96368 15264 96688 15265
rect 96368 15200 96376 15264
rect 96440 15200 96456 15264
rect 96520 15200 96536 15264
rect 96600 15200 96616 15264
rect 96680 15200 96688 15264
rect 96368 15199 96688 15200
rect 20713 15194 20779 15197
rect 19382 15192 20779 15194
rect 19382 15136 20718 15192
rect 20774 15136 20779 15192
rect 19382 15134 20779 15136
rect 19382 15061 19442 15134
rect 20713 15131 20779 15134
rect 70025 15194 70091 15197
rect 70301 15194 70367 15197
rect 70025 15192 70367 15194
rect 70025 15136 70030 15192
rect 70086 15136 70306 15192
rect 70362 15136 70367 15192
rect 70025 15134 70367 15136
rect 70025 15131 70091 15134
rect 70301 15131 70367 15134
rect 19333 15056 19442 15061
rect 19333 15000 19338 15056
rect 19394 15000 19442 15056
rect 19333 14998 19442 15000
rect 19517 15058 19583 15061
rect 19701 15058 19767 15061
rect 98085 15058 98151 15061
rect 19517 15056 19626 15058
rect 19517 15000 19522 15056
rect 19578 15000 19626 15056
rect 19333 14995 19399 14998
rect 19517 14995 19626 15000
rect 19701 15056 98151 15058
rect 19701 15000 19706 15056
rect 19762 15000 98090 15056
rect 98146 15000 98151 15056
rect 19701 14998 98151 15000
rect 19701 14995 19767 14998
rect 98085 14995 98151 14998
rect 19425 14922 19491 14925
rect 19382 14920 19491 14922
rect 19382 14864 19430 14920
rect 19486 14864 19491 14920
rect 19382 14859 19491 14864
rect 19566 14922 19626 14995
rect 20529 14922 20595 14925
rect 19566 14920 20595 14922
rect 19566 14864 20534 14920
rect 20590 14864 20595 14920
rect 19566 14862 20595 14864
rect 20529 14859 20595 14862
rect 33685 14922 33751 14925
rect 36261 14922 36327 14925
rect 33685 14920 36327 14922
rect 33685 14864 33690 14920
rect 33746 14864 36266 14920
rect 36322 14864 36327 14920
rect 33685 14862 36327 14864
rect 33685 14859 33751 14862
rect 36261 14859 36327 14862
rect 51073 14922 51139 14925
rect 57789 14922 57855 14925
rect 51073 14920 57855 14922
rect 51073 14864 51078 14920
rect 51134 14864 57794 14920
rect 57850 14864 57855 14920
rect 51073 14862 57855 14864
rect 51073 14859 51139 14862
rect 57789 14859 57855 14862
rect 58341 14922 58407 14925
rect 62389 14922 62455 14925
rect 58341 14920 62455 14922
rect 58341 14864 58346 14920
rect 58402 14864 62394 14920
rect 62450 14864 62455 14920
rect 58341 14862 62455 14864
rect 58341 14859 58407 14862
rect 62389 14859 62455 14862
rect 19382 14653 19442 14859
rect 69657 14786 69723 14789
rect 71037 14786 71103 14789
rect 69657 14784 71103 14786
rect 69657 14728 69662 14784
rect 69718 14728 71042 14784
rect 71098 14728 71103 14784
rect 69657 14726 71103 14728
rect 69657 14723 69723 14726
rect 71037 14723 71103 14726
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 50288 14720 50608 14721
rect 50288 14656 50296 14720
rect 50360 14656 50376 14720
rect 50440 14656 50456 14720
rect 50520 14656 50536 14720
rect 50600 14656 50608 14720
rect 50288 14655 50608 14656
rect 81008 14720 81328 14721
rect 81008 14656 81016 14720
rect 81080 14656 81096 14720
rect 81160 14656 81176 14720
rect 81240 14656 81256 14720
rect 81320 14656 81328 14720
rect 81008 14655 81328 14656
rect 19333 14648 19442 14653
rect 19333 14592 19338 14648
rect 19394 14592 19442 14648
rect 19333 14590 19442 14592
rect 19333 14587 19399 14590
rect 61009 14514 61075 14517
rect 63677 14514 63743 14517
rect 61009 14512 63743 14514
rect 61009 14456 61014 14512
rect 61070 14456 63682 14512
rect 63738 14456 63743 14512
rect 61009 14454 63743 14456
rect 61009 14451 61075 14454
rect 63677 14451 63743 14454
rect 40401 14378 40467 14381
rect 47209 14378 47275 14381
rect 40401 14376 47275 14378
rect 40401 14320 40406 14376
rect 40462 14320 47214 14376
rect 47270 14320 47275 14376
rect 40401 14318 47275 14320
rect 40401 14315 40467 14318
rect 47209 14315 47275 14318
rect 60273 14378 60339 14381
rect 61101 14378 61167 14381
rect 60273 14376 61167 14378
rect 60273 14320 60278 14376
rect 60334 14320 61106 14376
rect 61162 14320 61167 14376
rect 60273 14318 61167 14320
rect 60273 14315 60339 14318
rect 61101 14315 61167 14318
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 65648 14176 65968 14177
rect 65648 14112 65656 14176
rect 65720 14112 65736 14176
rect 65800 14112 65816 14176
rect 65880 14112 65896 14176
rect 65960 14112 65968 14176
rect 65648 14111 65968 14112
rect 96368 14176 96688 14177
rect 96368 14112 96376 14176
rect 96440 14112 96456 14176
rect 96520 14112 96536 14176
rect 96600 14112 96616 14176
rect 96680 14112 96688 14176
rect 96368 14111 96688 14112
rect 41137 13970 41203 13973
rect 44081 13970 44147 13973
rect 41137 13968 44147 13970
rect 41137 13912 41142 13968
rect 41198 13912 44086 13968
rect 44142 13912 44147 13968
rect 41137 13910 44147 13912
rect 41137 13907 41203 13910
rect 44081 13907 44147 13910
rect 53097 13970 53163 13973
rect 56869 13970 56935 13973
rect 53097 13968 56935 13970
rect 53097 13912 53102 13968
rect 53158 13912 56874 13968
rect 56930 13912 56935 13968
rect 53097 13910 56935 13912
rect 53097 13907 53163 13910
rect 56869 13907 56935 13910
rect 40401 13834 40467 13837
rect 44265 13834 44331 13837
rect 40401 13832 44331 13834
rect 40401 13776 40406 13832
rect 40462 13776 44270 13832
rect 44326 13776 44331 13832
rect 40401 13774 44331 13776
rect 40401 13771 40467 13774
rect 44265 13771 44331 13774
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 50288 13632 50608 13633
rect 50288 13568 50296 13632
rect 50360 13568 50376 13632
rect 50440 13568 50456 13632
rect 50520 13568 50536 13632
rect 50600 13568 50608 13632
rect 50288 13567 50608 13568
rect 81008 13632 81328 13633
rect 81008 13568 81016 13632
rect 81080 13568 81096 13632
rect 81160 13568 81176 13632
rect 81240 13568 81256 13632
rect 81320 13568 81328 13632
rect 81008 13567 81328 13568
rect 22461 13426 22527 13429
rect 27705 13426 27771 13429
rect 22461 13424 27771 13426
rect 22461 13368 22466 13424
rect 22522 13368 27710 13424
rect 27766 13368 27771 13424
rect 22461 13366 27771 13368
rect 22461 13363 22527 13366
rect 27705 13363 27771 13366
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 65648 13088 65968 13089
rect 65648 13024 65656 13088
rect 65720 13024 65736 13088
rect 65800 13024 65816 13088
rect 65880 13024 65896 13088
rect 65960 13024 65968 13088
rect 65648 13023 65968 13024
rect 96368 13088 96688 13089
rect 96368 13024 96376 13088
rect 96440 13024 96456 13088
rect 96520 13024 96536 13088
rect 96600 13024 96616 13088
rect 96680 13024 96688 13088
rect 96368 13023 96688 13024
rect 85573 12882 85639 12885
rect 86033 12882 86099 12885
rect 85573 12880 86099 12882
rect 85573 12824 85578 12880
rect 85634 12824 86038 12880
rect 86094 12824 86099 12880
rect 85573 12822 86099 12824
rect 85573 12819 85639 12822
rect 86033 12819 86099 12822
rect 43529 12746 43595 12749
rect 46197 12746 46263 12749
rect 43529 12744 46263 12746
rect 43529 12688 43534 12744
rect 43590 12688 46202 12744
rect 46258 12688 46263 12744
rect 43529 12686 46263 12688
rect 43529 12683 43595 12686
rect 46197 12683 46263 12686
rect 70209 12610 70275 12613
rect 75913 12610 75979 12613
rect 70209 12608 75979 12610
rect 70209 12552 70214 12608
rect 70270 12552 75918 12608
rect 75974 12552 75979 12608
rect 70209 12550 75979 12552
rect 70209 12547 70275 12550
rect 75913 12547 75979 12550
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 50288 12544 50608 12545
rect 50288 12480 50296 12544
rect 50360 12480 50376 12544
rect 50440 12480 50456 12544
rect 50520 12480 50536 12544
rect 50600 12480 50608 12544
rect 50288 12479 50608 12480
rect 81008 12544 81328 12545
rect 81008 12480 81016 12544
rect 81080 12480 81096 12544
rect 81160 12480 81176 12544
rect 81240 12480 81256 12544
rect 81320 12480 81328 12544
rect 81008 12479 81328 12480
rect 35341 12474 35407 12477
rect 35341 12472 35450 12474
rect 35341 12416 35346 12472
rect 35402 12416 35450 12472
rect 35341 12411 35450 12416
rect 35390 12338 35450 12411
rect 35525 12338 35591 12341
rect 35390 12336 35591 12338
rect 35390 12280 35530 12336
rect 35586 12280 35591 12336
rect 35390 12278 35591 12280
rect 35525 12275 35591 12278
rect 38653 12340 38719 12341
rect 38653 12336 38700 12340
rect 38764 12338 38770 12340
rect 38653 12280 38658 12336
rect 38653 12276 38700 12280
rect 38764 12278 38810 12338
rect 38764 12276 38770 12278
rect 38653 12275 38719 12276
rect 37917 12202 37983 12205
rect 39389 12202 39455 12205
rect 37917 12200 39455 12202
rect 37917 12144 37922 12200
rect 37978 12144 39394 12200
rect 39450 12144 39455 12200
rect 37917 12142 39455 12144
rect 37917 12139 37983 12142
rect 39389 12139 39455 12142
rect 41689 12202 41755 12205
rect 48037 12202 48103 12205
rect 41689 12200 48103 12202
rect 41689 12144 41694 12200
rect 41750 12144 48042 12200
rect 48098 12144 48103 12200
rect 41689 12142 48103 12144
rect 41689 12139 41755 12142
rect 48037 12139 48103 12142
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 65648 12000 65968 12001
rect 65648 11936 65656 12000
rect 65720 11936 65736 12000
rect 65800 11936 65816 12000
rect 65880 11936 65896 12000
rect 65960 11936 65968 12000
rect 65648 11935 65968 11936
rect 96368 12000 96688 12001
rect 96368 11936 96376 12000
rect 96440 11936 96456 12000
rect 96520 11936 96536 12000
rect 96600 11936 96616 12000
rect 96680 11936 96688 12000
rect 96368 11935 96688 11936
rect 38837 11930 38903 11933
rect 38702 11928 38903 11930
rect 38702 11872 38842 11928
rect 38898 11872 38903 11928
rect 38702 11870 38903 11872
rect 34789 11522 34855 11525
rect 38561 11522 38627 11525
rect 34789 11520 38627 11522
rect 34789 11464 34794 11520
rect 34850 11464 38566 11520
rect 38622 11464 38627 11520
rect 34789 11462 38627 11464
rect 34789 11459 34855 11462
rect 38561 11459 38627 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 38702 11389 38762 11870
rect 38837 11867 38903 11870
rect 50288 11456 50608 11457
rect 50288 11392 50296 11456
rect 50360 11392 50376 11456
rect 50440 11392 50456 11456
rect 50520 11392 50536 11456
rect 50600 11392 50608 11456
rect 50288 11391 50608 11392
rect 81008 11456 81328 11457
rect 81008 11392 81016 11456
rect 81080 11392 81096 11456
rect 81160 11392 81176 11456
rect 81240 11392 81256 11456
rect 81320 11392 81328 11456
rect 81008 11391 81328 11392
rect 38009 11386 38075 11389
rect 38469 11388 38535 11389
rect 38469 11386 38516 11388
rect 38009 11384 38516 11386
rect 38009 11328 38014 11384
rect 38070 11328 38474 11384
rect 38009 11326 38516 11328
rect 38009 11323 38075 11326
rect 38469 11324 38516 11326
rect 38580 11324 38586 11388
rect 38653 11384 38762 11389
rect 38653 11328 38658 11384
rect 38714 11328 38762 11384
rect 38653 11326 38762 11328
rect 38929 11386 38995 11389
rect 39389 11386 39455 11389
rect 38929 11384 39455 11386
rect 38929 11328 38934 11384
rect 38990 11328 39394 11384
rect 39450 11328 39455 11384
rect 38929 11326 39455 11328
rect 38469 11323 38535 11324
rect 38653 11323 38719 11326
rect 38929 11323 38995 11326
rect 39389 11323 39455 11326
rect 12341 11250 12407 11253
rect 12801 11250 12867 11253
rect 12341 11248 12867 11250
rect 12341 11192 12346 11248
rect 12402 11192 12806 11248
rect 12862 11192 12867 11248
rect 12341 11190 12867 11192
rect 12341 11187 12407 11190
rect 12801 11187 12867 11190
rect 13077 11250 13143 11253
rect 89253 11250 89319 11253
rect 13077 11248 89319 11250
rect 13077 11192 13082 11248
rect 13138 11192 89258 11248
rect 89314 11192 89319 11248
rect 13077 11190 89319 11192
rect 13077 11187 13143 11190
rect 89253 11187 89319 11190
rect 12525 11114 12591 11117
rect 16021 11114 16087 11117
rect 38745 11116 38811 11117
rect 12525 11112 16087 11114
rect 12525 11056 12530 11112
rect 12586 11056 16026 11112
rect 16082 11056 16087 11112
rect 12525 11054 16087 11056
rect 12525 11051 12591 11054
rect 16021 11051 16087 11054
rect 38694 11052 38700 11116
rect 38764 11114 38811 11116
rect 62941 11114 63007 11117
rect 65057 11114 65123 11117
rect 38764 11112 38856 11114
rect 38806 11056 38856 11112
rect 38764 11054 38856 11056
rect 62941 11112 65123 11114
rect 62941 11056 62946 11112
rect 63002 11056 65062 11112
rect 65118 11056 65123 11112
rect 62941 11054 65123 11056
rect 38764 11052 38811 11054
rect 38745 11051 38811 11052
rect 62941 11051 63007 11054
rect 65057 11051 65123 11054
rect 37917 10978 37983 10981
rect 39573 10978 39639 10981
rect 37917 10976 39639 10978
rect 37917 10920 37922 10976
rect 37978 10920 39578 10976
rect 39634 10920 39639 10976
rect 37917 10918 39639 10920
rect 37917 10915 37983 10918
rect 39573 10915 39639 10918
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 65648 10912 65968 10913
rect 65648 10848 65656 10912
rect 65720 10848 65736 10912
rect 65800 10848 65816 10912
rect 65880 10848 65896 10912
rect 65960 10848 65968 10912
rect 65648 10847 65968 10848
rect 96368 10912 96688 10913
rect 96368 10848 96376 10912
rect 96440 10848 96456 10912
rect 96520 10848 96536 10912
rect 96600 10848 96616 10912
rect 96680 10848 96688 10912
rect 96368 10847 96688 10848
rect 41137 10706 41203 10709
rect 41689 10706 41755 10709
rect 41137 10704 41755 10706
rect 41137 10648 41142 10704
rect 41198 10648 41694 10704
rect 41750 10648 41755 10704
rect 41137 10646 41755 10648
rect 41137 10643 41203 10646
rect 41689 10643 41755 10646
rect 44265 10706 44331 10709
rect 46565 10706 46631 10709
rect 44265 10704 46631 10706
rect 44265 10648 44270 10704
rect 44326 10648 46570 10704
rect 46626 10648 46631 10704
rect 44265 10646 46631 10648
rect 44265 10643 44331 10646
rect 46565 10643 46631 10646
rect 41781 10570 41847 10573
rect 44633 10570 44699 10573
rect 41781 10568 44699 10570
rect 41781 10512 41786 10568
rect 41842 10512 44638 10568
rect 44694 10512 44699 10568
rect 41781 10510 44699 10512
rect 41781 10507 41847 10510
rect 44633 10507 44699 10510
rect 68277 10570 68343 10573
rect 69105 10570 69171 10573
rect 68277 10568 69171 10570
rect 68277 10512 68282 10568
rect 68338 10512 69110 10568
rect 69166 10512 69171 10568
rect 68277 10510 69171 10512
rect 68277 10507 68343 10510
rect 69105 10507 69171 10510
rect 36445 10434 36511 10437
rect 37181 10434 37247 10437
rect 44081 10434 44147 10437
rect 36445 10432 44147 10434
rect 36445 10376 36450 10432
rect 36506 10376 37186 10432
rect 37242 10376 44086 10432
rect 44142 10376 44147 10432
rect 36445 10374 44147 10376
rect 36445 10371 36511 10374
rect 37181 10371 37247 10374
rect 44081 10371 44147 10374
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 50288 10368 50608 10369
rect 50288 10304 50296 10368
rect 50360 10304 50376 10368
rect 50440 10304 50456 10368
rect 50520 10304 50536 10368
rect 50600 10304 50608 10368
rect 50288 10303 50608 10304
rect 81008 10368 81328 10369
rect 81008 10304 81016 10368
rect 81080 10304 81096 10368
rect 81160 10304 81176 10368
rect 81240 10304 81256 10368
rect 81320 10304 81328 10368
rect 81008 10303 81328 10304
rect 25129 10298 25195 10301
rect 26325 10298 26391 10301
rect 25129 10296 26391 10298
rect 25129 10240 25134 10296
rect 25190 10240 26330 10296
rect 26386 10240 26391 10296
rect 25129 10238 26391 10240
rect 25129 10235 25195 10238
rect 26325 10235 26391 10238
rect 33225 10162 33291 10165
rect 38193 10162 38259 10165
rect 33225 10160 38259 10162
rect 33225 10104 33230 10160
rect 33286 10104 38198 10160
rect 38254 10104 38259 10160
rect 33225 10102 38259 10104
rect 33225 10099 33291 10102
rect 38193 10099 38259 10102
rect 68645 10162 68711 10165
rect 71681 10162 71747 10165
rect 68645 10160 71747 10162
rect 68645 10104 68650 10160
rect 68706 10104 71686 10160
rect 71742 10104 71747 10160
rect 68645 10102 71747 10104
rect 68645 10099 68711 10102
rect 71681 10099 71747 10102
rect 43989 10026 44055 10029
rect 46657 10026 46723 10029
rect 43989 10024 46723 10026
rect 43989 9968 43994 10024
rect 44050 9968 46662 10024
rect 46718 9968 46723 10024
rect 43989 9966 46723 9968
rect 43989 9963 44055 9966
rect 46657 9963 46723 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 65648 9824 65968 9825
rect 65648 9760 65656 9824
rect 65720 9760 65736 9824
rect 65800 9760 65816 9824
rect 65880 9760 65896 9824
rect 65960 9760 65968 9824
rect 65648 9759 65968 9760
rect 96368 9824 96688 9825
rect 96368 9760 96376 9824
rect 96440 9760 96456 9824
rect 96520 9760 96536 9824
rect 96600 9760 96616 9824
rect 96680 9760 96688 9824
rect 96368 9759 96688 9760
rect 68277 9754 68343 9757
rect 69933 9754 69999 9757
rect 68277 9752 69999 9754
rect 68277 9696 68282 9752
rect 68338 9696 69938 9752
rect 69994 9696 69999 9752
rect 68277 9694 69999 9696
rect 68277 9691 68343 9694
rect 69933 9691 69999 9694
rect 35985 9618 36051 9621
rect 37273 9618 37339 9621
rect 35985 9616 37339 9618
rect 35985 9560 35990 9616
rect 36046 9560 37278 9616
rect 37334 9560 37339 9616
rect 35985 9558 37339 9560
rect 35985 9555 36051 9558
rect 37273 9555 37339 9558
rect 3233 9482 3299 9485
rect 51809 9482 51875 9485
rect 3233 9480 51875 9482
rect 3233 9424 3238 9480
rect 3294 9424 51814 9480
rect 51870 9424 51875 9480
rect 3233 9422 51875 9424
rect 3233 9419 3299 9422
rect 51809 9419 51875 9422
rect 62389 9482 62455 9485
rect 65517 9482 65583 9485
rect 62389 9480 65583 9482
rect 62389 9424 62394 9480
rect 62450 9424 65522 9480
rect 65578 9424 65583 9480
rect 62389 9422 65583 9424
rect 62389 9419 62455 9422
rect 65517 9419 65583 9422
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 50288 9280 50608 9281
rect 50288 9216 50296 9280
rect 50360 9216 50376 9280
rect 50440 9216 50456 9280
rect 50520 9216 50536 9280
rect 50600 9216 50608 9280
rect 50288 9215 50608 9216
rect 81008 9280 81328 9281
rect 81008 9216 81016 9280
rect 81080 9216 81096 9280
rect 81160 9216 81176 9280
rect 81240 9216 81256 9280
rect 81320 9216 81328 9280
rect 81008 9215 81328 9216
rect 11789 9074 11855 9077
rect 95969 9074 96035 9077
rect 11789 9072 96035 9074
rect 11789 9016 11794 9072
rect 11850 9016 95974 9072
rect 96030 9016 96035 9072
rect 11789 9014 96035 9016
rect 11789 9011 11855 9014
rect 95969 9011 96035 9014
rect 61653 8938 61719 8941
rect 65057 8938 65123 8941
rect 61653 8936 65123 8938
rect 61653 8880 61658 8936
rect 61714 8880 65062 8936
rect 65118 8880 65123 8936
rect 61653 8878 65123 8880
rect 61653 8875 61719 8878
rect 65057 8875 65123 8878
rect 51809 8802 51875 8805
rect 56501 8802 56567 8805
rect 51809 8800 56567 8802
rect 51809 8744 51814 8800
rect 51870 8744 56506 8800
rect 56562 8744 56567 8800
rect 51809 8742 56567 8744
rect 51809 8739 51875 8742
rect 56501 8739 56567 8742
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 65648 8736 65968 8737
rect 65648 8672 65656 8736
rect 65720 8672 65736 8736
rect 65800 8672 65816 8736
rect 65880 8672 65896 8736
rect 65960 8672 65968 8736
rect 65648 8671 65968 8672
rect 96368 8736 96688 8737
rect 96368 8672 96376 8736
rect 96440 8672 96456 8736
rect 96520 8672 96536 8736
rect 96600 8672 96616 8736
rect 96680 8672 96688 8736
rect 96368 8671 96688 8672
rect 59261 8666 59327 8669
rect 60825 8666 60891 8669
rect 59261 8664 60891 8666
rect 59261 8608 59266 8664
rect 59322 8608 60830 8664
rect 60886 8608 60891 8664
rect 59261 8606 60891 8608
rect 59261 8603 59327 8606
rect 60825 8603 60891 8606
rect 61653 8666 61719 8669
rect 63309 8666 63375 8669
rect 61653 8664 63375 8666
rect 61653 8608 61658 8664
rect 61714 8608 63314 8664
rect 63370 8608 63375 8664
rect 61653 8606 63375 8608
rect 61653 8603 61719 8606
rect 63309 8603 63375 8606
rect 50797 8530 50863 8533
rect 51073 8530 51139 8533
rect 50797 8528 51139 8530
rect 50797 8472 50802 8528
rect 50858 8472 51078 8528
rect 51134 8472 51139 8528
rect 50797 8470 51139 8472
rect 50797 8467 50863 8470
rect 51073 8467 51139 8470
rect 60733 8530 60799 8533
rect 62205 8530 62271 8533
rect 60733 8528 62271 8530
rect 60733 8472 60738 8528
rect 60794 8472 62210 8528
rect 62266 8472 62271 8528
rect 60733 8470 62271 8472
rect 60733 8467 60799 8470
rect 62205 8467 62271 8470
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 50288 8192 50608 8193
rect 50288 8128 50296 8192
rect 50360 8128 50376 8192
rect 50440 8128 50456 8192
rect 50520 8128 50536 8192
rect 50600 8128 50608 8192
rect 50288 8127 50608 8128
rect 81008 8192 81328 8193
rect 81008 8128 81016 8192
rect 81080 8128 81096 8192
rect 81160 8128 81176 8192
rect 81240 8128 81256 8192
rect 81320 8128 81328 8192
rect 81008 8127 81328 8128
rect 38837 8122 38903 8125
rect 39481 8122 39547 8125
rect 38837 8120 39547 8122
rect 38837 8064 38842 8120
rect 38898 8064 39486 8120
rect 39542 8064 39547 8120
rect 38837 8062 39547 8064
rect 38837 8059 38903 8062
rect 39481 8059 39547 8062
rect 10041 7986 10107 7989
rect 65149 7986 65215 7989
rect 10041 7984 65215 7986
rect 10041 7928 10046 7984
rect 10102 7928 65154 7984
rect 65210 7928 65215 7984
rect 10041 7926 65215 7928
rect 10041 7923 10107 7926
rect 65149 7923 65215 7926
rect 2681 7850 2747 7853
rect 47393 7850 47459 7853
rect 2681 7848 47459 7850
rect 2681 7792 2686 7848
rect 2742 7792 47398 7848
rect 47454 7792 47459 7848
rect 2681 7790 47459 7792
rect 2681 7787 2747 7790
rect 47393 7787 47459 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 65648 7648 65968 7649
rect 65648 7584 65656 7648
rect 65720 7584 65736 7648
rect 65800 7584 65816 7648
rect 65880 7584 65896 7648
rect 65960 7584 65968 7648
rect 65648 7583 65968 7584
rect 96368 7648 96688 7649
rect 96368 7584 96376 7648
rect 96440 7584 96456 7648
rect 96520 7584 96536 7648
rect 96600 7584 96616 7648
rect 96680 7584 96688 7648
rect 96368 7583 96688 7584
rect 12157 7442 12223 7445
rect 74165 7442 74231 7445
rect 12157 7440 74231 7442
rect 12157 7384 12162 7440
rect 12218 7384 74170 7440
rect 74226 7384 74231 7440
rect 12157 7382 74231 7384
rect 12157 7379 12223 7382
rect 74165 7379 74231 7382
rect 24761 7306 24827 7309
rect 25681 7306 25747 7309
rect 25957 7306 26023 7309
rect 85573 7306 85639 7309
rect 24761 7304 85639 7306
rect 24761 7248 24766 7304
rect 24822 7248 25686 7304
rect 25742 7248 25962 7304
rect 26018 7248 85578 7304
rect 85634 7248 85639 7304
rect 24761 7246 85639 7248
rect 24761 7243 24827 7246
rect 25681 7243 25747 7246
rect 25957 7243 26023 7246
rect 85573 7243 85639 7246
rect 24117 7170 24183 7173
rect 25957 7170 26023 7173
rect 24117 7168 26023 7170
rect 24117 7112 24122 7168
rect 24178 7112 25962 7168
rect 26018 7112 26023 7168
rect 24117 7110 26023 7112
rect 24117 7107 24183 7110
rect 25957 7107 26023 7110
rect 48865 7170 48931 7173
rect 50153 7170 50219 7173
rect 48865 7168 50219 7170
rect 48865 7112 48870 7168
rect 48926 7112 50158 7168
rect 50214 7112 50219 7168
rect 48865 7110 50219 7112
rect 48865 7107 48931 7110
rect 50153 7107 50219 7110
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 50288 7104 50608 7105
rect 50288 7040 50296 7104
rect 50360 7040 50376 7104
rect 50440 7040 50456 7104
rect 50520 7040 50536 7104
rect 50600 7040 50608 7104
rect 50288 7039 50608 7040
rect 81008 7104 81328 7105
rect 81008 7040 81016 7104
rect 81080 7040 81096 7104
rect 81160 7040 81176 7104
rect 81240 7040 81256 7104
rect 81320 7040 81328 7104
rect 81008 7039 81328 7040
rect 21817 6762 21883 6765
rect 74533 6762 74599 6765
rect 21817 6760 74599 6762
rect 21817 6704 21822 6760
rect 21878 6704 74538 6760
rect 74594 6704 74599 6760
rect 21817 6702 74599 6704
rect 21817 6699 21883 6702
rect 74533 6699 74599 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 65648 6560 65968 6561
rect 65648 6496 65656 6560
rect 65720 6496 65736 6560
rect 65800 6496 65816 6560
rect 65880 6496 65896 6560
rect 65960 6496 65968 6560
rect 65648 6495 65968 6496
rect 96368 6560 96688 6561
rect 96368 6496 96376 6560
rect 96440 6496 96456 6560
rect 96520 6496 96536 6560
rect 96600 6496 96616 6560
rect 96680 6496 96688 6560
rect 96368 6495 96688 6496
rect 5441 6354 5507 6357
rect 52361 6354 52427 6357
rect 5441 6352 52427 6354
rect 5441 6296 5446 6352
rect 5502 6296 52366 6352
rect 52422 6296 52427 6352
rect 5441 6294 52427 6296
rect 5441 6291 5507 6294
rect 52361 6291 52427 6294
rect 52729 6354 52795 6357
rect 53189 6354 53255 6357
rect 52729 6352 53255 6354
rect 52729 6296 52734 6352
rect 52790 6296 53194 6352
rect 53250 6296 53255 6352
rect 52729 6294 53255 6296
rect 52729 6291 52795 6294
rect 53189 6291 53255 6294
rect 3049 6218 3115 6221
rect 75637 6218 75703 6221
rect 3049 6216 75703 6218
rect 3049 6160 3054 6216
rect 3110 6160 75642 6216
rect 75698 6160 75703 6216
rect 3049 6158 75703 6160
rect 3049 6155 3115 6158
rect 75637 6155 75703 6158
rect 20345 6082 20411 6085
rect 21817 6082 21883 6085
rect 20345 6080 21883 6082
rect 20345 6024 20350 6080
rect 20406 6024 21822 6080
rect 21878 6024 21883 6080
rect 20345 6022 21883 6024
rect 20345 6019 20411 6022
rect 21817 6019 21883 6022
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 50288 6016 50608 6017
rect 50288 5952 50296 6016
rect 50360 5952 50376 6016
rect 50440 5952 50456 6016
rect 50520 5952 50536 6016
rect 50600 5952 50608 6016
rect 50288 5951 50608 5952
rect 81008 6016 81328 6017
rect 81008 5952 81016 6016
rect 81080 5952 81096 6016
rect 81160 5952 81176 6016
rect 81240 5952 81256 6016
rect 81320 5952 81328 6016
rect 81008 5951 81328 5952
rect 7649 5674 7715 5677
rect 8753 5674 8819 5677
rect 7649 5672 8819 5674
rect 7649 5616 7654 5672
rect 7710 5616 8758 5672
rect 8814 5616 8819 5672
rect 7649 5614 8819 5616
rect 7649 5611 7715 5614
rect 8753 5611 8819 5614
rect 5073 5538 5139 5541
rect 8477 5538 8543 5541
rect 5073 5536 8543 5538
rect 5073 5480 5078 5536
rect 5134 5480 8482 5536
rect 8538 5480 8543 5536
rect 5073 5478 8543 5480
rect 5073 5475 5139 5478
rect 8477 5475 8543 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 65648 5472 65968 5473
rect 65648 5408 65656 5472
rect 65720 5408 65736 5472
rect 65800 5408 65816 5472
rect 65880 5408 65896 5472
rect 65960 5408 65968 5472
rect 65648 5407 65968 5408
rect 96368 5472 96688 5473
rect 96368 5408 96376 5472
rect 96440 5408 96456 5472
rect 96520 5408 96536 5472
rect 96600 5408 96616 5472
rect 96680 5408 96688 5472
rect 96368 5407 96688 5408
rect 18873 5266 18939 5269
rect 90449 5266 90515 5269
rect 90817 5266 90883 5269
rect 18873 5264 90883 5266
rect 18873 5208 18878 5264
rect 18934 5208 90454 5264
rect 90510 5208 90822 5264
rect 90878 5208 90883 5264
rect 18873 5206 90883 5208
rect 18873 5203 18939 5206
rect 90449 5203 90515 5206
rect 90817 5203 90883 5206
rect 59077 5130 59143 5133
rect 65149 5130 65215 5133
rect 59077 5128 65215 5130
rect 59077 5072 59082 5128
rect 59138 5072 65154 5128
rect 65210 5072 65215 5128
rect 59077 5070 65215 5072
rect 59077 5067 59143 5070
rect 65149 5067 65215 5070
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 50288 4928 50608 4929
rect 50288 4864 50296 4928
rect 50360 4864 50376 4928
rect 50440 4864 50456 4928
rect 50520 4864 50536 4928
rect 50600 4864 50608 4928
rect 50288 4863 50608 4864
rect 81008 4928 81328 4929
rect 81008 4864 81016 4928
rect 81080 4864 81096 4928
rect 81160 4864 81176 4928
rect 81240 4864 81256 4928
rect 81320 4864 81328 4928
rect 81008 4863 81328 4864
rect 62021 4722 62087 4725
rect 64413 4722 64479 4725
rect 62021 4720 64479 4722
rect 62021 4664 62026 4720
rect 62082 4664 64418 4720
rect 64474 4664 64479 4720
rect 62021 4662 64479 4664
rect 62021 4659 62087 4662
rect 64413 4659 64479 4662
rect 61745 4586 61811 4589
rect 62849 4586 62915 4589
rect 61745 4584 62915 4586
rect 61745 4528 61750 4584
rect 61806 4528 62854 4584
rect 62910 4528 62915 4584
rect 61745 4526 62915 4528
rect 61745 4523 61811 4526
rect 62849 4523 62915 4526
rect 62021 4450 62087 4453
rect 64965 4450 65031 4453
rect 62021 4448 65031 4450
rect 62021 4392 62026 4448
rect 62082 4392 64970 4448
rect 65026 4392 65031 4448
rect 62021 4390 65031 4392
rect 62021 4387 62087 4390
rect 64965 4387 65031 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 65648 4384 65968 4385
rect 65648 4320 65656 4384
rect 65720 4320 65736 4384
rect 65800 4320 65816 4384
rect 65880 4320 65896 4384
rect 65960 4320 65968 4384
rect 65648 4319 65968 4320
rect 96368 4384 96688 4385
rect 96368 4320 96376 4384
rect 96440 4320 96456 4384
rect 96520 4320 96536 4384
rect 96600 4320 96616 4384
rect 96680 4320 96688 4384
rect 96368 4319 96688 4320
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 50288 3840 50608 3841
rect 50288 3776 50296 3840
rect 50360 3776 50376 3840
rect 50440 3776 50456 3840
rect 50520 3776 50536 3840
rect 50600 3776 50608 3840
rect 50288 3775 50608 3776
rect 81008 3840 81328 3841
rect 81008 3776 81016 3840
rect 81080 3776 81096 3840
rect 81160 3776 81176 3840
rect 81240 3776 81256 3840
rect 81320 3776 81328 3840
rect 81008 3775 81328 3776
rect 20161 3770 20227 3773
rect 26417 3770 26483 3773
rect 49785 3770 49851 3773
rect 20161 3768 26483 3770
rect 20161 3712 20166 3768
rect 20222 3712 26422 3768
rect 26478 3712 26483 3768
rect 20161 3710 26483 3712
rect 20161 3707 20227 3710
rect 26417 3707 26483 3710
rect 49742 3768 49851 3770
rect 49742 3712 49790 3768
rect 49846 3712 49851 3768
rect 49742 3707 49851 3712
rect 17585 3634 17651 3637
rect 18137 3634 18203 3637
rect 17585 3632 18203 3634
rect 17585 3576 17590 3632
rect 17646 3576 18142 3632
rect 18198 3576 18203 3632
rect 17585 3574 18203 3576
rect 17585 3571 17651 3574
rect 18137 3571 18203 3574
rect 20621 3634 20687 3637
rect 22277 3634 22343 3637
rect 20621 3632 22343 3634
rect 20621 3576 20626 3632
rect 20682 3576 22282 3632
rect 22338 3576 22343 3632
rect 20621 3574 22343 3576
rect 20621 3571 20687 3574
rect 22277 3571 22343 3574
rect 49742 3501 49802 3707
rect 17217 3498 17283 3501
rect 18229 3498 18295 3501
rect 17217 3496 18295 3498
rect 17217 3440 17222 3496
rect 17278 3440 18234 3496
rect 18290 3440 18295 3496
rect 17217 3438 18295 3440
rect 17217 3435 17283 3438
rect 18229 3435 18295 3438
rect 21725 3498 21791 3501
rect 21725 3496 21834 3498
rect 21725 3440 21730 3496
rect 21786 3440 21834 3496
rect 21725 3435 21834 3440
rect 49742 3496 49851 3501
rect 49742 3440 49790 3496
rect 49846 3440 49851 3496
rect 49742 3438 49851 3440
rect 49785 3435 49851 3438
rect 17861 3362 17927 3365
rect 18137 3362 18203 3365
rect 17861 3360 18203 3362
rect 17861 3304 17866 3360
rect 17922 3304 18142 3360
rect 18198 3304 18203 3360
rect 17861 3302 18203 3304
rect 21774 3362 21834 3435
rect 22001 3362 22067 3365
rect 21774 3360 22067 3362
rect 21774 3304 22006 3360
rect 22062 3304 22067 3360
rect 21774 3302 22067 3304
rect 17861 3299 17927 3302
rect 18137 3299 18203 3302
rect 22001 3299 22067 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 65648 3296 65968 3297
rect 65648 3232 65656 3296
rect 65720 3232 65736 3296
rect 65800 3232 65816 3296
rect 65880 3232 65896 3296
rect 65960 3232 65968 3296
rect 65648 3231 65968 3232
rect 96368 3296 96688 3297
rect 96368 3232 96376 3296
rect 96440 3232 96456 3296
rect 96520 3232 96536 3296
rect 96600 3232 96616 3296
rect 96680 3232 96688 3296
rect 96368 3231 96688 3232
rect 19057 2954 19123 2957
rect 20069 2954 20135 2957
rect 26141 2954 26207 2957
rect 19057 2952 20135 2954
rect 19057 2896 19062 2952
rect 19118 2896 20074 2952
rect 20130 2896 20135 2952
rect 19057 2894 20135 2896
rect 19057 2891 19123 2894
rect 20069 2891 20135 2894
rect 25638 2952 26207 2954
rect 25638 2896 26146 2952
rect 26202 2896 26207 2952
rect 25638 2894 26207 2896
rect 25638 2821 25698 2894
rect 26141 2891 26207 2894
rect 25589 2816 25698 2821
rect 25589 2760 25594 2816
rect 25650 2760 25698 2816
rect 25589 2758 25698 2760
rect 25589 2755 25655 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 50288 2752 50608 2753
rect 50288 2688 50296 2752
rect 50360 2688 50376 2752
rect 50440 2688 50456 2752
rect 50520 2688 50536 2752
rect 50600 2688 50608 2752
rect 50288 2687 50608 2688
rect 81008 2752 81328 2753
rect 81008 2688 81016 2752
rect 81080 2688 81096 2752
rect 81160 2688 81176 2752
rect 81240 2688 81256 2752
rect 81320 2688 81328 2752
rect 81008 2687 81328 2688
rect 20161 2682 20227 2685
rect 21173 2682 21239 2685
rect 20161 2680 21239 2682
rect 20161 2624 20166 2680
rect 20222 2624 21178 2680
rect 21234 2624 21239 2680
rect 20161 2622 21239 2624
rect 20161 2619 20227 2622
rect 21173 2619 21239 2622
rect 71957 2546 72023 2549
rect 72325 2546 72391 2549
rect 71957 2544 72391 2546
rect 71957 2488 71962 2544
rect 72018 2488 72330 2544
rect 72386 2488 72391 2544
rect 71957 2486 72391 2488
rect 71957 2483 72023 2486
rect 72325 2483 72391 2486
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 65648 2208 65968 2209
rect 65648 2144 65656 2208
rect 65720 2144 65736 2208
rect 65800 2144 65816 2208
rect 65880 2144 65896 2208
rect 65960 2144 65968 2208
rect 65648 2143 65968 2144
rect 96368 2208 96688 2209
rect 96368 2144 96376 2208
rect 96440 2144 96456 2208
rect 96520 2144 96536 2208
rect 96600 2144 96616 2208
rect 96680 2144 96688 2208
rect 96368 2143 96688 2144
rect 46473 1322 46539 1325
rect 87965 1322 88031 1325
rect 46473 1320 88031 1322
rect 46473 1264 46478 1320
rect 46534 1264 87970 1320
rect 88026 1264 88031 1320
rect 46473 1262 88031 1264
rect 46473 1259 46539 1262
rect 87965 1259 88031 1262
rect 17493 1186 17559 1189
rect 88425 1186 88491 1189
rect 17493 1184 88491 1186
rect 17493 1128 17498 1184
rect 17554 1128 88430 1184
rect 88486 1128 88491 1184
rect 17493 1126 88491 1128
rect 17493 1123 17559 1126
rect 88425 1123 88491 1126
rect 21541 1050 21607 1053
rect 85113 1050 85179 1053
rect 21541 1048 85179 1050
rect 21541 992 21546 1048
rect 21602 992 85118 1048
rect 85174 992 85179 1048
rect 21541 990 85179 992
rect 21541 987 21607 990
rect 85113 987 85179 990
rect 20713 914 20779 917
rect 77753 914 77819 917
rect 20713 912 77819 914
rect 20713 856 20718 912
rect 20774 856 77758 912
rect 77814 856 77819 912
rect 20713 854 77819 856
rect 20713 851 20779 854
rect 77753 851 77819 854
rect 2221 778 2287 781
rect 55489 778 55555 781
rect 2221 776 55555 778
rect 2221 720 2226 776
rect 2282 720 55494 776
rect 55550 720 55555 776
rect 2221 718 55555 720
rect 2221 715 2287 718
rect 55489 715 55555 718
rect 33041 642 33107 645
rect 82077 642 82143 645
rect 33041 640 82143 642
rect 33041 584 33046 640
rect 33102 584 82082 640
rect 82138 584 82143 640
rect 33041 582 82143 584
rect 33041 579 33107 582
rect 82077 579 82143 582
rect 27429 506 27495 509
rect 67449 506 67515 509
rect 27429 504 67515 506
rect 27429 448 27434 504
rect 27490 448 67454 504
rect 67510 448 67515 504
rect 27429 446 67515 448
rect 27429 443 27495 446
rect 67449 443 67515 446
rect 38561 370 38627 373
rect 77385 370 77451 373
rect 38561 368 77451 370
rect 38561 312 38566 368
rect 38622 312 77390 368
rect 77446 312 77451 368
rect 38561 310 77451 312
rect 38561 307 38627 310
rect 77385 307 77451 310
rect 2405 234 2471 237
rect 75545 234 75611 237
rect 2405 232 75611 234
rect 2405 176 2410 232
rect 2466 176 75550 232
rect 75606 176 75611 232
rect 2405 174 75611 176
rect 2405 171 2471 174
rect 75545 171 75611 174
<< via3 >>
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 50296 37564 50360 37568
rect 50296 37508 50300 37564
rect 50300 37508 50356 37564
rect 50356 37508 50360 37564
rect 50296 37504 50360 37508
rect 50376 37564 50440 37568
rect 50376 37508 50380 37564
rect 50380 37508 50436 37564
rect 50436 37508 50440 37564
rect 50376 37504 50440 37508
rect 50456 37564 50520 37568
rect 50456 37508 50460 37564
rect 50460 37508 50516 37564
rect 50516 37508 50520 37564
rect 50456 37504 50520 37508
rect 50536 37564 50600 37568
rect 50536 37508 50540 37564
rect 50540 37508 50596 37564
rect 50596 37508 50600 37564
rect 50536 37504 50600 37508
rect 81016 37564 81080 37568
rect 81016 37508 81020 37564
rect 81020 37508 81076 37564
rect 81076 37508 81080 37564
rect 81016 37504 81080 37508
rect 81096 37564 81160 37568
rect 81096 37508 81100 37564
rect 81100 37508 81156 37564
rect 81156 37508 81160 37564
rect 81096 37504 81160 37508
rect 81176 37564 81240 37568
rect 81176 37508 81180 37564
rect 81180 37508 81236 37564
rect 81236 37508 81240 37564
rect 81176 37504 81240 37508
rect 81256 37564 81320 37568
rect 81256 37508 81260 37564
rect 81260 37508 81316 37564
rect 81316 37508 81320 37564
rect 81256 37504 81320 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 65656 37020 65720 37024
rect 65656 36964 65660 37020
rect 65660 36964 65716 37020
rect 65716 36964 65720 37020
rect 65656 36960 65720 36964
rect 65736 37020 65800 37024
rect 65736 36964 65740 37020
rect 65740 36964 65796 37020
rect 65796 36964 65800 37020
rect 65736 36960 65800 36964
rect 65816 37020 65880 37024
rect 65816 36964 65820 37020
rect 65820 36964 65876 37020
rect 65876 36964 65880 37020
rect 65816 36960 65880 36964
rect 65896 37020 65960 37024
rect 65896 36964 65900 37020
rect 65900 36964 65956 37020
rect 65956 36964 65960 37020
rect 65896 36960 65960 36964
rect 96376 37020 96440 37024
rect 96376 36964 96380 37020
rect 96380 36964 96436 37020
rect 96436 36964 96440 37020
rect 96376 36960 96440 36964
rect 96456 37020 96520 37024
rect 96456 36964 96460 37020
rect 96460 36964 96516 37020
rect 96516 36964 96520 37020
rect 96456 36960 96520 36964
rect 96536 37020 96600 37024
rect 96536 36964 96540 37020
rect 96540 36964 96596 37020
rect 96596 36964 96600 37020
rect 96536 36960 96600 36964
rect 96616 37020 96680 37024
rect 96616 36964 96620 37020
rect 96620 36964 96676 37020
rect 96676 36964 96680 37020
rect 96616 36960 96680 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 50296 36476 50360 36480
rect 50296 36420 50300 36476
rect 50300 36420 50356 36476
rect 50356 36420 50360 36476
rect 50296 36416 50360 36420
rect 50376 36476 50440 36480
rect 50376 36420 50380 36476
rect 50380 36420 50436 36476
rect 50436 36420 50440 36476
rect 50376 36416 50440 36420
rect 50456 36476 50520 36480
rect 50456 36420 50460 36476
rect 50460 36420 50516 36476
rect 50516 36420 50520 36476
rect 50456 36416 50520 36420
rect 50536 36476 50600 36480
rect 50536 36420 50540 36476
rect 50540 36420 50596 36476
rect 50596 36420 50600 36476
rect 50536 36416 50600 36420
rect 81016 36476 81080 36480
rect 81016 36420 81020 36476
rect 81020 36420 81076 36476
rect 81076 36420 81080 36476
rect 81016 36416 81080 36420
rect 81096 36476 81160 36480
rect 81096 36420 81100 36476
rect 81100 36420 81156 36476
rect 81156 36420 81160 36476
rect 81096 36416 81160 36420
rect 81176 36476 81240 36480
rect 81176 36420 81180 36476
rect 81180 36420 81236 36476
rect 81236 36420 81240 36476
rect 81176 36416 81240 36420
rect 81256 36476 81320 36480
rect 81256 36420 81260 36476
rect 81260 36420 81316 36476
rect 81316 36420 81320 36476
rect 81256 36416 81320 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 65656 35932 65720 35936
rect 65656 35876 65660 35932
rect 65660 35876 65716 35932
rect 65716 35876 65720 35932
rect 65656 35872 65720 35876
rect 65736 35932 65800 35936
rect 65736 35876 65740 35932
rect 65740 35876 65796 35932
rect 65796 35876 65800 35932
rect 65736 35872 65800 35876
rect 65816 35932 65880 35936
rect 65816 35876 65820 35932
rect 65820 35876 65876 35932
rect 65876 35876 65880 35932
rect 65816 35872 65880 35876
rect 65896 35932 65960 35936
rect 65896 35876 65900 35932
rect 65900 35876 65956 35932
rect 65956 35876 65960 35932
rect 65896 35872 65960 35876
rect 96376 35932 96440 35936
rect 96376 35876 96380 35932
rect 96380 35876 96436 35932
rect 96436 35876 96440 35932
rect 96376 35872 96440 35876
rect 96456 35932 96520 35936
rect 96456 35876 96460 35932
rect 96460 35876 96516 35932
rect 96516 35876 96520 35932
rect 96456 35872 96520 35876
rect 96536 35932 96600 35936
rect 96536 35876 96540 35932
rect 96540 35876 96596 35932
rect 96596 35876 96600 35932
rect 96536 35872 96600 35876
rect 96616 35932 96680 35936
rect 96616 35876 96620 35932
rect 96620 35876 96676 35932
rect 96676 35876 96680 35932
rect 96616 35872 96680 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 50296 35388 50360 35392
rect 50296 35332 50300 35388
rect 50300 35332 50356 35388
rect 50356 35332 50360 35388
rect 50296 35328 50360 35332
rect 50376 35388 50440 35392
rect 50376 35332 50380 35388
rect 50380 35332 50436 35388
rect 50436 35332 50440 35388
rect 50376 35328 50440 35332
rect 50456 35388 50520 35392
rect 50456 35332 50460 35388
rect 50460 35332 50516 35388
rect 50516 35332 50520 35388
rect 50456 35328 50520 35332
rect 50536 35388 50600 35392
rect 50536 35332 50540 35388
rect 50540 35332 50596 35388
rect 50596 35332 50600 35388
rect 50536 35328 50600 35332
rect 81016 35388 81080 35392
rect 81016 35332 81020 35388
rect 81020 35332 81076 35388
rect 81076 35332 81080 35388
rect 81016 35328 81080 35332
rect 81096 35388 81160 35392
rect 81096 35332 81100 35388
rect 81100 35332 81156 35388
rect 81156 35332 81160 35388
rect 81096 35328 81160 35332
rect 81176 35388 81240 35392
rect 81176 35332 81180 35388
rect 81180 35332 81236 35388
rect 81236 35332 81240 35388
rect 81176 35328 81240 35332
rect 81256 35388 81320 35392
rect 81256 35332 81260 35388
rect 81260 35332 81316 35388
rect 81316 35332 81320 35388
rect 81256 35328 81320 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 65656 34844 65720 34848
rect 65656 34788 65660 34844
rect 65660 34788 65716 34844
rect 65716 34788 65720 34844
rect 65656 34784 65720 34788
rect 65736 34844 65800 34848
rect 65736 34788 65740 34844
rect 65740 34788 65796 34844
rect 65796 34788 65800 34844
rect 65736 34784 65800 34788
rect 65816 34844 65880 34848
rect 65816 34788 65820 34844
rect 65820 34788 65876 34844
rect 65876 34788 65880 34844
rect 65816 34784 65880 34788
rect 65896 34844 65960 34848
rect 65896 34788 65900 34844
rect 65900 34788 65956 34844
rect 65956 34788 65960 34844
rect 65896 34784 65960 34788
rect 96376 34844 96440 34848
rect 96376 34788 96380 34844
rect 96380 34788 96436 34844
rect 96436 34788 96440 34844
rect 96376 34784 96440 34788
rect 96456 34844 96520 34848
rect 96456 34788 96460 34844
rect 96460 34788 96516 34844
rect 96516 34788 96520 34844
rect 96456 34784 96520 34788
rect 96536 34844 96600 34848
rect 96536 34788 96540 34844
rect 96540 34788 96596 34844
rect 96596 34788 96600 34844
rect 96536 34784 96600 34788
rect 96616 34844 96680 34848
rect 96616 34788 96620 34844
rect 96620 34788 96676 34844
rect 96676 34788 96680 34844
rect 96616 34784 96680 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 50296 34300 50360 34304
rect 50296 34244 50300 34300
rect 50300 34244 50356 34300
rect 50356 34244 50360 34300
rect 50296 34240 50360 34244
rect 50376 34300 50440 34304
rect 50376 34244 50380 34300
rect 50380 34244 50436 34300
rect 50436 34244 50440 34300
rect 50376 34240 50440 34244
rect 50456 34300 50520 34304
rect 50456 34244 50460 34300
rect 50460 34244 50516 34300
rect 50516 34244 50520 34300
rect 50456 34240 50520 34244
rect 50536 34300 50600 34304
rect 50536 34244 50540 34300
rect 50540 34244 50596 34300
rect 50596 34244 50600 34300
rect 50536 34240 50600 34244
rect 81016 34300 81080 34304
rect 81016 34244 81020 34300
rect 81020 34244 81076 34300
rect 81076 34244 81080 34300
rect 81016 34240 81080 34244
rect 81096 34300 81160 34304
rect 81096 34244 81100 34300
rect 81100 34244 81156 34300
rect 81156 34244 81160 34300
rect 81096 34240 81160 34244
rect 81176 34300 81240 34304
rect 81176 34244 81180 34300
rect 81180 34244 81236 34300
rect 81236 34244 81240 34300
rect 81176 34240 81240 34244
rect 81256 34300 81320 34304
rect 81256 34244 81260 34300
rect 81260 34244 81316 34300
rect 81316 34244 81320 34300
rect 81256 34240 81320 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 65656 33756 65720 33760
rect 65656 33700 65660 33756
rect 65660 33700 65716 33756
rect 65716 33700 65720 33756
rect 65656 33696 65720 33700
rect 65736 33756 65800 33760
rect 65736 33700 65740 33756
rect 65740 33700 65796 33756
rect 65796 33700 65800 33756
rect 65736 33696 65800 33700
rect 65816 33756 65880 33760
rect 65816 33700 65820 33756
rect 65820 33700 65876 33756
rect 65876 33700 65880 33756
rect 65816 33696 65880 33700
rect 65896 33756 65960 33760
rect 65896 33700 65900 33756
rect 65900 33700 65956 33756
rect 65956 33700 65960 33756
rect 65896 33696 65960 33700
rect 96376 33756 96440 33760
rect 96376 33700 96380 33756
rect 96380 33700 96436 33756
rect 96436 33700 96440 33756
rect 96376 33696 96440 33700
rect 96456 33756 96520 33760
rect 96456 33700 96460 33756
rect 96460 33700 96516 33756
rect 96516 33700 96520 33756
rect 96456 33696 96520 33700
rect 96536 33756 96600 33760
rect 96536 33700 96540 33756
rect 96540 33700 96596 33756
rect 96596 33700 96600 33756
rect 96536 33696 96600 33700
rect 96616 33756 96680 33760
rect 96616 33700 96620 33756
rect 96620 33700 96676 33756
rect 96676 33700 96680 33756
rect 96616 33696 96680 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 50296 33212 50360 33216
rect 50296 33156 50300 33212
rect 50300 33156 50356 33212
rect 50356 33156 50360 33212
rect 50296 33152 50360 33156
rect 50376 33212 50440 33216
rect 50376 33156 50380 33212
rect 50380 33156 50436 33212
rect 50436 33156 50440 33212
rect 50376 33152 50440 33156
rect 50456 33212 50520 33216
rect 50456 33156 50460 33212
rect 50460 33156 50516 33212
rect 50516 33156 50520 33212
rect 50456 33152 50520 33156
rect 50536 33212 50600 33216
rect 50536 33156 50540 33212
rect 50540 33156 50596 33212
rect 50596 33156 50600 33212
rect 50536 33152 50600 33156
rect 81016 33212 81080 33216
rect 81016 33156 81020 33212
rect 81020 33156 81076 33212
rect 81076 33156 81080 33212
rect 81016 33152 81080 33156
rect 81096 33212 81160 33216
rect 81096 33156 81100 33212
rect 81100 33156 81156 33212
rect 81156 33156 81160 33212
rect 81096 33152 81160 33156
rect 81176 33212 81240 33216
rect 81176 33156 81180 33212
rect 81180 33156 81236 33212
rect 81236 33156 81240 33212
rect 81176 33152 81240 33156
rect 81256 33212 81320 33216
rect 81256 33156 81260 33212
rect 81260 33156 81316 33212
rect 81316 33156 81320 33212
rect 81256 33152 81320 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 65656 32668 65720 32672
rect 65656 32612 65660 32668
rect 65660 32612 65716 32668
rect 65716 32612 65720 32668
rect 65656 32608 65720 32612
rect 65736 32668 65800 32672
rect 65736 32612 65740 32668
rect 65740 32612 65796 32668
rect 65796 32612 65800 32668
rect 65736 32608 65800 32612
rect 65816 32668 65880 32672
rect 65816 32612 65820 32668
rect 65820 32612 65876 32668
rect 65876 32612 65880 32668
rect 65816 32608 65880 32612
rect 65896 32668 65960 32672
rect 65896 32612 65900 32668
rect 65900 32612 65956 32668
rect 65956 32612 65960 32668
rect 65896 32608 65960 32612
rect 96376 32668 96440 32672
rect 96376 32612 96380 32668
rect 96380 32612 96436 32668
rect 96436 32612 96440 32668
rect 96376 32608 96440 32612
rect 96456 32668 96520 32672
rect 96456 32612 96460 32668
rect 96460 32612 96516 32668
rect 96516 32612 96520 32668
rect 96456 32608 96520 32612
rect 96536 32668 96600 32672
rect 96536 32612 96540 32668
rect 96540 32612 96596 32668
rect 96596 32612 96600 32668
rect 96536 32608 96600 32612
rect 96616 32668 96680 32672
rect 96616 32612 96620 32668
rect 96620 32612 96676 32668
rect 96676 32612 96680 32668
rect 96616 32608 96680 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 50296 32124 50360 32128
rect 50296 32068 50300 32124
rect 50300 32068 50356 32124
rect 50356 32068 50360 32124
rect 50296 32064 50360 32068
rect 50376 32124 50440 32128
rect 50376 32068 50380 32124
rect 50380 32068 50436 32124
rect 50436 32068 50440 32124
rect 50376 32064 50440 32068
rect 50456 32124 50520 32128
rect 50456 32068 50460 32124
rect 50460 32068 50516 32124
rect 50516 32068 50520 32124
rect 50456 32064 50520 32068
rect 50536 32124 50600 32128
rect 50536 32068 50540 32124
rect 50540 32068 50596 32124
rect 50596 32068 50600 32124
rect 50536 32064 50600 32068
rect 81016 32124 81080 32128
rect 81016 32068 81020 32124
rect 81020 32068 81076 32124
rect 81076 32068 81080 32124
rect 81016 32064 81080 32068
rect 81096 32124 81160 32128
rect 81096 32068 81100 32124
rect 81100 32068 81156 32124
rect 81156 32068 81160 32124
rect 81096 32064 81160 32068
rect 81176 32124 81240 32128
rect 81176 32068 81180 32124
rect 81180 32068 81236 32124
rect 81236 32068 81240 32124
rect 81176 32064 81240 32068
rect 81256 32124 81320 32128
rect 81256 32068 81260 32124
rect 81260 32068 81316 32124
rect 81316 32068 81320 32124
rect 81256 32064 81320 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 65656 31580 65720 31584
rect 65656 31524 65660 31580
rect 65660 31524 65716 31580
rect 65716 31524 65720 31580
rect 65656 31520 65720 31524
rect 65736 31580 65800 31584
rect 65736 31524 65740 31580
rect 65740 31524 65796 31580
rect 65796 31524 65800 31580
rect 65736 31520 65800 31524
rect 65816 31580 65880 31584
rect 65816 31524 65820 31580
rect 65820 31524 65876 31580
rect 65876 31524 65880 31580
rect 65816 31520 65880 31524
rect 65896 31580 65960 31584
rect 65896 31524 65900 31580
rect 65900 31524 65956 31580
rect 65956 31524 65960 31580
rect 65896 31520 65960 31524
rect 96376 31580 96440 31584
rect 96376 31524 96380 31580
rect 96380 31524 96436 31580
rect 96436 31524 96440 31580
rect 96376 31520 96440 31524
rect 96456 31580 96520 31584
rect 96456 31524 96460 31580
rect 96460 31524 96516 31580
rect 96516 31524 96520 31580
rect 96456 31520 96520 31524
rect 96536 31580 96600 31584
rect 96536 31524 96540 31580
rect 96540 31524 96596 31580
rect 96596 31524 96600 31580
rect 96536 31520 96600 31524
rect 96616 31580 96680 31584
rect 96616 31524 96620 31580
rect 96620 31524 96676 31580
rect 96676 31524 96680 31580
rect 96616 31520 96680 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 50296 31036 50360 31040
rect 50296 30980 50300 31036
rect 50300 30980 50356 31036
rect 50356 30980 50360 31036
rect 50296 30976 50360 30980
rect 50376 31036 50440 31040
rect 50376 30980 50380 31036
rect 50380 30980 50436 31036
rect 50436 30980 50440 31036
rect 50376 30976 50440 30980
rect 50456 31036 50520 31040
rect 50456 30980 50460 31036
rect 50460 30980 50516 31036
rect 50516 30980 50520 31036
rect 50456 30976 50520 30980
rect 50536 31036 50600 31040
rect 50536 30980 50540 31036
rect 50540 30980 50596 31036
rect 50596 30980 50600 31036
rect 50536 30976 50600 30980
rect 81016 31036 81080 31040
rect 81016 30980 81020 31036
rect 81020 30980 81076 31036
rect 81076 30980 81080 31036
rect 81016 30976 81080 30980
rect 81096 31036 81160 31040
rect 81096 30980 81100 31036
rect 81100 30980 81156 31036
rect 81156 30980 81160 31036
rect 81096 30976 81160 30980
rect 81176 31036 81240 31040
rect 81176 30980 81180 31036
rect 81180 30980 81236 31036
rect 81236 30980 81240 31036
rect 81176 30976 81240 30980
rect 81256 31036 81320 31040
rect 81256 30980 81260 31036
rect 81260 30980 81316 31036
rect 81316 30980 81320 31036
rect 81256 30976 81320 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 65656 30492 65720 30496
rect 65656 30436 65660 30492
rect 65660 30436 65716 30492
rect 65716 30436 65720 30492
rect 65656 30432 65720 30436
rect 65736 30492 65800 30496
rect 65736 30436 65740 30492
rect 65740 30436 65796 30492
rect 65796 30436 65800 30492
rect 65736 30432 65800 30436
rect 65816 30492 65880 30496
rect 65816 30436 65820 30492
rect 65820 30436 65876 30492
rect 65876 30436 65880 30492
rect 65816 30432 65880 30436
rect 65896 30492 65960 30496
rect 65896 30436 65900 30492
rect 65900 30436 65956 30492
rect 65956 30436 65960 30492
rect 65896 30432 65960 30436
rect 96376 30492 96440 30496
rect 96376 30436 96380 30492
rect 96380 30436 96436 30492
rect 96436 30436 96440 30492
rect 96376 30432 96440 30436
rect 96456 30492 96520 30496
rect 96456 30436 96460 30492
rect 96460 30436 96516 30492
rect 96516 30436 96520 30492
rect 96456 30432 96520 30436
rect 96536 30492 96600 30496
rect 96536 30436 96540 30492
rect 96540 30436 96596 30492
rect 96596 30436 96600 30492
rect 96536 30432 96600 30436
rect 96616 30492 96680 30496
rect 96616 30436 96620 30492
rect 96620 30436 96676 30492
rect 96676 30436 96680 30492
rect 96616 30432 96680 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 50296 29948 50360 29952
rect 50296 29892 50300 29948
rect 50300 29892 50356 29948
rect 50356 29892 50360 29948
rect 50296 29888 50360 29892
rect 50376 29948 50440 29952
rect 50376 29892 50380 29948
rect 50380 29892 50436 29948
rect 50436 29892 50440 29948
rect 50376 29888 50440 29892
rect 50456 29948 50520 29952
rect 50456 29892 50460 29948
rect 50460 29892 50516 29948
rect 50516 29892 50520 29948
rect 50456 29888 50520 29892
rect 50536 29948 50600 29952
rect 50536 29892 50540 29948
rect 50540 29892 50596 29948
rect 50596 29892 50600 29948
rect 50536 29888 50600 29892
rect 81016 29948 81080 29952
rect 81016 29892 81020 29948
rect 81020 29892 81076 29948
rect 81076 29892 81080 29948
rect 81016 29888 81080 29892
rect 81096 29948 81160 29952
rect 81096 29892 81100 29948
rect 81100 29892 81156 29948
rect 81156 29892 81160 29948
rect 81096 29888 81160 29892
rect 81176 29948 81240 29952
rect 81176 29892 81180 29948
rect 81180 29892 81236 29948
rect 81236 29892 81240 29948
rect 81176 29888 81240 29892
rect 81256 29948 81320 29952
rect 81256 29892 81260 29948
rect 81260 29892 81316 29948
rect 81316 29892 81320 29948
rect 81256 29888 81320 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 65656 29404 65720 29408
rect 65656 29348 65660 29404
rect 65660 29348 65716 29404
rect 65716 29348 65720 29404
rect 65656 29344 65720 29348
rect 65736 29404 65800 29408
rect 65736 29348 65740 29404
rect 65740 29348 65796 29404
rect 65796 29348 65800 29404
rect 65736 29344 65800 29348
rect 65816 29404 65880 29408
rect 65816 29348 65820 29404
rect 65820 29348 65876 29404
rect 65876 29348 65880 29404
rect 65816 29344 65880 29348
rect 65896 29404 65960 29408
rect 65896 29348 65900 29404
rect 65900 29348 65956 29404
rect 65956 29348 65960 29404
rect 65896 29344 65960 29348
rect 96376 29404 96440 29408
rect 96376 29348 96380 29404
rect 96380 29348 96436 29404
rect 96436 29348 96440 29404
rect 96376 29344 96440 29348
rect 96456 29404 96520 29408
rect 96456 29348 96460 29404
rect 96460 29348 96516 29404
rect 96516 29348 96520 29404
rect 96456 29344 96520 29348
rect 96536 29404 96600 29408
rect 96536 29348 96540 29404
rect 96540 29348 96596 29404
rect 96596 29348 96600 29404
rect 96536 29344 96600 29348
rect 96616 29404 96680 29408
rect 96616 29348 96620 29404
rect 96620 29348 96676 29404
rect 96676 29348 96680 29404
rect 96616 29344 96680 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 50296 28860 50360 28864
rect 50296 28804 50300 28860
rect 50300 28804 50356 28860
rect 50356 28804 50360 28860
rect 50296 28800 50360 28804
rect 50376 28860 50440 28864
rect 50376 28804 50380 28860
rect 50380 28804 50436 28860
rect 50436 28804 50440 28860
rect 50376 28800 50440 28804
rect 50456 28860 50520 28864
rect 50456 28804 50460 28860
rect 50460 28804 50516 28860
rect 50516 28804 50520 28860
rect 50456 28800 50520 28804
rect 50536 28860 50600 28864
rect 50536 28804 50540 28860
rect 50540 28804 50596 28860
rect 50596 28804 50600 28860
rect 50536 28800 50600 28804
rect 81016 28860 81080 28864
rect 81016 28804 81020 28860
rect 81020 28804 81076 28860
rect 81076 28804 81080 28860
rect 81016 28800 81080 28804
rect 81096 28860 81160 28864
rect 81096 28804 81100 28860
rect 81100 28804 81156 28860
rect 81156 28804 81160 28860
rect 81096 28800 81160 28804
rect 81176 28860 81240 28864
rect 81176 28804 81180 28860
rect 81180 28804 81236 28860
rect 81236 28804 81240 28860
rect 81176 28800 81240 28804
rect 81256 28860 81320 28864
rect 81256 28804 81260 28860
rect 81260 28804 81316 28860
rect 81316 28804 81320 28860
rect 81256 28800 81320 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 65656 28316 65720 28320
rect 65656 28260 65660 28316
rect 65660 28260 65716 28316
rect 65716 28260 65720 28316
rect 65656 28256 65720 28260
rect 65736 28316 65800 28320
rect 65736 28260 65740 28316
rect 65740 28260 65796 28316
rect 65796 28260 65800 28316
rect 65736 28256 65800 28260
rect 65816 28316 65880 28320
rect 65816 28260 65820 28316
rect 65820 28260 65876 28316
rect 65876 28260 65880 28316
rect 65816 28256 65880 28260
rect 65896 28316 65960 28320
rect 65896 28260 65900 28316
rect 65900 28260 65956 28316
rect 65956 28260 65960 28316
rect 65896 28256 65960 28260
rect 96376 28316 96440 28320
rect 96376 28260 96380 28316
rect 96380 28260 96436 28316
rect 96436 28260 96440 28316
rect 96376 28256 96440 28260
rect 96456 28316 96520 28320
rect 96456 28260 96460 28316
rect 96460 28260 96516 28316
rect 96516 28260 96520 28316
rect 96456 28256 96520 28260
rect 96536 28316 96600 28320
rect 96536 28260 96540 28316
rect 96540 28260 96596 28316
rect 96596 28260 96600 28316
rect 96536 28256 96600 28260
rect 96616 28316 96680 28320
rect 96616 28260 96620 28316
rect 96620 28260 96676 28316
rect 96676 28260 96680 28316
rect 96616 28256 96680 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 50296 27772 50360 27776
rect 50296 27716 50300 27772
rect 50300 27716 50356 27772
rect 50356 27716 50360 27772
rect 50296 27712 50360 27716
rect 50376 27772 50440 27776
rect 50376 27716 50380 27772
rect 50380 27716 50436 27772
rect 50436 27716 50440 27772
rect 50376 27712 50440 27716
rect 50456 27772 50520 27776
rect 50456 27716 50460 27772
rect 50460 27716 50516 27772
rect 50516 27716 50520 27772
rect 50456 27712 50520 27716
rect 50536 27772 50600 27776
rect 50536 27716 50540 27772
rect 50540 27716 50596 27772
rect 50596 27716 50600 27772
rect 50536 27712 50600 27716
rect 81016 27772 81080 27776
rect 81016 27716 81020 27772
rect 81020 27716 81076 27772
rect 81076 27716 81080 27772
rect 81016 27712 81080 27716
rect 81096 27772 81160 27776
rect 81096 27716 81100 27772
rect 81100 27716 81156 27772
rect 81156 27716 81160 27772
rect 81096 27712 81160 27716
rect 81176 27772 81240 27776
rect 81176 27716 81180 27772
rect 81180 27716 81236 27772
rect 81236 27716 81240 27772
rect 81176 27712 81240 27716
rect 81256 27772 81320 27776
rect 81256 27716 81260 27772
rect 81260 27716 81316 27772
rect 81316 27716 81320 27772
rect 81256 27712 81320 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 65656 27228 65720 27232
rect 65656 27172 65660 27228
rect 65660 27172 65716 27228
rect 65716 27172 65720 27228
rect 65656 27168 65720 27172
rect 65736 27228 65800 27232
rect 65736 27172 65740 27228
rect 65740 27172 65796 27228
rect 65796 27172 65800 27228
rect 65736 27168 65800 27172
rect 65816 27228 65880 27232
rect 65816 27172 65820 27228
rect 65820 27172 65876 27228
rect 65876 27172 65880 27228
rect 65816 27168 65880 27172
rect 65896 27228 65960 27232
rect 65896 27172 65900 27228
rect 65900 27172 65956 27228
rect 65956 27172 65960 27228
rect 65896 27168 65960 27172
rect 96376 27228 96440 27232
rect 96376 27172 96380 27228
rect 96380 27172 96436 27228
rect 96436 27172 96440 27228
rect 96376 27168 96440 27172
rect 96456 27228 96520 27232
rect 96456 27172 96460 27228
rect 96460 27172 96516 27228
rect 96516 27172 96520 27228
rect 96456 27168 96520 27172
rect 96536 27228 96600 27232
rect 96536 27172 96540 27228
rect 96540 27172 96596 27228
rect 96596 27172 96600 27228
rect 96536 27168 96600 27172
rect 96616 27228 96680 27232
rect 96616 27172 96620 27228
rect 96620 27172 96676 27228
rect 96676 27172 96680 27228
rect 96616 27168 96680 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 50296 26684 50360 26688
rect 50296 26628 50300 26684
rect 50300 26628 50356 26684
rect 50356 26628 50360 26684
rect 50296 26624 50360 26628
rect 50376 26684 50440 26688
rect 50376 26628 50380 26684
rect 50380 26628 50436 26684
rect 50436 26628 50440 26684
rect 50376 26624 50440 26628
rect 50456 26684 50520 26688
rect 50456 26628 50460 26684
rect 50460 26628 50516 26684
rect 50516 26628 50520 26684
rect 50456 26624 50520 26628
rect 50536 26684 50600 26688
rect 50536 26628 50540 26684
rect 50540 26628 50596 26684
rect 50596 26628 50600 26684
rect 50536 26624 50600 26628
rect 81016 26684 81080 26688
rect 81016 26628 81020 26684
rect 81020 26628 81076 26684
rect 81076 26628 81080 26684
rect 81016 26624 81080 26628
rect 81096 26684 81160 26688
rect 81096 26628 81100 26684
rect 81100 26628 81156 26684
rect 81156 26628 81160 26684
rect 81096 26624 81160 26628
rect 81176 26684 81240 26688
rect 81176 26628 81180 26684
rect 81180 26628 81236 26684
rect 81236 26628 81240 26684
rect 81176 26624 81240 26628
rect 81256 26684 81320 26688
rect 81256 26628 81260 26684
rect 81260 26628 81316 26684
rect 81316 26628 81320 26684
rect 81256 26624 81320 26628
rect 38516 26556 38580 26620
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 65656 26140 65720 26144
rect 65656 26084 65660 26140
rect 65660 26084 65716 26140
rect 65716 26084 65720 26140
rect 65656 26080 65720 26084
rect 65736 26140 65800 26144
rect 65736 26084 65740 26140
rect 65740 26084 65796 26140
rect 65796 26084 65800 26140
rect 65736 26080 65800 26084
rect 65816 26140 65880 26144
rect 65816 26084 65820 26140
rect 65820 26084 65876 26140
rect 65876 26084 65880 26140
rect 65816 26080 65880 26084
rect 65896 26140 65960 26144
rect 65896 26084 65900 26140
rect 65900 26084 65956 26140
rect 65956 26084 65960 26140
rect 65896 26080 65960 26084
rect 96376 26140 96440 26144
rect 96376 26084 96380 26140
rect 96380 26084 96436 26140
rect 96436 26084 96440 26140
rect 96376 26080 96440 26084
rect 96456 26140 96520 26144
rect 96456 26084 96460 26140
rect 96460 26084 96516 26140
rect 96516 26084 96520 26140
rect 96456 26080 96520 26084
rect 96536 26140 96600 26144
rect 96536 26084 96540 26140
rect 96540 26084 96596 26140
rect 96596 26084 96600 26140
rect 96536 26080 96600 26084
rect 96616 26140 96680 26144
rect 96616 26084 96620 26140
rect 96620 26084 96676 26140
rect 96676 26084 96680 26140
rect 96616 26080 96680 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 50296 25596 50360 25600
rect 50296 25540 50300 25596
rect 50300 25540 50356 25596
rect 50356 25540 50360 25596
rect 50296 25536 50360 25540
rect 50376 25596 50440 25600
rect 50376 25540 50380 25596
rect 50380 25540 50436 25596
rect 50436 25540 50440 25596
rect 50376 25536 50440 25540
rect 50456 25596 50520 25600
rect 50456 25540 50460 25596
rect 50460 25540 50516 25596
rect 50516 25540 50520 25596
rect 50456 25536 50520 25540
rect 50536 25596 50600 25600
rect 50536 25540 50540 25596
rect 50540 25540 50596 25596
rect 50596 25540 50600 25596
rect 50536 25536 50600 25540
rect 81016 25596 81080 25600
rect 81016 25540 81020 25596
rect 81020 25540 81076 25596
rect 81076 25540 81080 25596
rect 81016 25536 81080 25540
rect 81096 25596 81160 25600
rect 81096 25540 81100 25596
rect 81100 25540 81156 25596
rect 81156 25540 81160 25596
rect 81096 25536 81160 25540
rect 81176 25596 81240 25600
rect 81176 25540 81180 25596
rect 81180 25540 81236 25596
rect 81236 25540 81240 25596
rect 81176 25536 81240 25540
rect 81256 25596 81320 25600
rect 81256 25540 81260 25596
rect 81260 25540 81316 25596
rect 81316 25540 81320 25596
rect 81256 25536 81320 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 65656 25052 65720 25056
rect 65656 24996 65660 25052
rect 65660 24996 65716 25052
rect 65716 24996 65720 25052
rect 65656 24992 65720 24996
rect 65736 25052 65800 25056
rect 65736 24996 65740 25052
rect 65740 24996 65796 25052
rect 65796 24996 65800 25052
rect 65736 24992 65800 24996
rect 65816 25052 65880 25056
rect 65816 24996 65820 25052
rect 65820 24996 65876 25052
rect 65876 24996 65880 25052
rect 65816 24992 65880 24996
rect 65896 25052 65960 25056
rect 65896 24996 65900 25052
rect 65900 24996 65956 25052
rect 65956 24996 65960 25052
rect 65896 24992 65960 24996
rect 96376 25052 96440 25056
rect 96376 24996 96380 25052
rect 96380 24996 96436 25052
rect 96436 24996 96440 25052
rect 96376 24992 96440 24996
rect 96456 25052 96520 25056
rect 96456 24996 96460 25052
rect 96460 24996 96516 25052
rect 96516 24996 96520 25052
rect 96456 24992 96520 24996
rect 96536 25052 96600 25056
rect 96536 24996 96540 25052
rect 96540 24996 96596 25052
rect 96596 24996 96600 25052
rect 96536 24992 96600 24996
rect 96616 25052 96680 25056
rect 96616 24996 96620 25052
rect 96620 24996 96676 25052
rect 96676 24996 96680 25052
rect 96616 24992 96680 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 50296 24508 50360 24512
rect 50296 24452 50300 24508
rect 50300 24452 50356 24508
rect 50356 24452 50360 24508
rect 50296 24448 50360 24452
rect 50376 24508 50440 24512
rect 50376 24452 50380 24508
rect 50380 24452 50436 24508
rect 50436 24452 50440 24508
rect 50376 24448 50440 24452
rect 50456 24508 50520 24512
rect 50456 24452 50460 24508
rect 50460 24452 50516 24508
rect 50516 24452 50520 24508
rect 50456 24448 50520 24452
rect 50536 24508 50600 24512
rect 50536 24452 50540 24508
rect 50540 24452 50596 24508
rect 50596 24452 50600 24508
rect 50536 24448 50600 24452
rect 81016 24508 81080 24512
rect 81016 24452 81020 24508
rect 81020 24452 81076 24508
rect 81076 24452 81080 24508
rect 81016 24448 81080 24452
rect 81096 24508 81160 24512
rect 81096 24452 81100 24508
rect 81100 24452 81156 24508
rect 81156 24452 81160 24508
rect 81096 24448 81160 24452
rect 81176 24508 81240 24512
rect 81176 24452 81180 24508
rect 81180 24452 81236 24508
rect 81236 24452 81240 24508
rect 81176 24448 81240 24452
rect 81256 24508 81320 24512
rect 81256 24452 81260 24508
rect 81260 24452 81316 24508
rect 81316 24452 81320 24508
rect 81256 24448 81320 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 65656 23964 65720 23968
rect 65656 23908 65660 23964
rect 65660 23908 65716 23964
rect 65716 23908 65720 23964
rect 65656 23904 65720 23908
rect 65736 23964 65800 23968
rect 65736 23908 65740 23964
rect 65740 23908 65796 23964
rect 65796 23908 65800 23964
rect 65736 23904 65800 23908
rect 65816 23964 65880 23968
rect 65816 23908 65820 23964
rect 65820 23908 65876 23964
rect 65876 23908 65880 23964
rect 65816 23904 65880 23908
rect 65896 23964 65960 23968
rect 65896 23908 65900 23964
rect 65900 23908 65956 23964
rect 65956 23908 65960 23964
rect 65896 23904 65960 23908
rect 96376 23964 96440 23968
rect 96376 23908 96380 23964
rect 96380 23908 96436 23964
rect 96436 23908 96440 23964
rect 96376 23904 96440 23908
rect 96456 23964 96520 23968
rect 96456 23908 96460 23964
rect 96460 23908 96516 23964
rect 96516 23908 96520 23964
rect 96456 23904 96520 23908
rect 96536 23964 96600 23968
rect 96536 23908 96540 23964
rect 96540 23908 96596 23964
rect 96596 23908 96600 23964
rect 96536 23904 96600 23908
rect 96616 23964 96680 23968
rect 96616 23908 96620 23964
rect 96620 23908 96676 23964
rect 96676 23908 96680 23964
rect 96616 23904 96680 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 50296 23420 50360 23424
rect 50296 23364 50300 23420
rect 50300 23364 50356 23420
rect 50356 23364 50360 23420
rect 50296 23360 50360 23364
rect 50376 23420 50440 23424
rect 50376 23364 50380 23420
rect 50380 23364 50436 23420
rect 50436 23364 50440 23420
rect 50376 23360 50440 23364
rect 50456 23420 50520 23424
rect 50456 23364 50460 23420
rect 50460 23364 50516 23420
rect 50516 23364 50520 23420
rect 50456 23360 50520 23364
rect 50536 23420 50600 23424
rect 50536 23364 50540 23420
rect 50540 23364 50596 23420
rect 50596 23364 50600 23420
rect 50536 23360 50600 23364
rect 81016 23420 81080 23424
rect 81016 23364 81020 23420
rect 81020 23364 81076 23420
rect 81076 23364 81080 23420
rect 81016 23360 81080 23364
rect 81096 23420 81160 23424
rect 81096 23364 81100 23420
rect 81100 23364 81156 23420
rect 81156 23364 81160 23420
rect 81096 23360 81160 23364
rect 81176 23420 81240 23424
rect 81176 23364 81180 23420
rect 81180 23364 81236 23420
rect 81236 23364 81240 23420
rect 81176 23360 81240 23364
rect 81256 23420 81320 23424
rect 81256 23364 81260 23420
rect 81260 23364 81316 23420
rect 81316 23364 81320 23420
rect 81256 23360 81320 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 65656 22876 65720 22880
rect 65656 22820 65660 22876
rect 65660 22820 65716 22876
rect 65716 22820 65720 22876
rect 65656 22816 65720 22820
rect 65736 22876 65800 22880
rect 65736 22820 65740 22876
rect 65740 22820 65796 22876
rect 65796 22820 65800 22876
rect 65736 22816 65800 22820
rect 65816 22876 65880 22880
rect 65816 22820 65820 22876
rect 65820 22820 65876 22876
rect 65876 22820 65880 22876
rect 65816 22816 65880 22820
rect 65896 22876 65960 22880
rect 65896 22820 65900 22876
rect 65900 22820 65956 22876
rect 65956 22820 65960 22876
rect 65896 22816 65960 22820
rect 96376 22876 96440 22880
rect 96376 22820 96380 22876
rect 96380 22820 96436 22876
rect 96436 22820 96440 22876
rect 96376 22816 96440 22820
rect 96456 22876 96520 22880
rect 96456 22820 96460 22876
rect 96460 22820 96516 22876
rect 96516 22820 96520 22876
rect 96456 22816 96520 22820
rect 96536 22876 96600 22880
rect 96536 22820 96540 22876
rect 96540 22820 96596 22876
rect 96596 22820 96600 22876
rect 96536 22816 96600 22820
rect 96616 22876 96680 22880
rect 96616 22820 96620 22876
rect 96620 22820 96676 22876
rect 96676 22820 96680 22876
rect 96616 22816 96680 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 50296 22332 50360 22336
rect 50296 22276 50300 22332
rect 50300 22276 50356 22332
rect 50356 22276 50360 22332
rect 50296 22272 50360 22276
rect 50376 22332 50440 22336
rect 50376 22276 50380 22332
rect 50380 22276 50436 22332
rect 50436 22276 50440 22332
rect 50376 22272 50440 22276
rect 50456 22332 50520 22336
rect 50456 22276 50460 22332
rect 50460 22276 50516 22332
rect 50516 22276 50520 22332
rect 50456 22272 50520 22276
rect 50536 22332 50600 22336
rect 50536 22276 50540 22332
rect 50540 22276 50596 22332
rect 50596 22276 50600 22332
rect 50536 22272 50600 22276
rect 81016 22332 81080 22336
rect 81016 22276 81020 22332
rect 81020 22276 81076 22332
rect 81076 22276 81080 22332
rect 81016 22272 81080 22276
rect 81096 22332 81160 22336
rect 81096 22276 81100 22332
rect 81100 22276 81156 22332
rect 81156 22276 81160 22332
rect 81096 22272 81160 22276
rect 81176 22332 81240 22336
rect 81176 22276 81180 22332
rect 81180 22276 81236 22332
rect 81236 22276 81240 22332
rect 81176 22272 81240 22276
rect 81256 22332 81320 22336
rect 81256 22276 81260 22332
rect 81260 22276 81316 22332
rect 81316 22276 81320 22332
rect 81256 22272 81320 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 65656 21788 65720 21792
rect 65656 21732 65660 21788
rect 65660 21732 65716 21788
rect 65716 21732 65720 21788
rect 65656 21728 65720 21732
rect 65736 21788 65800 21792
rect 65736 21732 65740 21788
rect 65740 21732 65796 21788
rect 65796 21732 65800 21788
rect 65736 21728 65800 21732
rect 65816 21788 65880 21792
rect 65816 21732 65820 21788
rect 65820 21732 65876 21788
rect 65876 21732 65880 21788
rect 65816 21728 65880 21732
rect 65896 21788 65960 21792
rect 65896 21732 65900 21788
rect 65900 21732 65956 21788
rect 65956 21732 65960 21788
rect 65896 21728 65960 21732
rect 96376 21788 96440 21792
rect 96376 21732 96380 21788
rect 96380 21732 96436 21788
rect 96436 21732 96440 21788
rect 96376 21728 96440 21732
rect 96456 21788 96520 21792
rect 96456 21732 96460 21788
rect 96460 21732 96516 21788
rect 96516 21732 96520 21788
rect 96456 21728 96520 21732
rect 96536 21788 96600 21792
rect 96536 21732 96540 21788
rect 96540 21732 96596 21788
rect 96596 21732 96600 21788
rect 96536 21728 96600 21732
rect 96616 21788 96680 21792
rect 96616 21732 96620 21788
rect 96620 21732 96676 21788
rect 96676 21732 96680 21788
rect 96616 21728 96680 21732
rect 38516 21584 38580 21588
rect 38516 21528 38566 21584
rect 38566 21528 38580 21584
rect 38516 21524 38580 21528
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 50296 21244 50360 21248
rect 50296 21188 50300 21244
rect 50300 21188 50356 21244
rect 50356 21188 50360 21244
rect 50296 21184 50360 21188
rect 50376 21244 50440 21248
rect 50376 21188 50380 21244
rect 50380 21188 50436 21244
rect 50436 21188 50440 21244
rect 50376 21184 50440 21188
rect 50456 21244 50520 21248
rect 50456 21188 50460 21244
rect 50460 21188 50516 21244
rect 50516 21188 50520 21244
rect 50456 21184 50520 21188
rect 50536 21244 50600 21248
rect 50536 21188 50540 21244
rect 50540 21188 50596 21244
rect 50596 21188 50600 21244
rect 50536 21184 50600 21188
rect 81016 21244 81080 21248
rect 81016 21188 81020 21244
rect 81020 21188 81076 21244
rect 81076 21188 81080 21244
rect 81016 21184 81080 21188
rect 81096 21244 81160 21248
rect 81096 21188 81100 21244
rect 81100 21188 81156 21244
rect 81156 21188 81160 21244
rect 81096 21184 81160 21188
rect 81176 21244 81240 21248
rect 81176 21188 81180 21244
rect 81180 21188 81236 21244
rect 81236 21188 81240 21244
rect 81176 21184 81240 21188
rect 81256 21244 81320 21248
rect 81256 21188 81260 21244
rect 81260 21188 81316 21244
rect 81316 21188 81320 21244
rect 81256 21184 81320 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 65656 20700 65720 20704
rect 65656 20644 65660 20700
rect 65660 20644 65716 20700
rect 65716 20644 65720 20700
rect 65656 20640 65720 20644
rect 65736 20700 65800 20704
rect 65736 20644 65740 20700
rect 65740 20644 65796 20700
rect 65796 20644 65800 20700
rect 65736 20640 65800 20644
rect 65816 20700 65880 20704
rect 65816 20644 65820 20700
rect 65820 20644 65876 20700
rect 65876 20644 65880 20700
rect 65816 20640 65880 20644
rect 65896 20700 65960 20704
rect 65896 20644 65900 20700
rect 65900 20644 65956 20700
rect 65956 20644 65960 20700
rect 65896 20640 65960 20644
rect 96376 20700 96440 20704
rect 96376 20644 96380 20700
rect 96380 20644 96436 20700
rect 96436 20644 96440 20700
rect 96376 20640 96440 20644
rect 96456 20700 96520 20704
rect 96456 20644 96460 20700
rect 96460 20644 96516 20700
rect 96516 20644 96520 20700
rect 96456 20640 96520 20644
rect 96536 20700 96600 20704
rect 96536 20644 96540 20700
rect 96540 20644 96596 20700
rect 96596 20644 96600 20700
rect 96536 20640 96600 20644
rect 96616 20700 96680 20704
rect 96616 20644 96620 20700
rect 96620 20644 96676 20700
rect 96676 20644 96680 20700
rect 96616 20640 96680 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 50296 20156 50360 20160
rect 50296 20100 50300 20156
rect 50300 20100 50356 20156
rect 50356 20100 50360 20156
rect 50296 20096 50360 20100
rect 50376 20156 50440 20160
rect 50376 20100 50380 20156
rect 50380 20100 50436 20156
rect 50436 20100 50440 20156
rect 50376 20096 50440 20100
rect 50456 20156 50520 20160
rect 50456 20100 50460 20156
rect 50460 20100 50516 20156
rect 50516 20100 50520 20156
rect 50456 20096 50520 20100
rect 50536 20156 50600 20160
rect 50536 20100 50540 20156
rect 50540 20100 50596 20156
rect 50596 20100 50600 20156
rect 50536 20096 50600 20100
rect 81016 20156 81080 20160
rect 81016 20100 81020 20156
rect 81020 20100 81076 20156
rect 81076 20100 81080 20156
rect 81016 20096 81080 20100
rect 81096 20156 81160 20160
rect 81096 20100 81100 20156
rect 81100 20100 81156 20156
rect 81156 20100 81160 20156
rect 81096 20096 81160 20100
rect 81176 20156 81240 20160
rect 81176 20100 81180 20156
rect 81180 20100 81236 20156
rect 81236 20100 81240 20156
rect 81176 20096 81240 20100
rect 81256 20156 81320 20160
rect 81256 20100 81260 20156
rect 81260 20100 81316 20156
rect 81316 20100 81320 20156
rect 81256 20096 81320 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 65656 19612 65720 19616
rect 65656 19556 65660 19612
rect 65660 19556 65716 19612
rect 65716 19556 65720 19612
rect 65656 19552 65720 19556
rect 65736 19612 65800 19616
rect 65736 19556 65740 19612
rect 65740 19556 65796 19612
rect 65796 19556 65800 19612
rect 65736 19552 65800 19556
rect 65816 19612 65880 19616
rect 65816 19556 65820 19612
rect 65820 19556 65876 19612
rect 65876 19556 65880 19612
rect 65816 19552 65880 19556
rect 65896 19612 65960 19616
rect 65896 19556 65900 19612
rect 65900 19556 65956 19612
rect 65956 19556 65960 19612
rect 65896 19552 65960 19556
rect 96376 19612 96440 19616
rect 96376 19556 96380 19612
rect 96380 19556 96436 19612
rect 96436 19556 96440 19612
rect 96376 19552 96440 19556
rect 96456 19612 96520 19616
rect 96456 19556 96460 19612
rect 96460 19556 96516 19612
rect 96516 19556 96520 19612
rect 96456 19552 96520 19556
rect 96536 19612 96600 19616
rect 96536 19556 96540 19612
rect 96540 19556 96596 19612
rect 96596 19556 96600 19612
rect 96536 19552 96600 19556
rect 96616 19612 96680 19616
rect 96616 19556 96620 19612
rect 96620 19556 96676 19612
rect 96676 19556 96680 19612
rect 96616 19552 96680 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 50296 19068 50360 19072
rect 50296 19012 50300 19068
rect 50300 19012 50356 19068
rect 50356 19012 50360 19068
rect 50296 19008 50360 19012
rect 50376 19068 50440 19072
rect 50376 19012 50380 19068
rect 50380 19012 50436 19068
rect 50436 19012 50440 19068
rect 50376 19008 50440 19012
rect 50456 19068 50520 19072
rect 50456 19012 50460 19068
rect 50460 19012 50516 19068
rect 50516 19012 50520 19068
rect 50456 19008 50520 19012
rect 50536 19068 50600 19072
rect 50536 19012 50540 19068
rect 50540 19012 50596 19068
rect 50596 19012 50600 19068
rect 50536 19008 50600 19012
rect 81016 19068 81080 19072
rect 81016 19012 81020 19068
rect 81020 19012 81076 19068
rect 81076 19012 81080 19068
rect 81016 19008 81080 19012
rect 81096 19068 81160 19072
rect 81096 19012 81100 19068
rect 81100 19012 81156 19068
rect 81156 19012 81160 19068
rect 81096 19008 81160 19012
rect 81176 19068 81240 19072
rect 81176 19012 81180 19068
rect 81180 19012 81236 19068
rect 81236 19012 81240 19068
rect 81176 19008 81240 19012
rect 81256 19068 81320 19072
rect 81256 19012 81260 19068
rect 81260 19012 81316 19068
rect 81316 19012 81320 19068
rect 81256 19008 81320 19012
rect 38516 18804 38580 18868
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 65656 18524 65720 18528
rect 65656 18468 65660 18524
rect 65660 18468 65716 18524
rect 65716 18468 65720 18524
rect 65656 18464 65720 18468
rect 65736 18524 65800 18528
rect 65736 18468 65740 18524
rect 65740 18468 65796 18524
rect 65796 18468 65800 18524
rect 65736 18464 65800 18468
rect 65816 18524 65880 18528
rect 65816 18468 65820 18524
rect 65820 18468 65876 18524
rect 65876 18468 65880 18524
rect 65816 18464 65880 18468
rect 65896 18524 65960 18528
rect 65896 18468 65900 18524
rect 65900 18468 65956 18524
rect 65956 18468 65960 18524
rect 65896 18464 65960 18468
rect 96376 18524 96440 18528
rect 96376 18468 96380 18524
rect 96380 18468 96436 18524
rect 96436 18468 96440 18524
rect 96376 18464 96440 18468
rect 96456 18524 96520 18528
rect 96456 18468 96460 18524
rect 96460 18468 96516 18524
rect 96516 18468 96520 18524
rect 96456 18464 96520 18468
rect 96536 18524 96600 18528
rect 96536 18468 96540 18524
rect 96540 18468 96596 18524
rect 96596 18468 96600 18524
rect 96536 18464 96600 18468
rect 96616 18524 96680 18528
rect 96616 18468 96620 18524
rect 96620 18468 96676 18524
rect 96676 18468 96680 18524
rect 96616 18464 96680 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 50296 17980 50360 17984
rect 50296 17924 50300 17980
rect 50300 17924 50356 17980
rect 50356 17924 50360 17980
rect 50296 17920 50360 17924
rect 50376 17980 50440 17984
rect 50376 17924 50380 17980
rect 50380 17924 50436 17980
rect 50436 17924 50440 17980
rect 50376 17920 50440 17924
rect 50456 17980 50520 17984
rect 50456 17924 50460 17980
rect 50460 17924 50516 17980
rect 50516 17924 50520 17980
rect 50456 17920 50520 17924
rect 50536 17980 50600 17984
rect 50536 17924 50540 17980
rect 50540 17924 50596 17980
rect 50596 17924 50600 17980
rect 50536 17920 50600 17924
rect 81016 17980 81080 17984
rect 81016 17924 81020 17980
rect 81020 17924 81076 17980
rect 81076 17924 81080 17980
rect 81016 17920 81080 17924
rect 81096 17980 81160 17984
rect 81096 17924 81100 17980
rect 81100 17924 81156 17980
rect 81156 17924 81160 17980
rect 81096 17920 81160 17924
rect 81176 17980 81240 17984
rect 81176 17924 81180 17980
rect 81180 17924 81236 17980
rect 81236 17924 81240 17980
rect 81176 17920 81240 17924
rect 81256 17980 81320 17984
rect 81256 17924 81260 17980
rect 81260 17924 81316 17980
rect 81316 17924 81320 17980
rect 81256 17920 81320 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 65656 17436 65720 17440
rect 65656 17380 65660 17436
rect 65660 17380 65716 17436
rect 65716 17380 65720 17436
rect 65656 17376 65720 17380
rect 65736 17436 65800 17440
rect 65736 17380 65740 17436
rect 65740 17380 65796 17436
rect 65796 17380 65800 17436
rect 65736 17376 65800 17380
rect 65816 17436 65880 17440
rect 65816 17380 65820 17436
rect 65820 17380 65876 17436
rect 65876 17380 65880 17436
rect 65816 17376 65880 17380
rect 65896 17436 65960 17440
rect 65896 17380 65900 17436
rect 65900 17380 65956 17436
rect 65956 17380 65960 17436
rect 65896 17376 65960 17380
rect 96376 17436 96440 17440
rect 96376 17380 96380 17436
rect 96380 17380 96436 17436
rect 96436 17380 96440 17436
rect 96376 17376 96440 17380
rect 96456 17436 96520 17440
rect 96456 17380 96460 17436
rect 96460 17380 96516 17436
rect 96516 17380 96520 17436
rect 96456 17376 96520 17380
rect 96536 17436 96600 17440
rect 96536 17380 96540 17436
rect 96540 17380 96596 17436
rect 96596 17380 96600 17436
rect 96536 17376 96600 17380
rect 96616 17436 96680 17440
rect 96616 17380 96620 17436
rect 96620 17380 96676 17436
rect 96676 17380 96680 17436
rect 96616 17376 96680 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 50296 16892 50360 16896
rect 50296 16836 50300 16892
rect 50300 16836 50356 16892
rect 50356 16836 50360 16892
rect 50296 16832 50360 16836
rect 50376 16892 50440 16896
rect 50376 16836 50380 16892
rect 50380 16836 50436 16892
rect 50436 16836 50440 16892
rect 50376 16832 50440 16836
rect 50456 16892 50520 16896
rect 50456 16836 50460 16892
rect 50460 16836 50516 16892
rect 50516 16836 50520 16892
rect 50456 16832 50520 16836
rect 50536 16892 50600 16896
rect 50536 16836 50540 16892
rect 50540 16836 50596 16892
rect 50596 16836 50600 16892
rect 50536 16832 50600 16836
rect 81016 16892 81080 16896
rect 81016 16836 81020 16892
rect 81020 16836 81076 16892
rect 81076 16836 81080 16892
rect 81016 16832 81080 16836
rect 81096 16892 81160 16896
rect 81096 16836 81100 16892
rect 81100 16836 81156 16892
rect 81156 16836 81160 16892
rect 81096 16832 81160 16836
rect 81176 16892 81240 16896
rect 81176 16836 81180 16892
rect 81180 16836 81236 16892
rect 81236 16836 81240 16892
rect 81176 16832 81240 16836
rect 81256 16892 81320 16896
rect 81256 16836 81260 16892
rect 81260 16836 81316 16892
rect 81316 16836 81320 16892
rect 81256 16832 81320 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 65656 16348 65720 16352
rect 65656 16292 65660 16348
rect 65660 16292 65716 16348
rect 65716 16292 65720 16348
rect 65656 16288 65720 16292
rect 65736 16348 65800 16352
rect 65736 16292 65740 16348
rect 65740 16292 65796 16348
rect 65796 16292 65800 16348
rect 65736 16288 65800 16292
rect 65816 16348 65880 16352
rect 65816 16292 65820 16348
rect 65820 16292 65876 16348
rect 65876 16292 65880 16348
rect 65816 16288 65880 16292
rect 65896 16348 65960 16352
rect 65896 16292 65900 16348
rect 65900 16292 65956 16348
rect 65956 16292 65960 16348
rect 65896 16288 65960 16292
rect 96376 16348 96440 16352
rect 96376 16292 96380 16348
rect 96380 16292 96436 16348
rect 96436 16292 96440 16348
rect 96376 16288 96440 16292
rect 96456 16348 96520 16352
rect 96456 16292 96460 16348
rect 96460 16292 96516 16348
rect 96516 16292 96520 16348
rect 96456 16288 96520 16292
rect 96536 16348 96600 16352
rect 96536 16292 96540 16348
rect 96540 16292 96596 16348
rect 96596 16292 96600 16348
rect 96536 16288 96600 16292
rect 96616 16348 96680 16352
rect 96616 16292 96620 16348
rect 96620 16292 96676 16348
rect 96676 16292 96680 16348
rect 96616 16288 96680 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 50296 15804 50360 15808
rect 50296 15748 50300 15804
rect 50300 15748 50356 15804
rect 50356 15748 50360 15804
rect 50296 15744 50360 15748
rect 50376 15804 50440 15808
rect 50376 15748 50380 15804
rect 50380 15748 50436 15804
rect 50436 15748 50440 15804
rect 50376 15744 50440 15748
rect 50456 15804 50520 15808
rect 50456 15748 50460 15804
rect 50460 15748 50516 15804
rect 50516 15748 50520 15804
rect 50456 15744 50520 15748
rect 50536 15804 50600 15808
rect 50536 15748 50540 15804
rect 50540 15748 50596 15804
rect 50596 15748 50600 15804
rect 50536 15744 50600 15748
rect 81016 15804 81080 15808
rect 81016 15748 81020 15804
rect 81020 15748 81076 15804
rect 81076 15748 81080 15804
rect 81016 15744 81080 15748
rect 81096 15804 81160 15808
rect 81096 15748 81100 15804
rect 81100 15748 81156 15804
rect 81156 15748 81160 15804
rect 81096 15744 81160 15748
rect 81176 15804 81240 15808
rect 81176 15748 81180 15804
rect 81180 15748 81236 15804
rect 81236 15748 81240 15804
rect 81176 15744 81240 15748
rect 81256 15804 81320 15808
rect 81256 15748 81260 15804
rect 81260 15748 81316 15804
rect 81316 15748 81320 15804
rect 81256 15744 81320 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 65656 15260 65720 15264
rect 65656 15204 65660 15260
rect 65660 15204 65716 15260
rect 65716 15204 65720 15260
rect 65656 15200 65720 15204
rect 65736 15260 65800 15264
rect 65736 15204 65740 15260
rect 65740 15204 65796 15260
rect 65796 15204 65800 15260
rect 65736 15200 65800 15204
rect 65816 15260 65880 15264
rect 65816 15204 65820 15260
rect 65820 15204 65876 15260
rect 65876 15204 65880 15260
rect 65816 15200 65880 15204
rect 65896 15260 65960 15264
rect 65896 15204 65900 15260
rect 65900 15204 65956 15260
rect 65956 15204 65960 15260
rect 65896 15200 65960 15204
rect 96376 15260 96440 15264
rect 96376 15204 96380 15260
rect 96380 15204 96436 15260
rect 96436 15204 96440 15260
rect 96376 15200 96440 15204
rect 96456 15260 96520 15264
rect 96456 15204 96460 15260
rect 96460 15204 96516 15260
rect 96516 15204 96520 15260
rect 96456 15200 96520 15204
rect 96536 15260 96600 15264
rect 96536 15204 96540 15260
rect 96540 15204 96596 15260
rect 96596 15204 96600 15260
rect 96536 15200 96600 15204
rect 96616 15260 96680 15264
rect 96616 15204 96620 15260
rect 96620 15204 96676 15260
rect 96676 15204 96680 15260
rect 96616 15200 96680 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 50296 14716 50360 14720
rect 50296 14660 50300 14716
rect 50300 14660 50356 14716
rect 50356 14660 50360 14716
rect 50296 14656 50360 14660
rect 50376 14716 50440 14720
rect 50376 14660 50380 14716
rect 50380 14660 50436 14716
rect 50436 14660 50440 14716
rect 50376 14656 50440 14660
rect 50456 14716 50520 14720
rect 50456 14660 50460 14716
rect 50460 14660 50516 14716
rect 50516 14660 50520 14716
rect 50456 14656 50520 14660
rect 50536 14716 50600 14720
rect 50536 14660 50540 14716
rect 50540 14660 50596 14716
rect 50596 14660 50600 14716
rect 50536 14656 50600 14660
rect 81016 14716 81080 14720
rect 81016 14660 81020 14716
rect 81020 14660 81076 14716
rect 81076 14660 81080 14716
rect 81016 14656 81080 14660
rect 81096 14716 81160 14720
rect 81096 14660 81100 14716
rect 81100 14660 81156 14716
rect 81156 14660 81160 14716
rect 81096 14656 81160 14660
rect 81176 14716 81240 14720
rect 81176 14660 81180 14716
rect 81180 14660 81236 14716
rect 81236 14660 81240 14716
rect 81176 14656 81240 14660
rect 81256 14716 81320 14720
rect 81256 14660 81260 14716
rect 81260 14660 81316 14716
rect 81316 14660 81320 14716
rect 81256 14656 81320 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 65656 14172 65720 14176
rect 65656 14116 65660 14172
rect 65660 14116 65716 14172
rect 65716 14116 65720 14172
rect 65656 14112 65720 14116
rect 65736 14172 65800 14176
rect 65736 14116 65740 14172
rect 65740 14116 65796 14172
rect 65796 14116 65800 14172
rect 65736 14112 65800 14116
rect 65816 14172 65880 14176
rect 65816 14116 65820 14172
rect 65820 14116 65876 14172
rect 65876 14116 65880 14172
rect 65816 14112 65880 14116
rect 65896 14172 65960 14176
rect 65896 14116 65900 14172
rect 65900 14116 65956 14172
rect 65956 14116 65960 14172
rect 65896 14112 65960 14116
rect 96376 14172 96440 14176
rect 96376 14116 96380 14172
rect 96380 14116 96436 14172
rect 96436 14116 96440 14172
rect 96376 14112 96440 14116
rect 96456 14172 96520 14176
rect 96456 14116 96460 14172
rect 96460 14116 96516 14172
rect 96516 14116 96520 14172
rect 96456 14112 96520 14116
rect 96536 14172 96600 14176
rect 96536 14116 96540 14172
rect 96540 14116 96596 14172
rect 96596 14116 96600 14172
rect 96536 14112 96600 14116
rect 96616 14172 96680 14176
rect 96616 14116 96620 14172
rect 96620 14116 96676 14172
rect 96676 14116 96680 14172
rect 96616 14112 96680 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 50296 13628 50360 13632
rect 50296 13572 50300 13628
rect 50300 13572 50356 13628
rect 50356 13572 50360 13628
rect 50296 13568 50360 13572
rect 50376 13628 50440 13632
rect 50376 13572 50380 13628
rect 50380 13572 50436 13628
rect 50436 13572 50440 13628
rect 50376 13568 50440 13572
rect 50456 13628 50520 13632
rect 50456 13572 50460 13628
rect 50460 13572 50516 13628
rect 50516 13572 50520 13628
rect 50456 13568 50520 13572
rect 50536 13628 50600 13632
rect 50536 13572 50540 13628
rect 50540 13572 50596 13628
rect 50596 13572 50600 13628
rect 50536 13568 50600 13572
rect 81016 13628 81080 13632
rect 81016 13572 81020 13628
rect 81020 13572 81076 13628
rect 81076 13572 81080 13628
rect 81016 13568 81080 13572
rect 81096 13628 81160 13632
rect 81096 13572 81100 13628
rect 81100 13572 81156 13628
rect 81156 13572 81160 13628
rect 81096 13568 81160 13572
rect 81176 13628 81240 13632
rect 81176 13572 81180 13628
rect 81180 13572 81236 13628
rect 81236 13572 81240 13628
rect 81176 13568 81240 13572
rect 81256 13628 81320 13632
rect 81256 13572 81260 13628
rect 81260 13572 81316 13628
rect 81316 13572 81320 13628
rect 81256 13568 81320 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 65656 13084 65720 13088
rect 65656 13028 65660 13084
rect 65660 13028 65716 13084
rect 65716 13028 65720 13084
rect 65656 13024 65720 13028
rect 65736 13084 65800 13088
rect 65736 13028 65740 13084
rect 65740 13028 65796 13084
rect 65796 13028 65800 13084
rect 65736 13024 65800 13028
rect 65816 13084 65880 13088
rect 65816 13028 65820 13084
rect 65820 13028 65876 13084
rect 65876 13028 65880 13084
rect 65816 13024 65880 13028
rect 65896 13084 65960 13088
rect 65896 13028 65900 13084
rect 65900 13028 65956 13084
rect 65956 13028 65960 13084
rect 65896 13024 65960 13028
rect 96376 13084 96440 13088
rect 96376 13028 96380 13084
rect 96380 13028 96436 13084
rect 96436 13028 96440 13084
rect 96376 13024 96440 13028
rect 96456 13084 96520 13088
rect 96456 13028 96460 13084
rect 96460 13028 96516 13084
rect 96516 13028 96520 13084
rect 96456 13024 96520 13028
rect 96536 13084 96600 13088
rect 96536 13028 96540 13084
rect 96540 13028 96596 13084
rect 96596 13028 96600 13084
rect 96536 13024 96600 13028
rect 96616 13084 96680 13088
rect 96616 13028 96620 13084
rect 96620 13028 96676 13084
rect 96676 13028 96680 13084
rect 96616 13024 96680 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 50296 12540 50360 12544
rect 50296 12484 50300 12540
rect 50300 12484 50356 12540
rect 50356 12484 50360 12540
rect 50296 12480 50360 12484
rect 50376 12540 50440 12544
rect 50376 12484 50380 12540
rect 50380 12484 50436 12540
rect 50436 12484 50440 12540
rect 50376 12480 50440 12484
rect 50456 12540 50520 12544
rect 50456 12484 50460 12540
rect 50460 12484 50516 12540
rect 50516 12484 50520 12540
rect 50456 12480 50520 12484
rect 50536 12540 50600 12544
rect 50536 12484 50540 12540
rect 50540 12484 50596 12540
rect 50596 12484 50600 12540
rect 50536 12480 50600 12484
rect 81016 12540 81080 12544
rect 81016 12484 81020 12540
rect 81020 12484 81076 12540
rect 81076 12484 81080 12540
rect 81016 12480 81080 12484
rect 81096 12540 81160 12544
rect 81096 12484 81100 12540
rect 81100 12484 81156 12540
rect 81156 12484 81160 12540
rect 81096 12480 81160 12484
rect 81176 12540 81240 12544
rect 81176 12484 81180 12540
rect 81180 12484 81236 12540
rect 81236 12484 81240 12540
rect 81176 12480 81240 12484
rect 81256 12540 81320 12544
rect 81256 12484 81260 12540
rect 81260 12484 81316 12540
rect 81316 12484 81320 12540
rect 81256 12480 81320 12484
rect 38700 12336 38764 12340
rect 38700 12280 38714 12336
rect 38714 12280 38764 12336
rect 38700 12276 38764 12280
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 65656 11996 65720 12000
rect 65656 11940 65660 11996
rect 65660 11940 65716 11996
rect 65716 11940 65720 11996
rect 65656 11936 65720 11940
rect 65736 11996 65800 12000
rect 65736 11940 65740 11996
rect 65740 11940 65796 11996
rect 65796 11940 65800 11996
rect 65736 11936 65800 11940
rect 65816 11996 65880 12000
rect 65816 11940 65820 11996
rect 65820 11940 65876 11996
rect 65876 11940 65880 11996
rect 65816 11936 65880 11940
rect 65896 11996 65960 12000
rect 65896 11940 65900 11996
rect 65900 11940 65956 11996
rect 65956 11940 65960 11996
rect 65896 11936 65960 11940
rect 96376 11996 96440 12000
rect 96376 11940 96380 11996
rect 96380 11940 96436 11996
rect 96436 11940 96440 11996
rect 96376 11936 96440 11940
rect 96456 11996 96520 12000
rect 96456 11940 96460 11996
rect 96460 11940 96516 11996
rect 96516 11940 96520 11996
rect 96456 11936 96520 11940
rect 96536 11996 96600 12000
rect 96536 11940 96540 11996
rect 96540 11940 96596 11996
rect 96596 11940 96600 11996
rect 96536 11936 96600 11940
rect 96616 11996 96680 12000
rect 96616 11940 96620 11996
rect 96620 11940 96676 11996
rect 96676 11940 96680 11996
rect 96616 11936 96680 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 50296 11452 50360 11456
rect 50296 11396 50300 11452
rect 50300 11396 50356 11452
rect 50356 11396 50360 11452
rect 50296 11392 50360 11396
rect 50376 11452 50440 11456
rect 50376 11396 50380 11452
rect 50380 11396 50436 11452
rect 50436 11396 50440 11452
rect 50376 11392 50440 11396
rect 50456 11452 50520 11456
rect 50456 11396 50460 11452
rect 50460 11396 50516 11452
rect 50516 11396 50520 11452
rect 50456 11392 50520 11396
rect 50536 11452 50600 11456
rect 50536 11396 50540 11452
rect 50540 11396 50596 11452
rect 50596 11396 50600 11452
rect 50536 11392 50600 11396
rect 81016 11452 81080 11456
rect 81016 11396 81020 11452
rect 81020 11396 81076 11452
rect 81076 11396 81080 11452
rect 81016 11392 81080 11396
rect 81096 11452 81160 11456
rect 81096 11396 81100 11452
rect 81100 11396 81156 11452
rect 81156 11396 81160 11452
rect 81096 11392 81160 11396
rect 81176 11452 81240 11456
rect 81176 11396 81180 11452
rect 81180 11396 81236 11452
rect 81236 11396 81240 11452
rect 81176 11392 81240 11396
rect 81256 11452 81320 11456
rect 81256 11396 81260 11452
rect 81260 11396 81316 11452
rect 81316 11396 81320 11452
rect 81256 11392 81320 11396
rect 38516 11384 38580 11388
rect 38516 11328 38530 11384
rect 38530 11328 38580 11384
rect 38516 11324 38580 11328
rect 38700 11112 38764 11116
rect 38700 11056 38750 11112
rect 38750 11056 38764 11112
rect 38700 11052 38764 11056
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 65656 10908 65720 10912
rect 65656 10852 65660 10908
rect 65660 10852 65716 10908
rect 65716 10852 65720 10908
rect 65656 10848 65720 10852
rect 65736 10908 65800 10912
rect 65736 10852 65740 10908
rect 65740 10852 65796 10908
rect 65796 10852 65800 10908
rect 65736 10848 65800 10852
rect 65816 10908 65880 10912
rect 65816 10852 65820 10908
rect 65820 10852 65876 10908
rect 65876 10852 65880 10908
rect 65816 10848 65880 10852
rect 65896 10908 65960 10912
rect 65896 10852 65900 10908
rect 65900 10852 65956 10908
rect 65956 10852 65960 10908
rect 65896 10848 65960 10852
rect 96376 10908 96440 10912
rect 96376 10852 96380 10908
rect 96380 10852 96436 10908
rect 96436 10852 96440 10908
rect 96376 10848 96440 10852
rect 96456 10908 96520 10912
rect 96456 10852 96460 10908
rect 96460 10852 96516 10908
rect 96516 10852 96520 10908
rect 96456 10848 96520 10852
rect 96536 10908 96600 10912
rect 96536 10852 96540 10908
rect 96540 10852 96596 10908
rect 96596 10852 96600 10908
rect 96536 10848 96600 10852
rect 96616 10908 96680 10912
rect 96616 10852 96620 10908
rect 96620 10852 96676 10908
rect 96676 10852 96680 10908
rect 96616 10848 96680 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 50296 10364 50360 10368
rect 50296 10308 50300 10364
rect 50300 10308 50356 10364
rect 50356 10308 50360 10364
rect 50296 10304 50360 10308
rect 50376 10364 50440 10368
rect 50376 10308 50380 10364
rect 50380 10308 50436 10364
rect 50436 10308 50440 10364
rect 50376 10304 50440 10308
rect 50456 10364 50520 10368
rect 50456 10308 50460 10364
rect 50460 10308 50516 10364
rect 50516 10308 50520 10364
rect 50456 10304 50520 10308
rect 50536 10364 50600 10368
rect 50536 10308 50540 10364
rect 50540 10308 50596 10364
rect 50596 10308 50600 10364
rect 50536 10304 50600 10308
rect 81016 10364 81080 10368
rect 81016 10308 81020 10364
rect 81020 10308 81076 10364
rect 81076 10308 81080 10364
rect 81016 10304 81080 10308
rect 81096 10364 81160 10368
rect 81096 10308 81100 10364
rect 81100 10308 81156 10364
rect 81156 10308 81160 10364
rect 81096 10304 81160 10308
rect 81176 10364 81240 10368
rect 81176 10308 81180 10364
rect 81180 10308 81236 10364
rect 81236 10308 81240 10364
rect 81176 10304 81240 10308
rect 81256 10364 81320 10368
rect 81256 10308 81260 10364
rect 81260 10308 81316 10364
rect 81316 10308 81320 10364
rect 81256 10304 81320 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 65656 9820 65720 9824
rect 65656 9764 65660 9820
rect 65660 9764 65716 9820
rect 65716 9764 65720 9820
rect 65656 9760 65720 9764
rect 65736 9820 65800 9824
rect 65736 9764 65740 9820
rect 65740 9764 65796 9820
rect 65796 9764 65800 9820
rect 65736 9760 65800 9764
rect 65816 9820 65880 9824
rect 65816 9764 65820 9820
rect 65820 9764 65876 9820
rect 65876 9764 65880 9820
rect 65816 9760 65880 9764
rect 65896 9820 65960 9824
rect 65896 9764 65900 9820
rect 65900 9764 65956 9820
rect 65956 9764 65960 9820
rect 65896 9760 65960 9764
rect 96376 9820 96440 9824
rect 96376 9764 96380 9820
rect 96380 9764 96436 9820
rect 96436 9764 96440 9820
rect 96376 9760 96440 9764
rect 96456 9820 96520 9824
rect 96456 9764 96460 9820
rect 96460 9764 96516 9820
rect 96516 9764 96520 9820
rect 96456 9760 96520 9764
rect 96536 9820 96600 9824
rect 96536 9764 96540 9820
rect 96540 9764 96596 9820
rect 96596 9764 96600 9820
rect 96536 9760 96600 9764
rect 96616 9820 96680 9824
rect 96616 9764 96620 9820
rect 96620 9764 96676 9820
rect 96676 9764 96680 9820
rect 96616 9760 96680 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 50296 9276 50360 9280
rect 50296 9220 50300 9276
rect 50300 9220 50356 9276
rect 50356 9220 50360 9276
rect 50296 9216 50360 9220
rect 50376 9276 50440 9280
rect 50376 9220 50380 9276
rect 50380 9220 50436 9276
rect 50436 9220 50440 9276
rect 50376 9216 50440 9220
rect 50456 9276 50520 9280
rect 50456 9220 50460 9276
rect 50460 9220 50516 9276
rect 50516 9220 50520 9276
rect 50456 9216 50520 9220
rect 50536 9276 50600 9280
rect 50536 9220 50540 9276
rect 50540 9220 50596 9276
rect 50596 9220 50600 9276
rect 50536 9216 50600 9220
rect 81016 9276 81080 9280
rect 81016 9220 81020 9276
rect 81020 9220 81076 9276
rect 81076 9220 81080 9276
rect 81016 9216 81080 9220
rect 81096 9276 81160 9280
rect 81096 9220 81100 9276
rect 81100 9220 81156 9276
rect 81156 9220 81160 9276
rect 81096 9216 81160 9220
rect 81176 9276 81240 9280
rect 81176 9220 81180 9276
rect 81180 9220 81236 9276
rect 81236 9220 81240 9276
rect 81176 9216 81240 9220
rect 81256 9276 81320 9280
rect 81256 9220 81260 9276
rect 81260 9220 81316 9276
rect 81316 9220 81320 9276
rect 81256 9216 81320 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 65656 8732 65720 8736
rect 65656 8676 65660 8732
rect 65660 8676 65716 8732
rect 65716 8676 65720 8732
rect 65656 8672 65720 8676
rect 65736 8732 65800 8736
rect 65736 8676 65740 8732
rect 65740 8676 65796 8732
rect 65796 8676 65800 8732
rect 65736 8672 65800 8676
rect 65816 8732 65880 8736
rect 65816 8676 65820 8732
rect 65820 8676 65876 8732
rect 65876 8676 65880 8732
rect 65816 8672 65880 8676
rect 65896 8732 65960 8736
rect 65896 8676 65900 8732
rect 65900 8676 65956 8732
rect 65956 8676 65960 8732
rect 65896 8672 65960 8676
rect 96376 8732 96440 8736
rect 96376 8676 96380 8732
rect 96380 8676 96436 8732
rect 96436 8676 96440 8732
rect 96376 8672 96440 8676
rect 96456 8732 96520 8736
rect 96456 8676 96460 8732
rect 96460 8676 96516 8732
rect 96516 8676 96520 8732
rect 96456 8672 96520 8676
rect 96536 8732 96600 8736
rect 96536 8676 96540 8732
rect 96540 8676 96596 8732
rect 96596 8676 96600 8732
rect 96536 8672 96600 8676
rect 96616 8732 96680 8736
rect 96616 8676 96620 8732
rect 96620 8676 96676 8732
rect 96676 8676 96680 8732
rect 96616 8672 96680 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 50296 8188 50360 8192
rect 50296 8132 50300 8188
rect 50300 8132 50356 8188
rect 50356 8132 50360 8188
rect 50296 8128 50360 8132
rect 50376 8188 50440 8192
rect 50376 8132 50380 8188
rect 50380 8132 50436 8188
rect 50436 8132 50440 8188
rect 50376 8128 50440 8132
rect 50456 8188 50520 8192
rect 50456 8132 50460 8188
rect 50460 8132 50516 8188
rect 50516 8132 50520 8188
rect 50456 8128 50520 8132
rect 50536 8188 50600 8192
rect 50536 8132 50540 8188
rect 50540 8132 50596 8188
rect 50596 8132 50600 8188
rect 50536 8128 50600 8132
rect 81016 8188 81080 8192
rect 81016 8132 81020 8188
rect 81020 8132 81076 8188
rect 81076 8132 81080 8188
rect 81016 8128 81080 8132
rect 81096 8188 81160 8192
rect 81096 8132 81100 8188
rect 81100 8132 81156 8188
rect 81156 8132 81160 8188
rect 81096 8128 81160 8132
rect 81176 8188 81240 8192
rect 81176 8132 81180 8188
rect 81180 8132 81236 8188
rect 81236 8132 81240 8188
rect 81176 8128 81240 8132
rect 81256 8188 81320 8192
rect 81256 8132 81260 8188
rect 81260 8132 81316 8188
rect 81316 8132 81320 8188
rect 81256 8128 81320 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 65656 7644 65720 7648
rect 65656 7588 65660 7644
rect 65660 7588 65716 7644
rect 65716 7588 65720 7644
rect 65656 7584 65720 7588
rect 65736 7644 65800 7648
rect 65736 7588 65740 7644
rect 65740 7588 65796 7644
rect 65796 7588 65800 7644
rect 65736 7584 65800 7588
rect 65816 7644 65880 7648
rect 65816 7588 65820 7644
rect 65820 7588 65876 7644
rect 65876 7588 65880 7644
rect 65816 7584 65880 7588
rect 65896 7644 65960 7648
rect 65896 7588 65900 7644
rect 65900 7588 65956 7644
rect 65956 7588 65960 7644
rect 65896 7584 65960 7588
rect 96376 7644 96440 7648
rect 96376 7588 96380 7644
rect 96380 7588 96436 7644
rect 96436 7588 96440 7644
rect 96376 7584 96440 7588
rect 96456 7644 96520 7648
rect 96456 7588 96460 7644
rect 96460 7588 96516 7644
rect 96516 7588 96520 7644
rect 96456 7584 96520 7588
rect 96536 7644 96600 7648
rect 96536 7588 96540 7644
rect 96540 7588 96596 7644
rect 96596 7588 96600 7644
rect 96536 7584 96600 7588
rect 96616 7644 96680 7648
rect 96616 7588 96620 7644
rect 96620 7588 96676 7644
rect 96676 7588 96680 7644
rect 96616 7584 96680 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 50296 7100 50360 7104
rect 50296 7044 50300 7100
rect 50300 7044 50356 7100
rect 50356 7044 50360 7100
rect 50296 7040 50360 7044
rect 50376 7100 50440 7104
rect 50376 7044 50380 7100
rect 50380 7044 50436 7100
rect 50436 7044 50440 7100
rect 50376 7040 50440 7044
rect 50456 7100 50520 7104
rect 50456 7044 50460 7100
rect 50460 7044 50516 7100
rect 50516 7044 50520 7100
rect 50456 7040 50520 7044
rect 50536 7100 50600 7104
rect 50536 7044 50540 7100
rect 50540 7044 50596 7100
rect 50596 7044 50600 7100
rect 50536 7040 50600 7044
rect 81016 7100 81080 7104
rect 81016 7044 81020 7100
rect 81020 7044 81076 7100
rect 81076 7044 81080 7100
rect 81016 7040 81080 7044
rect 81096 7100 81160 7104
rect 81096 7044 81100 7100
rect 81100 7044 81156 7100
rect 81156 7044 81160 7100
rect 81096 7040 81160 7044
rect 81176 7100 81240 7104
rect 81176 7044 81180 7100
rect 81180 7044 81236 7100
rect 81236 7044 81240 7100
rect 81176 7040 81240 7044
rect 81256 7100 81320 7104
rect 81256 7044 81260 7100
rect 81260 7044 81316 7100
rect 81316 7044 81320 7100
rect 81256 7040 81320 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 65656 6556 65720 6560
rect 65656 6500 65660 6556
rect 65660 6500 65716 6556
rect 65716 6500 65720 6556
rect 65656 6496 65720 6500
rect 65736 6556 65800 6560
rect 65736 6500 65740 6556
rect 65740 6500 65796 6556
rect 65796 6500 65800 6556
rect 65736 6496 65800 6500
rect 65816 6556 65880 6560
rect 65816 6500 65820 6556
rect 65820 6500 65876 6556
rect 65876 6500 65880 6556
rect 65816 6496 65880 6500
rect 65896 6556 65960 6560
rect 65896 6500 65900 6556
rect 65900 6500 65956 6556
rect 65956 6500 65960 6556
rect 65896 6496 65960 6500
rect 96376 6556 96440 6560
rect 96376 6500 96380 6556
rect 96380 6500 96436 6556
rect 96436 6500 96440 6556
rect 96376 6496 96440 6500
rect 96456 6556 96520 6560
rect 96456 6500 96460 6556
rect 96460 6500 96516 6556
rect 96516 6500 96520 6556
rect 96456 6496 96520 6500
rect 96536 6556 96600 6560
rect 96536 6500 96540 6556
rect 96540 6500 96596 6556
rect 96596 6500 96600 6556
rect 96536 6496 96600 6500
rect 96616 6556 96680 6560
rect 96616 6500 96620 6556
rect 96620 6500 96676 6556
rect 96676 6500 96680 6556
rect 96616 6496 96680 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 50296 6012 50360 6016
rect 50296 5956 50300 6012
rect 50300 5956 50356 6012
rect 50356 5956 50360 6012
rect 50296 5952 50360 5956
rect 50376 6012 50440 6016
rect 50376 5956 50380 6012
rect 50380 5956 50436 6012
rect 50436 5956 50440 6012
rect 50376 5952 50440 5956
rect 50456 6012 50520 6016
rect 50456 5956 50460 6012
rect 50460 5956 50516 6012
rect 50516 5956 50520 6012
rect 50456 5952 50520 5956
rect 50536 6012 50600 6016
rect 50536 5956 50540 6012
rect 50540 5956 50596 6012
rect 50596 5956 50600 6012
rect 50536 5952 50600 5956
rect 81016 6012 81080 6016
rect 81016 5956 81020 6012
rect 81020 5956 81076 6012
rect 81076 5956 81080 6012
rect 81016 5952 81080 5956
rect 81096 6012 81160 6016
rect 81096 5956 81100 6012
rect 81100 5956 81156 6012
rect 81156 5956 81160 6012
rect 81096 5952 81160 5956
rect 81176 6012 81240 6016
rect 81176 5956 81180 6012
rect 81180 5956 81236 6012
rect 81236 5956 81240 6012
rect 81176 5952 81240 5956
rect 81256 6012 81320 6016
rect 81256 5956 81260 6012
rect 81260 5956 81316 6012
rect 81316 5956 81320 6012
rect 81256 5952 81320 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 65656 5468 65720 5472
rect 65656 5412 65660 5468
rect 65660 5412 65716 5468
rect 65716 5412 65720 5468
rect 65656 5408 65720 5412
rect 65736 5468 65800 5472
rect 65736 5412 65740 5468
rect 65740 5412 65796 5468
rect 65796 5412 65800 5468
rect 65736 5408 65800 5412
rect 65816 5468 65880 5472
rect 65816 5412 65820 5468
rect 65820 5412 65876 5468
rect 65876 5412 65880 5468
rect 65816 5408 65880 5412
rect 65896 5468 65960 5472
rect 65896 5412 65900 5468
rect 65900 5412 65956 5468
rect 65956 5412 65960 5468
rect 65896 5408 65960 5412
rect 96376 5468 96440 5472
rect 96376 5412 96380 5468
rect 96380 5412 96436 5468
rect 96436 5412 96440 5468
rect 96376 5408 96440 5412
rect 96456 5468 96520 5472
rect 96456 5412 96460 5468
rect 96460 5412 96516 5468
rect 96516 5412 96520 5468
rect 96456 5408 96520 5412
rect 96536 5468 96600 5472
rect 96536 5412 96540 5468
rect 96540 5412 96596 5468
rect 96596 5412 96600 5468
rect 96536 5408 96600 5412
rect 96616 5468 96680 5472
rect 96616 5412 96620 5468
rect 96620 5412 96676 5468
rect 96676 5412 96680 5468
rect 96616 5408 96680 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 50296 4924 50360 4928
rect 50296 4868 50300 4924
rect 50300 4868 50356 4924
rect 50356 4868 50360 4924
rect 50296 4864 50360 4868
rect 50376 4924 50440 4928
rect 50376 4868 50380 4924
rect 50380 4868 50436 4924
rect 50436 4868 50440 4924
rect 50376 4864 50440 4868
rect 50456 4924 50520 4928
rect 50456 4868 50460 4924
rect 50460 4868 50516 4924
rect 50516 4868 50520 4924
rect 50456 4864 50520 4868
rect 50536 4924 50600 4928
rect 50536 4868 50540 4924
rect 50540 4868 50596 4924
rect 50596 4868 50600 4924
rect 50536 4864 50600 4868
rect 81016 4924 81080 4928
rect 81016 4868 81020 4924
rect 81020 4868 81076 4924
rect 81076 4868 81080 4924
rect 81016 4864 81080 4868
rect 81096 4924 81160 4928
rect 81096 4868 81100 4924
rect 81100 4868 81156 4924
rect 81156 4868 81160 4924
rect 81096 4864 81160 4868
rect 81176 4924 81240 4928
rect 81176 4868 81180 4924
rect 81180 4868 81236 4924
rect 81236 4868 81240 4924
rect 81176 4864 81240 4868
rect 81256 4924 81320 4928
rect 81256 4868 81260 4924
rect 81260 4868 81316 4924
rect 81316 4868 81320 4924
rect 81256 4864 81320 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 65656 4380 65720 4384
rect 65656 4324 65660 4380
rect 65660 4324 65716 4380
rect 65716 4324 65720 4380
rect 65656 4320 65720 4324
rect 65736 4380 65800 4384
rect 65736 4324 65740 4380
rect 65740 4324 65796 4380
rect 65796 4324 65800 4380
rect 65736 4320 65800 4324
rect 65816 4380 65880 4384
rect 65816 4324 65820 4380
rect 65820 4324 65876 4380
rect 65876 4324 65880 4380
rect 65816 4320 65880 4324
rect 65896 4380 65960 4384
rect 65896 4324 65900 4380
rect 65900 4324 65956 4380
rect 65956 4324 65960 4380
rect 65896 4320 65960 4324
rect 96376 4380 96440 4384
rect 96376 4324 96380 4380
rect 96380 4324 96436 4380
rect 96436 4324 96440 4380
rect 96376 4320 96440 4324
rect 96456 4380 96520 4384
rect 96456 4324 96460 4380
rect 96460 4324 96516 4380
rect 96516 4324 96520 4380
rect 96456 4320 96520 4324
rect 96536 4380 96600 4384
rect 96536 4324 96540 4380
rect 96540 4324 96596 4380
rect 96596 4324 96600 4380
rect 96536 4320 96600 4324
rect 96616 4380 96680 4384
rect 96616 4324 96620 4380
rect 96620 4324 96676 4380
rect 96676 4324 96680 4380
rect 96616 4320 96680 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 50296 3836 50360 3840
rect 50296 3780 50300 3836
rect 50300 3780 50356 3836
rect 50356 3780 50360 3836
rect 50296 3776 50360 3780
rect 50376 3836 50440 3840
rect 50376 3780 50380 3836
rect 50380 3780 50436 3836
rect 50436 3780 50440 3836
rect 50376 3776 50440 3780
rect 50456 3836 50520 3840
rect 50456 3780 50460 3836
rect 50460 3780 50516 3836
rect 50516 3780 50520 3836
rect 50456 3776 50520 3780
rect 50536 3836 50600 3840
rect 50536 3780 50540 3836
rect 50540 3780 50596 3836
rect 50596 3780 50600 3836
rect 50536 3776 50600 3780
rect 81016 3836 81080 3840
rect 81016 3780 81020 3836
rect 81020 3780 81076 3836
rect 81076 3780 81080 3836
rect 81016 3776 81080 3780
rect 81096 3836 81160 3840
rect 81096 3780 81100 3836
rect 81100 3780 81156 3836
rect 81156 3780 81160 3836
rect 81096 3776 81160 3780
rect 81176 3836 81240 3840
rect 81176 3780 81180 3836
rect 81180 3780 81236 3836
rect 81236 3780 81240 3836
rect 81176 3776 81240 3780
rect 81256 3836 81320 3840
rect 81256 3780 81260 3836
rect 81260 3780 81316 3836
rect 81316 3780 81320 3836
rect 81256 3776 81320 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 65656 3292 65720 3296
rect 65656 3236 65660 3292
rect 65660 3236 65716 3292
rect 65716 3236 65720 3292
rect 65656 3232 65720 3236
rect 65736 3292 65800 3296
rect 65736 3236 65740 3292
rect 65740 3236 65796 3292
rect 65796 3236 65800 3292
rect 65736 3232 65800 3236
rect 65816 3292 65880 3296
rect 65816 3236 65820 3292
rect 65820 3236 65876 3292
rect 65876 3236 65880 3292
rect 65816 3232 65880 3236
rect 65896 3292 65960 3296
rect 65896 3236 65900 3292
rect 65900 3236 65956 3292
rect 65956 3236 65960 3292
rect 65896 3232 65960 3236
rect 96376 3292 96440 3296
rect 96376 3236 96380 3292
rect 96380 3236 96436 3292
rect 96436 3236 96440 3292
rect 96376 3232 96440 3236
rect 96456 3292 96520 3296
rect 96456 3236 96460 3292
rect 96460 3236 96516 3292
rect 96516 3236 96520 3292
rect 96456 3232 96520 3236
rect 96536 3292 96600 3296
rect 96536 3236 96540 3292
rect 96540 3236 96596 3292
rect 96596 3236 96600 3292
rect 96536 3232 96600 3236
rect 96616 3292 96680 3296
rect 96616 3236 96620 3292
rect 96620 3236 96676 3292
rect 96676 3236 96680 3292
rect 96616 3232 96680 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 50296 2748 50360 2752
rect 50296 2692 50300 2748
rect 50300 2692 50356 2748
rect 50356 2692 50360 2748
rect 50296 2688 50360 2692
rect 50376 2748 50440 2752
rect 50376 2692 50380 2748
rect 50380 2692 50436 2748
rect 50436 2692 50440 2748
rect 50376 2688 50440 2692
rect 50456 2748 50520 2752
rect 50456 2692 50460 2748
rect 50460 2692 50516 2748
rect 50516 2692 50520 2748
rect 50456 2688 50520 2692
rect 50536 2748 50600 2752
rect 50536 2692 50540 2748
rect 50540 2692 50596 2748
rect 50596 2692 50600 2748
rect 50536 2688 50600 2692
rect 81016 2748 81080 2752
rect 81016 2692 81020 2748
rect 81020 2692 81076 2748
rect 81076 2692 81080 2748
rect 81016 2688 81080 2692
rect 81096 2748 81160 2752
rect 81096 2692 81100 2748
rect 81100 2692 81156 2748
rect 81156 2692 81160 2748
rect 81096 2688 81160 2692
rect 81176 2748 81240 2752
rect 81176 2692 81180 2748
rect 81180 2692 81236 2748
rect 81236 2692 81240 2748
rect 81176 2688 81240 2692
rect 81256 2748 81320 2752
rect 81256 2692 81260 2748
rect 81260 2692 81316 2748
rect 81316 2692 81320 2748
rect 81256 2688 81320 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
rect 65656 2204 65720 2208
rect 65656 2148 65660 2204
rect 65660 2148 65716 2204
rect 65716 2148 65720 2204
rect 65656 2144 65720 2148
rect 65736 2204 65800 2208
rect 65736 2148 65740 2204
rect 65740 2148 65796 2204
rect 65796 2148 65800 2204
rect 65736 2144 65800 2148
rect 65816 2204 65880 2208
rect 65816 2148 65820 2204
rect 65820 2148 65876 2204
rect 65876 2148 65880 2204
rect 65816 2144 65880 2148
rect 65896 2204 65960 2208
rect 65896 2148 65900 2204
rect 65900 2148 65956 2204
rect 65956 2148 65960 2204
rect 65896 2144 65960 2148
rect 96376 2204 96440 2208
rect 96376 2148 96380 2204
rect 96380 2148 96436 2204
rect 96436 2148 96440 2204
rect 96376 2144 96440 2148
rect 96456 2204 96520 2208
rect 96456 2148 96460 2204
rect 96460 2148 96516 2204
rect 96516 2148 96520 2204
rect 96456 2144 96520 2148
rect 96536 2204 96600 2208
rect 96536 2148 96540 2204
rect 96540 2148 96596 2204
rect 96596 2148 96600 2204
rect 96536 2144 96600 2148
rect 96616 2204 96680 2208
rect 96616 2148 96620 2204
rect 96620 2148 96676 2204
rect 96676 2148 96680 2204
rect 96616 2144 96680 2148
<< metal4 >>
rect 4208 37024 4528 37584
rect 19568 37568 19888 37584
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4868 2176 5188 37536
rect 5528 2176 5848 37536
rect 6188 2176 6508 37536
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 4208 2128 4528 2144
rect 19568 2128 19888 2688
rect 20228 2176 20548 37536
rect 20888 2176 21208 37536
rect 21548 2176 21868 37536
rect 34928 37024 35248 37584
rect 50288 37568 50608 37584
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 35588 2176 35908 37536
rect 36248 2176 36568 37536
rect 36908 2176 37228 37536
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 36480 50608 37504
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 35392 50608 36416
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 34304 50608 35328
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 33216 50608 34240
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 32128 50608 33152
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 31040 50608 32064
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 29952 50608 30976
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 28864 50608 29888
rect 50288 28800 50296 28864
rect 50360 28800 50376 28864
rect 50440 28800 50456 28864
rect 50520 28800 50536 28864
rect 50600 28800 50608 28864
rect 50288 27776 50608 28800
rect 50288 27712 50296 27776
rect 50360 27712 50376 27776
rect 50440 27712 50456 27776
rect 50520 27712 50536 27776
rect 50600 27712 50608 27776
rect 50288 26688 50608 27712
rect 50288 26624 50296 26688
rect 50360 26624 50376 26688
rect 50440 26624 50456 26688
rect 50520 26624 50536 26688
rect 50600 26624 50608 26688
rect 38515 26620 38581 26621
rect 38515 26556 38516 26620
rect 38580 26556 38581 26620
rect 38515 26555 38581 26556
rect 38518 21589 38578 26555
rect 50288 25600 50608 26624
rect 50288 25536 50296 25600
rect 50360 25536 50376 25600
rect 50440 25536 50456 25600
rect 50520 25536 50536 25600
rect 50600 25536 50608 25600
rect 50288 24512 50608 25536
rect 50288 24448 50296 24512
rect 50360 24448 50376 24512
rect 50440 24448 50456 24512
rect 50520 24448 50536 24512
rect 50600 24448 50608 24512
rect 50288 23424 50608 24448
rect 50288 23360 50296 23424
rect 50360 23360 50376 23424
rect 50440 23360 50456 23424
rect 50520 23360 50536 23424
rect 50600 23360 50608 23424
rect 50288 22336 50608 23360
rect 50288 22272 50296 22336
rect 50360 22272 50376 22336
rect 50440 22272 50456 22336
rect 50520 22272 50536 22336
rect 50600 22272 50608 22336
rect 38515 21588 38581 21589
rect 38515 21524 38516 21588
rect 38580 21524 38581 21588
rect 38515 21523 38581 21524
rect 50288 21248 50608 22272
rect 50288 21184 50296 21248
rect 50360 21184 50376 21248
rect 50440 21184 50456 21248
rect 50520 21184 50536 21248
rect 50600 21184 50608 21248
rect 50288 20160 50608 21184
rect 50288 20096 50296 20160
rect 50360 20096 50376 20160
rect 50440 20096 50456 20160
rect 50520 20096 50536 20160
rect 50600 20096 50608 20160
rect 50288 19072 50608 20096
rect 50288 19008 50296 19072
rect 50360 19008 50376 19072
rect 50440 19008 50456 19072
rect 50520 19008 50536 19072
rect 50600 19008 50608 19072
rect 38515 18868 38581 18869
rect 38515 18804 38516 18868
rect 38580 18804 38581 18868
rect 38515 18803 38581 18804
rect 38518 11389 38578 18803
rect 50288 17984 50608 19008
rect 50288 17920 50296 17984
rect 50360 17920 50376 17984
rect 50440 17920 50456 17984
rect 50520 17920 50536 17984
rect 50600 17920 50608 17984
rect 50288 16896 50608 17920
rect 50288 16832 50296 16896
rect 50360 16832 50376 16896
rect 50440 16832 50456 16896
rect 50520 16832 50536 16896
rect 50600 16832 50608 16896
rect 50288 15808 50608 16832
rect 50288 15744 50296 15808
rect 50360 15744 50376 15808
rect 50440 15744 50456 15808
rect 50520 15744 50536 15808
rect 50600 15744 50608 15808
rect 50288 14720 50608 15744
rect 50288 14656 50296 14720
rect 50360 14656 50376 14720
rect 50440 14656 50456 14720
rect 50520 14656 50536 14720
rect 50600 14656 50608 14720
rect 50288 13632 50608 14656
rect 50288 13568 50296 13632
rect 50360 13568 50376 13632
rect 50440 13568 50456 13632
rect 50520 13568 50536 13632
rect 50600 13568 50608 13632
rect 50288 12544 50608 13568
rect 50288 12480 50296 12544
rect 50360 12480 50376 12544
rect 50440 12480 50456 12544
rect 50520 12480 50536 12544
rect 50600 12480 50608 12544
rect 38699 12340 38765 12341
rect 38699 12276 38700 12340
rect 38764 12276 38765 12340
rect 38699 12275 38765 12276
rect 38515 11388 38581 11389
rect 38515 11324 38516 11388
rect 38580 11324 38581 11388
rect 38515 11323 38581 11324
rect 38702 11117 38762 12275
rect 50288 11456 50608 12480
rect 50288 11392 50296 11456
rect 50360 11392 50376 11456
rect 50440 11392 50456 11456
rect 50520 11392 50536 11456
rect 50600 11392 50608 11456
rect 38699 11116 38765 11117
rect 38699 11052 38700 11116
rect 38764 11052 38765 11116
rect 38699 11051 38765 11052
rect 50288 10368 50608 11392
rect 50288 10304 50296 10368
rect 50360 10304 50376 10368
rect 50440 10304 50456 10368
rect 50520 10304 50536 10368
rect 50600 10304 50608 10368
rect 50288 9280 50608 10304
rect 50288 9216 50296 9280
rect 50360 9216 50376 9280
rect 50440 9216 50456 9280
rect 50520 9216 50536 9280
rect 50600 9216 50608 9280
rect 50288 8192 50608 9216
rect 50288 8128 50296 8192
rect 50360 8128 50376 8192
rect 50440 8128 50456 8192
rect 50520 8128 50536 8192
rect 50600 8128 50608 8192
rect 50288 7104 50608 8128
rect 50288 7040 50296 7104
rect 50360 7040 50376 7104
rect 50440 7040 50456 7104
rect 50520 7040 50536 7104
rect 50600 7040 50608 7104
rect 50288 6016 50608 7040
rect 50288 5952 50296 6016
rect 50360 5952 50376 6016
rect 50440 5952 50456 6016
rect 50520 5952 50536 6016
rect 50600 5952 50608 6016
rect 50288 4928 50608 5952
rect 50288 4864 50296 4928
rect 50360 4864 50376 4928
rect 50440 4864 50456 4928
rect 50520 4864 50536 4928
rect 50600 4864 50608 4928
rect 50288 3840 50608 4864
rect 50288 3776 50296 3840
rect 50360 3776 50376 3840
rect 50440 3776 50456 3840
rect 50520 3776 50536 3840
rect 50600 3776 50608 3840
rect 50288 2752 50608 3776
rect 50288 2688 50296 2752
rect 50360 2688 50376 2752
rect 50440 2688 50456 2752
rect 50520 2688 50536 2752
rect 50600 2688 50608 2752
rect 34928 2128 35248 2144
rect 50288 2128 50608 2688
rect 50948 2176 51268 37536
rect 51608 2176 51928 37536
rect 52268 2176 52588 37536
rect 65648 37024 65968 37584
rect 81008 37568 81328 37584
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 35936 65968 36960
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 34848 65968 35872
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 33760 65968 34784
rect 65648 33696 65656 33760
rect 65720 33696 65736 33760
rect 65800 33696 65816 33760
rect 65880 33696 65896 33760
rect 65960 33696 65968 33760
rect 65648 32672 65968 33696
rect 65648 32608 65656 32672
rect 65720 32608 65736 32672
rect 65800 32608 65816 32672
rect 65880 32608 65896 32672
rect 65960 32608 65968 32672
rect 65648 31584 65968 32608
rect 65648 31520 65656 31584
rect 65720 31520 65736 31584
rect 65800 31520 65816 31584
rect 65880 31520 65896 31584
rect 65960 31520 65968 31584
rect 65648 30496 65968 31520
rect 65648 30432 65656 30496
rect 65720 30432 65736 30496
rect 65800 30432 65816 30496
rect 65880 30432 65896 30496
rect 65960 30432 65968 30496
rect 65648 29408 65968 30432
rect 65648 29344 65656 29408
rect 65720 29344 65736 29408
rect 65800 29344 65816 29408
rect 65880 29344 65896 29408
rect 65960 29344 65968 29408
rect 65648 28320 65968 29344
rect 65648 28256 65656 28320
rect 65720 28256 65736 28320
rect 65800 28256 65816 28320
rect 65880 28256 65896 28320
rect 65960 28256 65968 28320
rect 65648 27232 65968 28256
rect 65648 27168 65656 27232
rect 65720 27168 65736 27232
rect 65800 27168 65816 27232
rect 65880 27168 65896 27232
rect 65960 27168 65968 27232
rect 65648 26144 65968 27168
rect 65648 26080 65656 26144
rect 65720 26080 65736 26144
rect 65800 26080 65816 26144
rect 65880 26080 65896 26144
rect 65960 26080 65968 26144
rect 65648 25056 65968 26080
rect 65648 24992 65656 25056
rect 65720 24992 65736 25056
rect 65800 24992 65816 25056
rect 65880 24992 65896 25056
rect 65960 24992 65968 25056
rect 65648 23968 65968 24992
rect 65648 23904 65656 23968
rect 65720 23904 65736 23968
rect 65800 23904 65816 23968
rect 65880 23904 65896 23968
rect 65960 23904 65968 23968
rect 65648 22880 65968 23904
rect 65648 22816 65656 22880
rect 65720 22816 65736 22880
rect 65800 22816 65816 22880
rect 65880 22816 65896 22880
rect 65960 22816 65968 22880
rect 65648 21792 65968 22816
rect 65648 21728 65656 21792
rect 65720 21728 65736 21792
rect 65800 21728 65816 21792
rect 65880 21728 65896 21792
rect 65960 21728 65968 21792
rect 65648 20704 65968 21728
rect 65648 20640 65656 20704
rect 65720 20640 65736 20704
rect 65800 20640 65816 20704
rect 65880 20640 65896 20704
rect 65960 20640 65968 20704
rect 65648 19616 65968 20640
rect 65648 19552 65656 19616
rect 65720 19552 65736 19616
rect 65800 19552 65816 19616
rect 65880 19552 65896 19616
rect 65960 19552 65968 19616
rect 65648 18528 65968 19552
rect 65648 18464 65656 18528
rect 65720 18464 65736 18528
rect 65800 18464 65816 18528
rect 65880 18464 65896 18528
rect 65960 18464 65968 18528
rect 65648 17440 65968 18464
rect 65648 17376 65656 17440
rect 65720 17376 65736 17440
rect 65800 17376 65816 17440
rect 65880 17376 65896 17440
rect 65960 17376 65968 17440
rect 65648 16352 65968 17376
rect 65648 16288 65656 16352
rect 65720 16288 65736 16352
rect 65800 16288 65816 16352
rect 65880 16288 65896 16352
rect 65960 16288 65968 16352
rect 65648 15264 65968 16288
rect 65648 15200 65656 15264
rect 65720 15200 65736 15264
rect 65800 15200 65816 15264
rect 65880 15200 65896 15264
rect 65960 15200 65968 15264
rect 65648 14176 65968 15200
rect 65648 14112 65656 14176
rect 65720 14112 65736 14176
rect 65800 14112 65816 14176
rect 65880 14112 65896 14176
rect 65960 14112 65968 14176
rect 65648 13088 65968 14112
rect 65648 13024 65656 13088
rect 65720 13024 65736 13088
rect 65800 13024 65816 13088
rect 65880 13024 65896 13088
rect 65960 13024 65968 13088
rect 65648 12000 65968 13024
rect 65648 11936 65656 12000
rect 65720 11936 65736 12000
rect 65800 11936 65816 12000
rect 65880 11936 65896 12000
rect 65960 11936 65968 12000
rect 65648 10912 65968 11936
rect 65648 10848 65656 10912
rect 65720 10848 65736 10912
rect 65800 10848 65816 10912
rect 65880 10848 65896 10912
rect 65960 10848 65968 10912
rect 65648 9824 65968 10848
rect 65648 9760 65656 9824
rect 65720 9760 65736 9824
rect 65800 9760 65816 9824
rect 65880 9760 65896 9824
rect 65960 9760 65968 9824
rect 65648 8736 65968 9760
rect 65648 8672 65656 8736
rect 65720 8672 65736 8736
rect 65800 8672 65816 8736
rect 65880 8672 65896 8736
rect 65960 8672 65968 8736
rect 65648 7648 65968 8672
rect 65648 7584 65656 7648
rect 65720 7584 65736 7648
rect 65800 7584 65816 7648
rect 65880 7584 65896 7648
rect 65960 7584 65968 7648
rect 65648 6560 65968 7584
rect 65648 6496 65656 6560
rect 65720 6496 65736 6560
rect 65800 6496 65816 6560
rect 65880 6496 65896 6560
rect 65960 6496 65968 6560
rect 65648 5472 65968 6496
rect 65648 5408 65656 5472
rect 65720 5408 65736 5472
rect 65800 5408 65816 5472
rect 65880 5408 65896 5472
rect 65960 5408 65968 5472
rect 65648 4384 65968 5408
rect 65648 4320 65656 4384
rect 65720 4320 65736 4384
rect 65800 4320 65816 4384
rect 65880 4320 65896 4384
rect 65960 4320 65968 4384
rect 65648 3296 65968 4320
rect 65648 3232 65656 3296
rect 65720 3232 65736 3296
rect 65800 3232 65816 3296
rect 65880 3232 65896 3296
rect 65960 3232 65968 3296
rect 65648 2208 65968 3232
rect 65648 2144 65656 2208
rect 65720 2144 65736 2208
rect 65800 2144 65816 2208
rect 65880 2144 65896 2208
rect 65960 2144 65968 2208
rect 66308 2176 66628 37536
rect 66968 2176 67288 37536
rect 67628 2176 67948 37536
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 36480 81328 37504
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 35392 81328 36416
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 34304 81328 35328
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 33216 81328 34240
rect 81008 33152 81016 33216
rect 81080 33152 81096 33216
rect 81160 33152 81176 33216
rect 81240 33152 81256 33216
rect 81320 33152 81328 33216
rect 81008 32128 81328 33152
rect 81008 32064 81016 32128
rect 81080 32064 81096 32128
rect 81160 32064 81176 32128
rect 81240 32064 81256 32128
rect 81320 32064 81328 32128
rect 81008 31040 81328 32064
rect 81008 30976 81016 31040
rect 81080 30976 81096 31040
rect 81160 30976 81176 31040
rect 81240 30976 81256 31040
rect 81320 30976 81328 31040
rect 81008 29952 81328 30976
rect 81008 29888 81016 29952
rect 81080 29888 81096 29952
rect 81160 29888 81176 29952
rect 81240 29888 81256 29952
rect 81320 29888 81328 29952
rect 81008 28864 81328 29888
rect 81008 28800 81016 28864
rect 81080 28800 81096 28864
rect 81160 28800 81176 28864
rect 81240 28800 81256 28864
rect 81320 28800 81328 28864
rect 81008 27776 81328 28800
rect 81008 27712 81016 27776
rect 81080 27712 81096 27776
rect 81160 27712 81176 27776
rect 81240 27712 81256 27776
rect 81320 27712 81328 27776
rect 81008 26688 81328 27712
rect 81008 26624 81016 26688
rect 81080 26624 81096 26688
rect 81160 26624 81176 26688
rect 81240 26624 81256 26688
rect 81320 26624 81328 26688
rect 81008 25600 81328 26624
rect 81008 25536 81016 25600
rect 81080 25536 81096 25600
rect 81160 25536 81176 25600
rect 81240 25536 81256 25600
rect 81320 25536 81328 25600
rect 81008 24512 81328 25536
rect 81008 24448 81016 24512
rect 81080 24448 81096 24512
rect 81160 24448 81176 24512
rect 81240 24448 81256 24512
rect 81320 24448 81328 24512
rect 81008 23424 81328 24448
rect 81008 23360 81016 23424
rect 81080 23360 81096 23424
rect 81160 23360 81176 23424
rect 81240 23360 81256 23424
rect 81320 23360 81328 23424
rect 81008 22336 81328 23360
rect 81008 22272 81016 22336
rect 81080 22272 81096 22336
rect 81160 22272 81176 22336
rect 81240 22272 81256 22336
rect 81320 22272 81328 22336
rect 81008 21248 81328 22272
rect 81008 21184 81016 21248
rect 81080 21184 81096 21248
rect 81160 21184 81176 21248
rect 81240 21184 81256 21248
rect 81320 21184 81328 21248
rect 81008 20160 81328 21184
rect 81008 20096 81016 20160
rect 81080 20096 81096 20160
rect 81160 20096 81176 20160
rect 81240 20096 81256 20160
rect 81320 20096 81328 20160
rect 81008 19072 81328 20096
rect 81008 19008 81016 19072
rect 81080 19008 81096 19072
rect 81160 19008 81176 19072
rect 81240 19008 81256 19072
rect 81320 19008 81328 19072
rect 81008 17984 81328 19008
rect 81008 17920 81016 17984
rect 81080 17920 81096 17984
rect 81160 17920 81176 17984
rect 81240 17920 81256 17984
rect 81320 17920 81328 17984
rect 81008 16896 81328 17920
rect 81008 16832 81016 16896
rect 81080 16832 81096 16896
rect 81160 16832 81176 16896
rect 81240 16832 81256 16896
rect 81320 16832 81328 16896
rect 81008 15808 81328 16832
rect 81008 15744 81016 15808
rect 81080 15744 81096 15808
rect 81160 15744 81176 15808
rect 81240 15744 81256 15808
rect 81320 15744 81328 15808
rect 81008 14720 81328 15744
rect 81008 14656 81016 14720
rect 81080 14656 81096 14720
rect 81160 14656 81176 14720
rect 81240 14656 81256 14720
rect 81320 14656 81328 14720
rect 81008 13632 81328 14656
rect 81008 13568 81016 13632
rect 81080 13568 81096 13632
rect 81160 13568 81176 13632
rect 81240 13568 81256 13632
rect 81320 13568 81328 13632
rect 81008 12544 81328 13568
rect 81008 12480 81016 12544
rect 81080 12480 81096 12544
rect 81160 12480 81176 12544
rect 81240 12480 81256 12544
rect 81320 12480 81328 12544
rect 81008 11456 81328 12480
rect 81008 11392 81016 11456
rect 81080 11392 81096 11456
rect 81160 11392 81176 11456
rect 81240 11392 81256 11456
rect 81320 11392 81328 11456
rect 81008 10368 81328 11392
rect 81008 10304 81016 10368
rect 81080 10304 81096 10368
rect 81160 10304 81176 10368
rect 81240 10304 81256 10368
rect 81320 10304 81328 10368
rect 81008 9280 81328 10304
rect 81008 9216 81016 9280
rect 81080 9216 81096 9280
rect 81160 9216 81176 9280
rect 81240 9216 81256 9280
rect 81320 9216 81328 9280
rect 81008 8192 81328 9216
rect 81008 8128 81016 8192
rect 81080 8128 81096 8192
rect 81160 8128 81176 8192
rect 81240 8128 81256 8192
rect 81320 8128 81328 8192
rect 81008 7104 81328 8128
rect 81008 7040 81016 7104
rect 81080 7040 81096 7104
rect 81160 7040 81176 7104
rect 81240 7040 81256 7104
rect 81320 7040 81328 7104
rect 81008 6016 81328 7040
rect 81008 5952 81016 6016
rect 81080 5952 81096 6016
rect 81160 5952 81176 6016
rect 81240 5952 81256 6016
rect 81320 5952 81328 6016
rect 81008 4928 81328 5952
rect 81008 4864 81016 4928
rect 81080 4864 81096 4928
rect 81160 4864 81176 4928
rect 81240 4864 81256 4928
rect 81320 4864 81328 4928
rect 81008 3840 81328 4864
rect 81008 3776 81016 3840
rect 81080 3776 81096 3840
rect 81160 3776 81176 3840
rect 81240 3776 81256 3840
rect 81320 3776 81328 3840
rect 81008 2752 81328 3776
rect 81008 2688 81016 2752
rect 81080 2688 81096 2752
rect 81160 2688 81176 2752
rect 81240 2688 81256 2752
rect 81320 2688 81328 2752
rect 65648 2128 65968 2144
rect 81008 2128 81328 2688
rect 81668 2176 81988 37536
rect 82328 2176 82648 37536
rect 82988 2176 83308 37536
rect 96368 37024 96688 37584
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 35936 96688 36960
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 34848 96688 35872
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 33760 96688 34784
rect 96368 33696 96376 33760
rect 96440 33696 96456 33760
rect 96520 33696 96536 33760
rect 96600 33696 96616 33760
rect 96680 33696 96688 33760
rect 96368 32672 96688 33696
rect 96368 32608 96376 32672
rect 96440 32608 96456 32672
rect 96520 32608 96536 32672
rect 96600 32608 96616 32672
rect 96680 32608 96688 32672
rect 96368 31584 96688 32608
rect 96368 31520 96376 31584
rect 96440 31520 96456 31584
rect 96520 31520 96536 31584
rect 96600 31520 96616 31584
rect 96680 31520 96688 31584
rect 96368 30496 96688 31520
rect 96368 30432 96376 30496
rect 96440 30432 96456 30496
rect 96520 30432 96536 30496
rect 96600 30432 96616 30496
rect 96680 30432 96688 30496
rect 96368 29408 96688 30432
rect 96368 29344 96376 29408
rect 96440 29344 96456 29408
rect 96520 29344 96536 29408
rect 96600 29344 96616 29408
rect 96680 29344 96688 29408
rect 96368 28320 96688 29344
rect 96368 28256 96376 28320
rect 96440 28256 96456 28320
rect 96520 28256 96536 28320
rect 96600 28256 96616 28320
rect 96680 28256 96688 28320
rect 96368 27232 96688 28256
rect 96368 27168 96376 27232
rect 96440 27168 96456 27232
rect 96520 27168 96536 27232
rect 96600 27168 96616 27232
rect 96680 27168 96688 27232
rect 96368 26144 96688 27168
rect 96368 26080 96376 26144
rect 96440 26080 96456 26144
rect 96520 26080 96536 26144
rect 96600 26080 96616 26144
rect 96680 26080 96688 26144
rect 96368 25056 96688 26080
rect 96368 24992 96376 25056
rect 96440 24992 96456 25056
rect 96520 24992 96536 25056
rect 96600 24992 96616 25056
rect 96680 24992 96688 25056
rect 96368 23968 96688 24992
rect 96368 23904 96376 23968
rect 96440 23904 96456 23968
rect 96520 23904 96536 23968
rect 96600 23904 96616 23968
rect 96680 23904 96688 23968
rect 96368 22880 96688 23904
rect 96368 22816 96376 22880
rect 96440 22816 96456 22880
rect 96520 22816 96536 22880
rect 96600 22816 96616 22880
rect 96680 22816 96688 22880
rect 96368 21792 96688 22816
rect 96368 21728 96376 21792
rect 96440 21728 96456 21792
rect 96520 21728 96536 21792
rect 96600 21728 96616 21792
rect 96680 21728 96688 21792
rect 96368 20704 96688 21728
rect 96368 20640 96376 20704
rect 96440 20640 96456 20704
rect 96520 20640 96536 20704
rect 96600 20640 96616 20704
rect 96680 20640 96688 20704
rect 96368 19616 96688 20640
rect 96368 19552 96376 19616
rect 96440 19552 96456 19616
rect 96520 19552 96536 19616
rect 96600 19552 96616 19616
rect 96680 19552 96688 19616
rect 96368 18528 96688 19552
rect 96368 18464 96376 18528
rect 96440 18464 96456 18528
rect 96520 18464 96536 18528
rect 96600 18464 96616 18528
rect 96680 18464 96688 18528
rect 96368 17440 96688 18464
rect 96368 17376 96376 17440
rect 96440 17376 96456 17440
rect 96520 17376 96536 17440
rect 96600 17376 96616 17440
rect 96680 17376 96688 17440
rect 96368 16352 96688 17376
rect 96368 16288 96376 16352
rect 96440 16288 96456 16352
rect 96520 16288 96536 16352
rect 96600 16288 96616 16352
rect 96680 16288 96688 16352
rect 96368 15264 96688 16288
rect 96368 15200 96376 15264
rect 96440 15200 96456 15264
rect 96520 15200 96536 15264
rect 96600 15200 96616 15264
rect 96680 15200 96688 15264
rect 96368 14176 96688 15200
rect 96368 14112 96376 14176
rect 96440 14112 96456 14176
rect 96520 14112 96536 14176
rect 96600 14112 96616 14176
rect 96680 14112 96688 14176
rect 96368 13088 96688 14112
rect 96368 13024 96376 13088
rect 96440 13024 96456 13088
rect 96520 13024 96536 13088
rect 96600 13024 96616 13088
rect 96680 13024 96688 13088
rect 96368 12000 96688 13024
rect 96368 11936 96376 12000
rect 96440 11936 96456 12000
rect 96520 11936 96536 12000
rect 96600 11936 96616 12000
rect 96680 11936 96688 12000
rect 96368 10912 96688 11936
rect 96368 10848 96376 10912
rect 96440 10848 96456 10912
rect 96520 10848 96536 10912
rect 96600 10848 96616 10912
rect 96680 10848 96688 10912
rect 96368 9824 96688 10848
rect 96368 9760 96376 9824
rect 96440 9760 96456 9824
rect 96520 9760 96536 9824
rect 96600 9760 96616 9824
rect 96680 9760 96688 9824
rect 96368 8736 96688 9760
rect 96368 8672 96376 8736
rect 96440 8672 96456 8736
rect 96520 8672 96536 8736
rect 96600 8672 96616 8736
rect 96680 8672 96688 8736
rect 96368 7648 96688 8672
rect 96368 7584 96376 7648
rect 96440 7584 96456 7648
rect 96520 7584 96536 7648
rect 96600 7584 96616 7648
rect 96680 7584 96688 7648
rect 96368 6560 96688 7584
rect 96368 6496 96376 6560
rect 96440 6496 96456 6560
rect 96520 6496 96536 6560
rect 96600 6496 96616 6560
rect 96680 6496 96688 6560
rect 96368 5472 96688 6496
rect 96368 5408 96376 5472
rect 96440 5408 96456 5472
rect 96520 5408 96536 5472
rect 96600 5408 96616 5472
rect 96680 5408 96688 5472
rect 96368 4384 96688 5408
rect 96368 4320 96376 4384
rect 96440 4320 96456 4384
rect 96520 4320 96536 4384
rect 96600 4320 96616 4384
rect 96680 4320 96688 4384
rect 96368 3296 96688 4320
rect 96368 3232 96376 3296
rect 96440 3232 96456 3296
rect 96520 3232 96536 3296
rect 96600 3232 96616 3296
rect 96680 3232 96688 3296
rect 96368 2208 96688 3232
rect 96368 2144 96376 2208
rect 96440 2144 96456 2208
rect 96520 2144 96536 2208
rect 96600 2144 96616 2208
rect 96680 2144 96688 2208
rect 97028 2176 97348 37536
rect 97688 2176 98008 37536
rect 96368 2128 96688 2144
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1623939100
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  input296 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 1748 0 -1 2720
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  input330 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 1472 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input341
timestamp 1623939100
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 2760 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1623939100
transform 1 0 2300 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input319 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 3864 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input322
timestamp 1623939100
transform 1 0 4232 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input323
timestamp 1623939100
transform 1 0 4784 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26
timestamp 1623939100
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1623939100
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1623939100
transform 1 0 3496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36
timestamp 1623939100
transform 1 0 4416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1623939100
transform 1 0 5336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43
timestamp 1623939100
transform 1 0 5060 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input324
timestamp 1623939100
transform 1 0 5428 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_53
timestamp 1623939100
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53
timestamp 1623939100
transform 1 0 5980 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input298 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_58
timestamp 1623939100
transform 1 0 6440 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1623939100
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1623939100
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input326
timestamp 1623939100
transform 1 0 6808 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1623939100
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1623939100
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input325
timestamp 1623939100
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input331
timestamp 1623939100
transform 1 0 8188 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input358 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 7728 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69
timestamp 1623939100
transform 1 0 7452 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1623939100
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1623939100
transform 1 0 7360 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_78
timestamp 1623939100
transform 1 0 8280 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1623939100
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input332
timestamp 1623939100
transform 1 0 9016 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input333
timestamp 1623939100
transform 1 0 9568 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input334
timestamp 1623939100
transform 1 0 10212 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1623939100
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101
timestamp 1623939100
transform 1 0 10396 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_92 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 9568 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_98
timestamp 1623939100
transform 1 0 10120 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_108
timestamp 1623939100
transform 1 0 11040 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_110
timestamp 1623939100
transform 1 0 11224 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105
timestamp 1623939100
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input335 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 10856 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1623939100
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1623939100
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1623939100
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1623939100
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input337
timestamp 1623939100
transform 1 0 12052 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input336
timestamp 1623939100
transform 1 0 12236 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_125
timestamp 1623939100
transform 1 0 12604 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1623939100
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input338
timestamp 1623939100
transform 1 0 13156 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input339
timestamp 1623939100
transform 1 0 13248 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input340
timestamp 1623939100
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127
timestamp 1623939100
transform 1 0 12788 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137
timestamp 1623939100
transform 1 0 13708 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_131
timestamp 1623939100
transform 1 0 13156 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1623939100
transform 1 0 13800 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_154
timestamp 1623939100
transform 1 0 15272 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_146
timestamp 1623939100
transform 1 0 14536 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1623939100
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output585 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 14904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input342
timestamp 1623939100
transform 1 0 14904 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_163
timestamp 1623939100
transform 1 0 16100 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_158
timestamp 1623939100
transform 1 0 15640 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1623939100
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input344
timestamp 1623939100
transform 1 0 15732 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input343
timestamp 1623939100
transform 1 0 15824 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_166
timestamp 1623939100
transform 1 0 16376 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1623939100
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1623939100
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input345
timestamp 1623939100
transform 1 0 17572 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input346
timestamp 1623939100
transform 1 0 17296 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input348
timestamp 1623939100
transform 1 0 18216 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1623939100
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_185
timestamp 1623939100
transform 1 0 18124 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1623939100
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_182
timestamp 1623939100
transform 1 0 17848 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1623939100
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input347
timestamp 1623939100
transform 1 0 18492 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input349
timestamp 1623939100
transform 1 0 19136 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input350
timestamp 1623939100
transform 1 0 20056 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input351
timestamp 1623939100
transform 1 0 20240 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_195
timestamp 1623939100
transform 1 0 19044 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1623939100
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1623939100
transform 1 0 18768 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1623939100
transform 1 0 19688 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1623939100
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input353
timestamp 1623939100
transform 1 0 20792 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input354
timestamp 1623939100
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_214
timestamp 1623939100
transform 1 0 20792 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_224
timestamp 1623939100
transform 1 0 21712 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_210
timestamp 1623939100
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_218
timestamp 1623939100
transform 1 0 21160 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_226 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1623939100
transform 1 0 22172 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_233
timestamp 1623939100
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output600
timestamp 1623939100
transform 1 0 22540 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1623939100
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1623939100
transform 1 0 22908 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_253 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform -1 0 22908 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output447
timestamp 1623939100
transform -1 0 23276 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1623939100
transform 1 0 23276 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input78
timestamp 1623939100
transform 1 0 23276 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1623939100
transform 1 0 23552 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output486
timestamp 1623939100
transform 1 0 23644 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 1623939100
transform 1 0 23920 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_249
timestamp 1623939100
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_251
timestamp 1623939100
transform 1 0 24196 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output497
timestamp 1623939100
transform 1 0 24380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_261
timestamp 1623939100
transform 1 0 25116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_257
timestamp 1623939100
transform 1 0 24748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1623939100
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1623939100
transform 1 0 24748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1623939100
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 24840 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1623939100
transform 1 0 25852 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_270
timestamp 1623939100
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_316
timestamp 1623939100
transform -1 0 25576 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output541
timestamp 1623939100
transform 1 0 25484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output508
timestamp 1623939100
transform -1 0 25944 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_277
timestamp 1623939100
transform 1 0 26588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1623939100
transform 1 0 26680 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_322
timestamp 1623939100
transform -1 0 26312 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output552
timestamp 1623939100
transform 1 0 26220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output519
timestamp 1623939100
transform -1 0 26680 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_286
timestamp 1623939100
transform 1 0 27416 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1623939100
transform 1 0 27416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_376
timestamp 1623939100
transform -1 0 27784 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_332
timestamp 1623939100
transform -1 0 27048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output530
timestamp 1623939100
transform -1 0 27416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1623939100
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_291
timestamp 1623939100
transform 1 0 27876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output574
timestamp 1623939100
transform -1 0 28152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1623939100
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_294
timestamp 1623939100
transform 1 0 28152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_273
timestamp 1623939100
transform -1 0 28244 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_235
timestamp 1623939100
transform 1 0 28336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output458
timestamp 1623939100
transform -1 0 28612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_301
timestamp 1623939100
transform 1 0 28796 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1623939100
transform 1 0 28612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _561_
timestamp 1623939100
transform 1 0 28520 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output469
timestamp 1623939100
transform 1 0 28980 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1623939100
transform 1 0 29164 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_308
timestamp 1623939100
transform 1 0 29440 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_307
timestamp 1623939100
transform 1 0 29348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output478
timestamp 1623939100
transform 1 0 29716 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1623939100
transform 1 0 29808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_315
timestamp 1623939100
transform 1 0 30084 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1623939100
transform 1 0 30084 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_322
timestamp 1623939100
transform 1 0 30728 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1623939100
transform 1 0 30544 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1623939100
transform 1 0 30452 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1623939100
transform 1 0 30452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output479
timestamp 1623939100
transform 1 0 30912 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1623939100
transform 1 0 31096 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_329
timestamp 1623939100
transform 1 0 31372 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_328
timestamp 1623939100
transform 1 0 31280 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output480
timestamp 1623939100
transform 1 0 31648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 1623939100
transform 1 0 31740 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_336
timestamp 1623939100
transform 1 0 32016 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_336
timestamp 1623939100
transform 1 0 32016 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output481
timestamp 1623939100
transform 1 0 32384 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_343
timestamp 1623939100
transform 1 0 32660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_344
timestamp 1623939100
transform 1 0 32752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1623939100
transform 1 0 33028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1623939100
transform 1 0 32568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_350
timestamp 1623939100
transform 1 0 33304 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1623939100
transform 1 0 33212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output482
timestamp 1623939100
transform 1 0 33580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1623939100
transform 1 0 33120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input77
timestamp 1623939100
transform 1 0 33672 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _281_
timestamp 1623939100
transform 1 0 35328 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 1623939100
transform 1 0 34316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output483
timestamp 1623939100
transform 1 0 34316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output484
timestamp 1623939100
transform 1 0 35052 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_357
timestamp 1623939100
transform 1 0 33948 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1623939100
transform 1 0 34684 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1623939100
transform 1 0 35420 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_357
timestamp 1623939100
transform 1 0 33948 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_364
timestamp 1623939100
transform 1 0 34592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_378
timestamp 1623939100
transform 1 0 35880 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_378
timestamp 1623939100
transform 1 0 35880 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_294
timestamp 1623939100
transform -1 0 36248 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1623939100
transform 1 0 35788 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_386
timestamp 1623939100
transform 1 0 36616 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_297
timestamp 1623939100
transform -1 0 36984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_295
timestamp 1623939100
transform -1 0 36800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output490
timestamp 1623939100
transform 1 0 36248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output485
timestamp 1623939100
transform -1 0 36616 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1623939100
transform 1 0 37260 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_394
timestamp 1623939100
transform 1 0 37352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output487
timestamp 1623939100
transform -1 0 37352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1623939100
transform 1 0 36984 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_400
timestamp 1623939100
transform 1 0 37904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_402
timestamp 1623939100
transform 1 0 38088 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_306
timestamp 1623939100
transform -1 0 38272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output493
timestamp 1623939100
transform -1 0 38640 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output488
timestamp 1623939100
transform 1 0 37720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1623939100
transform 1 0 37812 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_408
timestamp 1623939100
transform 1 0 38640 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_407
timestamp 1623939100
transform 1 0 38548 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_299
timestamp 1623939100
transform -1 0 38916 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output489
timestamp 1623939100
transform -1 0 39284 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1623939100
transform 1 0 39008 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1623939100
transform 1 0 38456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_415
timestamp 1623939100
transform 1 0 39284 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_415
timestamp 1623939100
transform 1 0 39284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_423
timestamp 1623939100
transform 1 0 40020 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_423
timestamp 1623939100
transform 1 0 40020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_303
timestamp 1623939100
transform -1 0 40388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_301
timestamp 1623939100
transform -1 0 39652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output498
timestamp 1623939100
transform 1 0 40112 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output491
timestamp 1623939100
transform -1 0 40020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_428
timestamp 1623939100
transform 1 0 40480 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_433
timestamp 1623939100
transform 1 0 40940 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_304
timestamp 1623939100
transform -1 0 40940 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output492
timestamp 1623939100
transform -1 0 40756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_436
timestamp 1623939100
transform 1 0 41216 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_436
timestamp 1623939100
transform 1 0 41216 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output500
timestamp 1623939100
transform 1 0 41308 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1623939100
transform 1 0 41124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_441
timestamp 1623939100
transform 1 0 41676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1623939100
transform 1 0 41952 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output494
timestamp 1623939100
transform 1 0 41584 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 1623939100
transform 1 0 42044 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_448
timestamp 1623939100
transform 1 0 42320 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1623939100
transform 1 0 42688 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output495
timestamp 1623939100
transform 1 0 42320 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_457
timestamp 1623939100
transform 1 0 43148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output496
timestamp 1623939100
transform 1 0 43056 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1623939100
transform 1 0 43056 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_460
timestamp 1623939100
transform 1 0 43424 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output503
timestamp 1623939100
transform 1 0 43516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_465
timestamp 1623939100
transform 1 0 43884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_465
timestamp 1623939100
transform 1 0 43884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_308
timestamp 1623939100
transform -1 0 44252 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1623939100
transform 1 0 43792 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_472
timestamp 1623939100
transform 1 0 44528 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output499
timestamp 1623939100
transform -1 0 44620 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 1623939100
transform 1 0 44252 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_473
timestamp 1623939100
transform 1 0 44620 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_309
timestamp 1623939100
transform -1 0 44988 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output501
timestamp 1623939100
transform -1 0 45356 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 1623939100
transform 1 0 44896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_479
timestamp 1623939100
transform 1 0 45172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_481
timestamp 1623939100
transform 1 0 45356 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_314
timestamp 1623939100
transform -1 0 45540 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output507
timestamp 1623939100
transform -1 0 45908 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1623939100
transform 1 0 45908 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output502
timestamp 1623939100
transform 1 0 45724 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1623939100
transform 1 0 46092 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output509
timestamp 1623939100
transform 1 0 46276 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1623939100
transform 1 0 46460 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_495
timestamp 1623939100
transform 1 0 46644 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_494
timestamp 1623939100
transform 1 0 46552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_318
timestamp 1623939100
transform -1 0 47012 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output504
timestamp 1623939100
transform 1 0 46920 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output510
timestamp 1623939100
transform -1 0 47380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_503
timestamp 1623939100
transform 1 0 47380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_502
timestamp 1623939100
transform 1 0 47288 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output505
timestamp 1623939100
transform 1 0 47656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_514
timestamp 1623939100
transform 1 0 48392 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_511
timestamp 1623939100
transform 1 0 48116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_510
timestamp 1623939100
transform 1 0 48024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_311
timestamp 1623939100
transform -1 0 48392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output506
timestamp 1623939100
transform -1 0 48760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1623939100
transform 1 0 48300 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_520
timestamp 1623939100
transform 1 0 48944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_312
timestamp 1623939100
transform -1 0 48944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output512
timestamp 1623939100
transform 1 0 48760 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_522
timestamp 1623939100
transform 1 0 49128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_523
timestamp 1623939100
transform 1 0 49220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_320
timestamp 1623939100
transform -1 0 49496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output514
timestamp 1623939100
transform -1 0 49864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1623939100
transform 1 0 49128 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_530
timestamp 1623939100
transform 1 0 49864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_529
timestamp 1623939100
transform 1 0 49772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input106
timestamp 1623939100
transform 1 0 50232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _385_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 49864 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_537
timestamp 1623939100
transform 1 0 50508 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1623939100
transform 1 0 50416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output511
timestamp 1623939100
transform 1 0 50784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_547
timestamp 1623939100
transform 1 0 51428 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_550
timestamp 1623939100
transform 1 0 51704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_544
timestamp 1623939100
transform 1 0 51152 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output517
timestamp 1623939100
transform 1 0 51060 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_554
timestamp 1623939100
transform 1 0 52072 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_552
timestamp 1623939100
transform 1 0 51888 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output513
timestamp 1623939100
transform 1 0 52256 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 1623939100
transform 1 0 52440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 1623939100
transform 1 0 51796 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1623939100
transform 1 0 51796 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_561
timestamp 1623939100
transform 1 0 52716 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_560
timestamp 1623939100
transform 1 0 52624 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1623939100
transform 1 0 53636 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_569
timestamp 1623939100
transform 1 0 53452 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_568
timestamp 1623939100
transform 1 0 53360 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output515
timestamp 1623939100
transform 1 0 52992 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1623939100
transform 1 0 53544 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_579
timestamp 1623939100
transform 1 0 54372 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_576
timestamp 1623939100
transform 1 0 54096 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output522
timestamp 1623939100
transform 1 0 54004 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output516
timestamp 1623939100
transform 1 0 53728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1623939100
transform 1 0 54464 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_581
timestamp 1623939100
transform 1 0 54556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_589
timestamp 1623939100
transform 1 0 55292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_327
timestamp 1623939100
transform -1 0 55292 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output525
timestamp 1623939100
transform -1 0 55660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output518
timestamp 1623939100
transform 1 0 54924 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_601
timestamp 1623939100
transform 1 0 56396 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_593
timestamp 1623939100
transform 1 0 55660 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_597
timestamp 1623939100
transform 1 0 56028 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output521
timestamp 1623939100
transform 1 0 56396 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output520
timestamp 1623939100
transform 1 0 55660 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output527
timestamp 1623939100
transform 1 0 56580 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_607
timestamp 1623939100
transform 1 0 56948 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_610
timestamp 1623939100
transform 1 0 57224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_605
timestamp 1623939100
transform 1 0 56764 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1623939100
transform 1 0 57316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1623939100
transform 1 0 57132 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_614
timestamp 1623939100
transform 1 0 57592 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_324
timestamp 1623939100
transform -1 0 57592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output523
timestamp 1623939100
transform -1 0 57960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_621
timestamp 1623939100
transform 1 0 58236 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_618
timestamp 1623939100
transform 1 0 57960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_325
timestamp 1623939100
transform -1 0 58328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output524
timestamp 1623939100
transform -1 0 58696 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input121
timestamp 1623939100
transform 1 0 57960 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_628
timestamp 1623939100
transform 1 0 58880 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_626
timestamp 1623939100
transform 1 0 58696 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1623939100
transform 1 0 58788 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_634
timestamp 1623939100
transform 1 0 59432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output532
timestamp 1623939100
transform 1 0 59248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output526
timestamp 1623939100
transform 1 0 59064 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_636
timestamp 1623939100
transform 1 0 59616 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_639
timestamp 1623939100
transform 1 0 59892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1623939100
transform 1 0 59800 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_643
timestamp 1623939100
transform 1 0 60260 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_328
timestamp 1623939100
transform -1 0 60260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output528
timestamp 1623939100
transform -1 0 60628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input125
timestamp 1623939100
transform 1 0 59984 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_650
timestamp 1623939100
transform 1 0 60904 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_647
timestamp 1623939100
transform 1 0 60628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_330
timestamp 1623939100
transform -1 0 60996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output529
timestamp 1623939100
transform -1 0 61364 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input126
timestamp 1623939100
transform 1 0 60628 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_660
timestamp 1623939100
transform 1 0 61824 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_663
timestamp 1623939100
transform 1 0 62100 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_655
timestamp 1623939100
transform 1 0 61364 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_333
timestamp 1623939100
transform -1 0 61732 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output536
timestamp 1623939100
transform 1 0 61456 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output531
timestamp 1623939100
transform -1 0 62100 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_668
timestamp 1623939100
transform 1 0 62560 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_668
timestamp 1623939100
transform 1 0 62560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_335
timestamp 1623939100
transform -1 0 62928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output538
timestamp 1623939100
transform 1 0 62652 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1623939100
transform 1 0 62468 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_673
timestamp 1623939100
transform 1 0 63020 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_676
timestamp 1623939100
transform 1 0 63296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output533
timestamp 1623939100
transform -1 0 63296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_680
timestamp 1623939100
transform 1 0 63664 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output534
timestamp 1623939100
transform 1 0 63664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _684_
timestamp 1623939100
transform 1 0 63388 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_685
timestamp 1623939100
transform 1 0 64124 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_684
timestamp 1623939100
transform 1 0 64032 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1623939100
transform 1 0 64032 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_342
timestamp 1623939100
transform -1 0 64492 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_693
timestamp 1623939100
transform 1 0 64860 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_692
timestamp 1623939100
transform 1 0 64768 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output542
timestamp 1623939100
transform -1 0 64860 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output535
timestamp 1623939100
transform 1 0 64400 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_700
timestamp 1623939100
transform 1 0 65504 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_697
timestamp 1623939100
transform 1 0 65228 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output537
timestamp 1623939100
transform 1 0 65596 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input134
timestamp 1623939100
transform 1 0 65228 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1623939100
transform 1 0 65136 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_707
timestamp 1623939100
transform 1 0 66148 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_705
timestamp 1623939100
transform 1 0 65964 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_337
timestamp 1623939100
transform -1 0 66332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input136
timestamp 1623939100
transform 1 0 65872 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_346
timestamp 1623939100
transform -1 0 66884 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_338
timestamp 1623939100
transform -1 0 66884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output539
timestamp 1623939100
transform -1 0 66700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_340
timestamp 1623939100
transform -1 0 67068 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output546
timestamp 1623939100
transform -1 0 67252 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output540
timestamp 1623939100
transform -1 0 67436 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_719
timestamp 1623939100
transform 1 0 67252 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_341
timestamp 1623939100
transform -1 0 67620 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_726
timestamp 1623939100
transform 1 0 67896 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_726
timestamp 1623939100
transform 1 0 67896 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_723
timestamp 1623939100
transform 1 0 67620 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1623939100
transform 1 0 67620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1623939100
transform 1 0 67804 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_344
timestamp 1623939100
transform -1 0 68264 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_733
timestamp 1623939100
transform 1 0 68540 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_734
timestamp 1623939100
transform 1 0 68632 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_345
timestamp 1623939100
transform -1 0 69000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output544
timestamp 1623939100
transform -1 0 69368 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output543
timestamp 1623939100
transform -1 0 68632 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input139
timestamp 1623939100
transform 1 0 68264 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_742
timestamp 1623939100
transform 1 0 69368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_742
timestamp 1623939100
transform 1 0 69368 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_350
timestamp 1623939100
transform -1 0 69736 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output550
timestamp 1623939100
transform -1 0 70104 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output545
timestamp 1623939100
transform 1 0 69736 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1623939100
transform 1 0 69276 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_750
timestamp 1623939100
transform 1 0 70104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_750
timestamp 1623939100
transform 1 0 70104 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 71300 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1623939100
transform 1 0 70472 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output547
timestamp 1623939100
transform 1 0 70932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output548
timestamp 1623939100
transform 1 0 71668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output553
timestamp 1623939100
transform -1 0 70932 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_352
timestamp 1623939100
transform -1 0 70564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_755
timestamp 1623939100
transform 1 0 70564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_763
timestamp 1623939100
transform 1 0 71300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_759
timestamp 1623939100
transform 1 0 70932 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_772
timestamp 1623939100
transform 1 0 72128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_771
timestamp 1623939100
transform 1 0 72036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_348
timestamp 1623939100
transform -1 0 72404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output549
timestamp 1623939100
transform -1 0 72772 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_780
timestamp 1623939100
transform 1 0 72864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_779
timestamp 1623939100
transform 1 0 72772 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output556
timestamp 1623939100
transform 1 0 72496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_784
timestamp 1623939100
transform 1 0 73232 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1623939100
transform 1 0 73232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1623939100
transform 1 0 73140 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_787
timestamp 1623939100
transform 1 0 73508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output551
timestamp 1623939100
transform 1 0 73600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input150
timestamp 1623939100
transform 1 0 73876 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_794
timestamp 1623939100
transform 1 0 74152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_792
timestamp 1623939100
transform 1 0 73968 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_353
timestamp 1623939100
transform -1 0 74336 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output554
timestamp 1623939100
transform -1 0 74704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_799
timestamp 1623939100
transform 1 0 74612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_800
timestamp 1623939100
transform 1 0 74704 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_357
timestamp 1623939100
transform -1 0 74980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1623939100
transform 1 0 74520 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_355
timestamp 1623939100
transform -1 0 75072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output560
timestamp 1623939100
transform -1 0 75348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output555
timestamp 1623939100
transform -1 0 75440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_807
timestamp 1623939100
transform 1 0 75348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_808
timestamp 1623939100
transform 1 0 75440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input153
timestamp 1623939100
transform 1 0 75716 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1623939100
transform 1 0 75808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_818
timestamp 1623939100
transform 1 0 76360 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_814
timestamp 1623939100
transform 1 0 75992 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_821
timestamp 1623939100
transform 1 0 76636 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_813
timestamp 1623939100
transform 1 0 75900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_362
timestamp 1623939100
transform -1 0 76636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output564
timestamp 1623939100
transform -1 0 77004 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output557
timestamp 1623939100
transform 1 0 76268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_825
timestamp 1623939100
transform 1 0 77004 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_829
timestamp 1623939100
transform 1 0 77372 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output558
timestamp 1623939100
transform 1 0 77004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_833
timestamp 1623939100
transform 1 0 77740 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output559
timestamp 1623939100
transform 1 0 77740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_839
timestamp 1623939100
transform 1 0 78292 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_842
timestamp 1623939100
transform 1 0 78568 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_837
timestamp 1623939100
transform 1 0 78108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_365
timestamp 1623939100
transform -1 0 78660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output566
timestamp 1623939100
transform 1 0 77924 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1623939100
transform 1 0 78476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_847
timestamp 1623939100
transform 1 0 79028 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_850
timestamp 1623939100
transform 1 0 79304 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_358
timestamp 1623939100
transform -1 0 78936 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output567
timestamp 1623939100
transform -1 0 79028 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output561
timestamp 1623939100
transform -1 0 79304 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_360
timestamp 1623939100
transform -1 0 79672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output562
timestamp 1623939100
transform -1 0 80040 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_856
timestamp 1623939100
transform 1 0 79856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_858
timestamp 1623939100
transform 1 0 80040 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_369
timestamp 1623939100
transform -1 0 80224 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_363
timestamp 1623939100
transform -1 0 80408 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output569
timestamp 1623939100
transform -1 0 80592 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1623939100
transform 1 0 79764 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_864
timestamp 1623939100
transform 1 0 80592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_866
timestamp 1623939100
transform 1 0 80776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_371
timestamp 1623939100
transform -1 0 80960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output565
timestamp 1623939100
transform -1 0 80776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_872
timestamp 1623939100
transform 1 0 81328 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_871
timestamp 1623939100
transform 1 0 81236 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_372
timestamp 1623939100
transform -1 0 81696 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output570
timestamp 1623939100
transform -1 0 81328 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1623939100
transform 1 0 81144 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_880
timestamp 1623939100
transform 1 0 82064 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_877
timestamp 1623939100
transform 1 0 81788 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_257
timestamp 1623939100
transform 1 0 81880 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output571
timestamp 1623939100
transform -1 0 82064 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output449
timestamp 1623939100
transform 1 0 82064 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_888
timestamp 1623939100
transform 1 0 82800 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_884
timestamp 1623939100
transform 1 0 82432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_255
timestamp 1623939100
transform -1 0 82800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output573
timestamp 1623939100
transform 1 0 82432 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output448
timestamp 1623939100
transform -1 0 83168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_895
timestamp 1623939100
transform 1 0 83444 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_892
timestamp 1623939100
transform 1 0 83168 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1623939100
transform 1 0 83168 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_902
timestamp 1623939100
transform 1 0 84088 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_904
timestamp 1623939100
transform 1 0 84272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_900
timestamp 1623939100
transform 1 0 83904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_898
timestamp 1623939100
transform 1 0 83720 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1623939100
transform 1 0 83812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1623939100
transform 1 0 83812 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_913
timestamp 1623939100
transform 1 0 85100 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_910
timestamp 1623939100
transform 1 0 84824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1623939100
transform 1 0 85008 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 84364 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_925
timestamp 1623939100
transform 1 0 86204 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_924
timestamp 1623939100
transform 1 0 86112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_263
timestamp 1623939100
transform -1 0 85836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output453
timestamp 1623939100
transform -1 0 86204 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_932
timestamp 1623939100
transform 1 0 86848 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_929
timestamp 1623939100
transform 1 0 86572 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output450
timestamp 1623939100
transform 1 0 86940 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1623939100
transform 1 0 86572 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1623939100
transform 1 0 86480 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_937
timestamp 1623939100
transform 1 0 87308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_940
timestamp 1623939100
transform 1 0 87584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_945
timestamp 1623939100
transform 1 0 88044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_260
timestamp 1623939100
transform -1 0 88412 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output451
timestamp 1623939100
transform 1 0 87676 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_958
timestamp 1623939100
transform 1 0 89240 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_955
timestamp 1623939100
transform 1 0 88964 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_261
timestamp 1623939100
transform -1 0 88964 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output452
timestamp 1623939100
transform -1 0 88780 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1623939100
transform 1 0 89148 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _739_
timestamp 1623939100
transform 1 0 87676 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_1_960
timestamp 1623939100
transform 1 0 89424 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_966
timestamp 1623939100
transform 1 0 89976 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_265
timestamp 1623939100
transform -1 0 89608 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output454
timestamp 1623939100
transform -1 0 89976 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_970
timestamp 1623939100
transform 1 0 90344 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_968
timestamp 1623939100
transform 1 0 90160 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_974
timestamp 1623939100
transform 1 0 90712 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_275
timestamp 1623939100
transform -1 0 90712 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_269
timestamp 1623939100
transform -1 0 91080 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_267
timestamp 1623939100
transform -1 0 90344 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output461
timestamp 1623939100
transform -1 0 91080 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output455
timestamp 1623939100
transform -1 0 90712 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1623939100
transform 1 0 90252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_978
timestamp 1623939100
transform 1 0 91080 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output456
timestamp 1623939100
transform -1 0 91448 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_982
timestamp 1623939100
transform 1 0 91448 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output462
timestamp 1623939100
transform 1 0 91448 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_986
timestamp 1623939100
transform 1 0 91816 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_987
timestamp 1623939100
transform 1 0 91908 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_271
timestamp 1623939100
transform -1 0 92276 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1623939100
transform 1 0 91816 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output464
timestamp 1623939100
transform 1 0 92184 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output457
timestamp 1623939100
transform -1 0 92644 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_994
timestamp 1623939100
transform 1 0 92552 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_995
timestamp 1623939100
transform 1 0 92644 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_279
timestamp 1623939100
transform -1 0 93104 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output466
timestamp 1623939100
transform -1 0 93472 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output459
timestamp 1623939100
transform 1 0 93012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1004
timestamp 1623939100
transform 1 0 93472 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1003
timestamp 1623939100
transform 1 0 93380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output460
timestamp 1623939100
transform 1 0 93748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1012
timestamp 1623939100
transform 1 0 94208 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1011
timestamp 1623939100
transform 1 0 94116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output467
timestamp 1623939100
transform 1 0 93840 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1020
timestamp 1623939100
transform 1 0 94944 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1016
timestamp 1623939100
transform 1 0 94576 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_281
timestamp 1623939100
transform -1 0 94576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_277
timestamp 1623939100
transform -1 0 94944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output468
timestamp 1623939100
transform -1 0 94944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output463
timestamp 1623939100
transform -1 0 95312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1623939100
transform 1 0 94484 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1024
timestamp 1623939100
transform 1 0 95312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1027
timestamp 1623939100
transform 1 0 95588 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_284
timestamp 1623939100
transform -1 0 95956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output465
timestamp 1623939100
transform 1 0 95680 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1623939100
transform 1 0 95496 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1035
timestamp 1623939100
transform 1 0 96324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1032
timestamp 1623939100
transform 1 0 96048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_249
timestamp 1623939100
transform 1 0 96232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output471
timestamp 1623939100
transform -1 0 96324 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1040
timestamp 1623939100
transform 1 0 96784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_285
timestamp 1623939100
transform -1 0 96692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output472
timestamp 1623939100
transform -1 0 97060 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output445
timestamp 1623939100
transform 1 0 96416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1043
timestamp 1623939100
transform 1 0 97060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1045
timestamp 1623939100
transform 1 0 97244 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_286
timestamp 1623939100
transform -1 0 97428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output473
timestamp 1623939100
transform -1 0 97796 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1623939100
transform 1 0 97152 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1051
timestamp 1623939100
transform 1 0 97796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1055
timestamp 1623939100
transform 1 0 98164 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output444
timestamp 1623939100
transform 1 0 97796 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1623939100
transform -1 0 98808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1623939100
transform -1 0 98808 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1623939100
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input297
timestamp 1623939100
transform 1 0 2760 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input308
timestamp 1623939100
transform 1 0 1840 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1623939100
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1623939100
transform 1 0 1748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1623939100
transform 1 0 2392 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1623939100
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input355
timestamp 1623939100
transform 1 0 4232 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1623939100
transform 1 0 3312 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_28
timestamp 1623939100
transform 1 0 3680 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_30
timestamp 1623939100
transform 1 0 3864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_40
timestamp 1623939100
transform 1 0 4784 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  _436_
timestamp 1623939100
transform 1 0 5520 0 -1 3808
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_2_59
timestamp 1623939100
transform 1 0 6532 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input357
timestamp 1623939100
transform 1 0 6900 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input360
timestamp 1623939100
transform 1 0 7820 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_69
timestamp 1623939100
transform 1 0 7452 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_79
timestamp 1623939100
transform 1 0 8372 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1623939100
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output578
timestamp 1623939100
transform 1 0 9476 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output579
timestamp 1623939100
transform 1 0 10212 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1623939100
transform 1 0 8924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1623939100
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_95
timestamp 1623939100
transform 1 0 9844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_103
timestamp 1623939100
transform 1 0 10580 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output580
timestamp 1623939100
transform 1 0 10948 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output581
timestamp 1623939100
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output582
timestamp 1623939100
transform 1 0 12420 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_111
timestamp 1623939100
transform 1 0 11316 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1623939100
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1623939100
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output584
timestamp 1623939100
transform 1 0 13156 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_127
timestamp 1623939100
transform 1 0 12788 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1623939100
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1623939100
transform 1 0 14352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output586
timestamp 1623939100
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output588
timestamp 1623939100
transform 1 0 15456 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output590
timestamp 1623939100
transform 1 0 16192 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_152
timestamp 1623939100
transform 1 0 15088 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_160
timestamp 1623939100
transform 1 0 15824 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output591
timestamp 1623939100
transform -1 0 17296 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output592
timestamp 1623939100
transform -1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_382
timestamp 1623939100
transform -1 0 16928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_384
timestamp 1623939100
transform -1 0 17664 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_168
timestamp 1623939100
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_176
timestamp 1623939100
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1623939100
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1623939100
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output593
timestamp 1623939100
transform 1 0 18400 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output596
timestamp 1623939100
transform 1 0 19964 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_192
timestamp 1623939100
transform 1 0 18768 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1623939100
transform 1 0 19596 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1623939100
transform 1 0 22172 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output597
timestamp 1623939100
transform 1 0 20700 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output599
timestamp 1623939100
transform 1 0 21436 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1623939100
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_217
timestamp 1623939100
transform 1 0 21068 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_225
timestamp 1623939100
transform 1 0 21804 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1623939100
transform 1 0 22816 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 1623939100
transform 1 0 24012 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_232
timestamp 1623939100
transform 1 0 22448 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_239
timestamp 1623939100
transform 1 0 23092 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_247
timestamp 1623939100
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1623939100
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input122
timestamp 1623939100
transform 1 0 25208 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input133
timestamp 1623939100
transform 1 0 25852 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_252
timestamp 1623939100
transform 1 0 24288 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_256
timestamp 1623939100
transform 1 0 24656 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1623939100
transform 1 0 24840 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1623939100
transform 1 0 25484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1623939100
transform 1 0 27692 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output563
timestamp 1623939100
transform 1 0 26680 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_272
timestamp 1623939100
transform 1 0 26128 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_282
timestamp 1623939100
transform 1 0 27048 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_288
timestamp 1623939100
transform 1 0 27600 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1623939100
transform 1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_292
timestamp 1623939100
transform 1 0 27968 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_300
timestamp 1623939100
transform 1 0 28704 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_305
timestamp 1623939100
transform 1 0 29164 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1623939100
transform 1 0 29992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input199
timestamp 1623939100
transform 1 0 30452 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input200
timestamp 1623939100
transform 1 0 31096 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_313
timestamp 1623939100
transform 1 0 29900 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_315
timestamp 1623939100
transform 1 0 30084 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp 1623939100
transform 1 0 30728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_329
timestamp 1623939100
transform 1 0 31372 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 1623939100
transform 1 0 31924 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input202
timestamp 1623939100
transform 1 0 32568 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input203
timestamp 1623939100
transform 1 0 33212 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_338
timestamp 1623939100
transform 1 0 32200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_345
timestamp 1623939100
transform 1 0 32844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_352
timestamp 1623939100
transform 1 0 33488 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1623939100
transform 1 0 35236 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 1623939100
transform 1 0 34408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_360
timestamp 1623939100
transform 1 0 34224 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_365
timestamp 1623939100
transform 1 0 34684 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_372
timestamp 1623939100
transform 1 0 35328 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 37352 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1623939100
transform 1 0 35696 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 1623939100
transform 1 0 36340 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_379
timestamp 1623939100
transform 1 0 35972 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_386
timestamp 1623939100
transform 1 0 36616 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1623939100
transform 1 0 38916 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_407
timestamp 1623939100
transform 1 0 38548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_414
timestamp 1623939100
transform 1 0 39192 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1623939100
transform 1 0 40480 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1623939100
transform 1 0 39560 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1623939100
transform 1 0 40940 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_421
timestamp 1623939100
transform 1 0 39836 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_427
timestamp 1623939100
transform 1 0 40388 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_429
timestamp 1623939100
transform 1 0 40572 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_436
timestamp 1623939100
transform 1 0 41216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1623939100
transform 1 0 41676 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input94
timestamp 1623939100
transform 1 0 42320 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input95
timestamp 1623939100
transform 1 0 42964 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_440
timestamp 1623939100
transform 1 0 41584 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_444
timestamp 1623939100
transform 1 0 41952 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_451
timestamp 1623939100
transform 1 0 42596 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_458
timestamp 1623939100
transform 1 0 43240 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 1623939100
transform 1 0 44804 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input221
timestamp 1623939100
transform 1 0 43608 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_465
timestamp 1623939100
transform 1 0 43884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_473
timestamp 1623939100
transform 1 0 44620 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_478
timestamp 1623939100
transform 1 0 45080 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _620_
timestamp 1623939100
transform 1 0 46552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1623939100
transform 1 0 45724 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_484
timestamp 1623939100
transform 1 0 45632 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_486
timestamp 1623939100
transform 1 0 45816 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_497
timestamp 1623939100
transform 1 0 46828 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 1623939100
transform 1 0 47196 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input103
timestamp 1623939100
transform 1 0 47840 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input104
timestamp 1623939100
transform 1 0 48484 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_504
timestamp 1623939100
transform 1 0 47472 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_511
timestamp 1623939100
transform 1 0 48116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_518
timestamp 1623939100
transform 1 0 48760 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input105
timestamp 1623939100
transform 1 0 49128 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input107
timestamp 1623939100
transform 1 0 49772 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_525
timestamp 1623939100
transform 1 0 49404 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_532
timestamp 1623939100
transform 1 0 50048 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_540
timestamp 1623939100
transform 1 0 50784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1623939100
transform 1 0 50968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input109
timestamp 1623939100
transform 1 0 51428 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input112
timestamp 1623939100
transform 1 0 52072 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1623939100
transform 1 0 52716 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_543
timestamp 1623939100
transform 1 0 51060 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_550
timestamp 1623939100
transform 1 0 51704 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_557
timestamp 1623939100
transform 1 0 52348 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input114
timestamp 1623939100
transform 1 0 53360 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input115
timestamp 1623939100
transform 1 0 54004 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input116
timestamp 1623939100
transform 1 0 54648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_564
timestamp 1623939100
transform 1 0 52992 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_571
timestamp 1623939100
transform 1 0 53636 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_578
timestamp 1623939100
transform 1 0 54280 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1623939100
transform 1 0 56212 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input117
timestamp 1623939100
transform 1 0 55292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input119
timestamp 1623939100
transform 1 0 56672 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_585
timestamp 1623939100
transform 1 0 54924 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_592
timestamp 1623939100
transform 1 0 55568 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_598
timestamp 1623939100
transform 1 0 56120 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_600
timestamp 1623939100
transform 1 0 56304 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input120
timestamp 1623939100
transform 1 0 57316 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input123
timestamp 1623939100
transform 1 0 58144 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_607
timestamp 1623939100
transform 1 0 56948 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_614
timestamp 1623939100
transform 1 0 57592 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_623
timestamp 1623939100
transform 1 0 58420 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input124
timestamp 1623939100
transform 1 0 58788 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input249
timestamp 1623939100
transform 1 0 59432 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_630
timestamp 1623939100
transform 1 0 59064 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_637
timestamp 1623939100
transform 1 0 59708 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_645
timestamp 1623939100
transform 1 0 60444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1623939100
transform 1 0 61456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input127
timestamp 1623939100
transform 1 0 60628 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input128
timestamp 1623939100
transform 1 0 61916 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_650
timestamp 1623939100
transform 1 0 60904 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_657
timestamp 1623939100
transform 1 0 61548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_664
timestamp 1623939100
transform 1 0 62192 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input129
timestamp 1623939100
transform 1 0 62560 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input130
timestamp 1623939100
transform 1 0 63204 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input131
timestamp 1623939100
transform 1 0 63848 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_671
timestamp 1623939100
transform 1 0 62836 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_678
timestamp 1623939100
transform 1 0 63480 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_685
timestamp 1623939100
transform 1 0 64124 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input132
timestamp 1623939100
transform 1 0 64492 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input135
timestamp 1623939100
transform 1 0 65136 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input260
timestamp 1623939100
transform 1 0 65780 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_692
timestamp 1623939100
transform 1 0 64768 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_699
timestamp 1623939100
transform 1 0 65412 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_706
timestamp 1623939100
transform 1 0 66056 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1623939100
transform 1 0 66700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1623939100
transform 1 0 67160 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input140
timestamp 1623939100
transform 1 0 67896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_712
timestamp 1623939100
transform 1 0 66608 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_714
timestamp 1623939100
transform 1 0 66792 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_721
timestamp 1623939100
transform 1 0 67436 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_725
timestamp 1623939100
transform 1 0 67804 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_729
timestamp 1623939100
transform 1 0 68172 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1623939100
transform 1 0 68540 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1623939100
transform 1 0 69184 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input143
timestamp 1623939100
transform 1 0 69828 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_736
timestamp 1623939100
transform 1 0 68816 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_743
timestamp 1623939100
transform 1 0 69460 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_750
timestamp 1623939100
transform 1 0 70104 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1623939100
transform 1 0 71944 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input145
timestamp 1623939100
transform 1 0 70472 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input146
timestamp 1623939100
transform 1 0 71116 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_757
timestamp 1623939100
transform 1 0 70748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_764
timestamp 1623939100
transform 1 0 71392 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input147
timestamp 1623939100
transform 1 0 72404 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input149
timestamp 1623939100
transform 1 0 73048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_771
timestamp 1623939100
transform 1 0 72036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_778
timestamp 1623939100
transform 1 0 72680 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_785
timestamp 1623939100
transform 1 0 73324 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input151
timestamp 1623939100
transform 1 0 74060 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input152
timestamp 1623939100
transform 1 0 74704 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_796
timestamp 1623939100
transform 1 0 74336 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_803
timestamp 1623939100
transform 1 0 74980 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_811
timestamp 1623939100
transform 1 0 75716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _595_
timestamp 1623939100
transform 1 0 77648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1623939100
transform 1 0 77188 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input154
timestamp 1623939100
transform 1 0 75900 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input156
timestamp 1623939100
transform 1 0 76544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_816
timestamp 1623939100
transform 1 0 76176 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_823
timestamp 1623939100
transform 1 0 76820 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_828
timestamp 1623939100
transform 1 0 77280 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input158
timestamp 1623939100
transform 1 0 78292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output568
timestamp 1623939100
transform -1 0 79488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_367
timestamp 1623939100
transform -1 0 79120 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_835
timestamp 1623939100
transform 1 0 77924 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_842
timestamp 1623939100
transform 1 0 78568 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_852
timestamp 1623939100
transform 1 0 79488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input161
timestamp 1623939100
transform 1 0 79856 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input162
timestamp 1623939100
transform 1 0 80500 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output572
timestamp 1623939100
transform -1 0 81880 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_374
timestamp 1623939100
transform -1 0 81512 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_859
timestamp 1623939100
transform 1 0 80132 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_866
timestamp 1623939100
transform 1 0 80776 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1623939100
transform 1 0 82432 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input168
timestamp 1623939100
transform 1 0 82984 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_878
timestamp 1623939100
transform 1 0 81880 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_885
timestamp 1623939100
transform 1 0 82524 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_889
timestamp 1623939100
transform 1 0 82892 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_893
timestamp 1623939100
transform 1 0 83260 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _579_
timestamp 1623939100
transform 1 0 83628 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1623939100
transform 1 0 84272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1623939100
transform 1 0 84916 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_900
timestamp 1623939100
transform 1 0 83904 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_907
timestamp 1623939100
transform 1 0 84548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_914
timestamp 1623939100
transform 1 0 85192 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1623939100
transform 1 0 85560 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1623939100
transform 1 0 86204 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1623939100
transform 1 0 86848 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_921
timestamp 1623939100
transform 1 0 85836 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_928
timestamp 1623939100
transform 1 0 86480 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_935
timestamp 1623939100
transform 1 0 87124 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1623939100
transform 1 0 87676 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1623939100
transform 1 0 88136 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1623939100
transform 1 0 88780 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_942
timestamp 1623939100
transform 1 0 87768 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_949
timestamp 1623939100
transform 1 0 88412 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_956
timestamp 1623939100
transform 1 0 89056 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1623939100
transform 1 0 89424 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1623939100
transform 1 0 90068 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1623939100
transform 1 0 90712 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_963
timestamp 1623939100
transform 1 0 89700 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_970
timestamp 1623939100
transform 1 0 90344 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_977
timestamp 1623939100
transform 1 0 90988 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1623939100
transform 1 0 92920 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1623939100
transform 1 0 91356 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1623939100
transform 1 0 92000 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_984
timestamp 1623939100
transform 1 0 91632 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_991
timestamp 1623939100
transform 1 0 92276 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_997
timestamp 1623939100
transform 1 0 92828 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_999
timestamp 1623939100
transform 1 0 93012 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1623939100
transform 1 0 93380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1623939100
transform 1 0 94024 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output470
timestamp 1623939100
transform -1 0 95312 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_283
timestamp 1623939100
transform -1 0 94944 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1006
timestamp 1623939100
transform 1 0 93656 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1013
timestamp 1623939100
transform 1 0 94300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1017
timestamp 1623939100
transform 1 0 94668 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1623939100
transform 1 0 95680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output476
timestamp 1623939100
transform 1 0 96692 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_290
timestamp 1623939100
transform 1 0 96508 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1024
timestamp 1623939100
transform 1 0 95312 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1031
timestamp 1623939100
transform 1 0 95956 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1623939100
transform -1 0 98808 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1623939100
transform 1 0 98164 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output474
timestamp 1623939100
transform 1 0 97428 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1043
timestamp 1623939100
transform 1 0 97060 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1051
timestamp 1623939100
transform 1 0 97796 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1056
timestamp 1623939100
transform 1 0 98256 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1623939100
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input329
timestamp 1623939100
transform 1 0 1748 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input367
timestamp 1623939100
transform 1 0 2668 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1623939100
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1623939100
transform 1 0 2300 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input352
timestamp 1623939100
transform 1 0 3588 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input356
timestamp 1623939100
transform 1 0 4692 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output598
timestamp 1623939100
transform 1 0 4232 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_23
timestamp 1623939100
transform 1 0 3220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_31
timestamp 1623939100
transform 1 0 3956 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_38
timestamp 1623939100
transform 1 0 4600 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1623939100
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input359
timestamp 1623939100
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output602
timestamp 1623939100
transform 1 0 5612 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1623939100
transform 1 0 5244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_53
timestamp 1623939100
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_58
timestamp 1623939100
transform 1 0 6440 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input361
timestamp 1623939100
transform 1 0 7728 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output577
timestamp 1623939100
transform 1 0 8556 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_66
timestamp 1623939100
transform 1 0 7176 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_76
timestamp 1623939100
transform 1 0 8096 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_80
timestamp 1623939100
transform 1 0 8464 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input300
timestamp 1623939100
transform 1 0 10028 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input301
timestamp 1623939100
transform 1 0 10672 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output607
timestamp 1623939100
transform 1 0 9292 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1623939100
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1623939100
transform 1 0 9660 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_100
timestamp 1623939100
transform 1 0 10304 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1623939100
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output583
timestamp 1623939100
transform 1 0 12236 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_107
timestamp 1623939100
transform 1 0 10948 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1623939100
transform 1 0 11500 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_115
timestamp 1623939100
transform 1 0 11684 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_125
timestamp 1623939100
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _662_
timestamp 1623939100
transform 1 0 12972 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input306
timestamp 1623939100
transform 1 0 13616 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input307
timestamp 1623939100
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_366
timestamp 1623939100
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1623939100
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1623939100
transform 1 0 13892 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input311
timestamp 1623939100
transform 1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output589
timestamp 1623939100
transform 1 0 15272 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_146
timestamp 1623939100
transform 1 0 14536 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_158
timestamp 1623939100
transform 1 0 15640 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_165
timestamp 1623939100
transform 1 0 16284 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1623939100
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input313
timestamp 1623939100
transform 1 0 17296 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output594
timestamp 1623939100
transform 1 0 18308 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1623939100
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_179
timestamp 1623939100
transform 1 0 17572 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _574_
timestamp 1623939100
transform 1 0 19780 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output595
timestamp 1623939100
transform 1 0 19044 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_191
timestamp 1623939100
transform 1 0 18676 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_199
timestamp 1623939100
transform 1 0 19412 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_206
timestamp 1623939100
transform 1 0 20056 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1623939100
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input317
timestamp 1623939100
transform 1 0 20424 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input320
timestamp 1623939100
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1623939100
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_220
timestamp 1623939100
transform 1 0 21344 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_229
timestamp 1623939100
transform 1 0 22172 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_8  _535_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 22540 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_249
timestamp 1623939100
transform 1 0 24012 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _685_
timestamp 1623939100
transform 1 0 25668 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input228
timestamp 1623939100
transform 1 0 24380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input239
timestamp 1623939100
transform 1 0 25024 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_278
timestamp 1623939100
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_256
timestamp 1623939100
transform 1 0 24656 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_263
timestamp 1623939100
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_270
timestamp 1623939100
transform 1 0 25944 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1623939100
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input144
timestamp 1623939100
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input155
timestamp 1623939100
transform 1 0 27784 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_277
timestamp 1623939100
transform 1 0 26588 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_286
timestamp 1623939100
transform 1 0 27416 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input178
timestamp 1623939100
transform 1 0 28428 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input189
timestamp 1623939100
transform 1 0 29072 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input198
timestamp 1623939100
transform 1 0 29716 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_293
timestamp 1623939100
transform 1 0 28060 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_300
timestamp 1623939100
transform 1 0 28704 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_307
timestamp 1623939100
transform 1 0 29348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input201
timestamp 1623939100
transform 1 0 31188 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_314 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 29992 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_326
timestamp 1623939100
transform 1 0 31096 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_330
timestamp 1623939100
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1623939100
transform 1 0 32568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input204
timestamp 1623939100
transform 1 0 33028 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input205
timestamp 1623939100
transform 1 0 33672 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_343
timestamp 1623939100
transform 1 0 32660 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_350
timestamp 1623939100
transform 1 0 33304 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _482_
timestamp 1623939100
transform 1 0 34316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input208
timestamp 1623939100
transform 1 0 35512 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_357
timestamp 1623939100
transform 1 0 33948 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_370
timestamp 1623939100
transform 1 0 35144 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 1623939100
transform 1 0 36800 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input209
timestamp 1623939100
transform 1 0 36156 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_377
timestamp 1623939100
transform 1 0 35788 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_384
timestamp 1623939100
transform 1 0 36432 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_391
timestamp 1623939100
transform 1 0 37076 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1623939100
transform 1 0 37812 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 1623939100
transform 1 0 38640 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input212
timestamp 1623939100
transform 1 0 39284 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_400
timestamp 1623939100
transform 1 0 37904 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_411
timestamp 1623939100
transform 1 0 38916 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1623939100
transform 1 0 39928 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input215
timestamp 1623939100
transform 1 0 40572 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input216
timestamp 1623939100
transform 1 0 41216 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_418
timestamp 1623939100
transform 1 0 39560 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_425
timestamp 1623939100
transform 1 0 40204 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_432
timestamp 1623939100
transform 1 0 40848 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1623939100
transform 1 0 43056 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input219
timestamp 1623939100
transform 1 0 41860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_439
timestamp 1623939100
transform 1 0 41492 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_446
timestamp 1623939100
transform 1 0 42136 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_454
timestamp 1623939100
transform 1 0 42872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_457
timestamp 1623939100
transform 1 0 43148 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input222
timestamp 1623939100
transform 1 0 43516 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input223
timestamp 1623939100
transform 1 0 44160 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_464
timestamp 1623939100
transform 1 0 43792 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_471
timestamp 1623939100
transform 1 0 44436 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_479
timestamp 1623939100
transform 1 0 45172 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 1623939100
transform 1 0 45356 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 1623939100
transform 1 0 46000 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input226
timestamp 1623939100
transform 1 0 46644 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_484
timestamp 1623939100
transform 1 0 45632 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_491
timestamp 1623939100
transform 1 0 46276 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_498
timestamp 1623939100
transform 1 0 46920 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1623939100
transform 1 0 48300 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input229
timestamp 1623939100
transform 1 0 47288 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input232
timestamp 1623939100
transform 1 0 48760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_505
timestamp 1623939100
transform 1 0 47564 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_514
timestamp 1623939100
transform 1 0 48392 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input233
timestamp 1623939100
transform 1 0 49404 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input234
timestamp 1623939100
transform 1 0 50048 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input235
timestamp 1623939100
transform 1 0 50692 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_521
timestamp 1623939100
transform 1 0 49036 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_528
timestamp 1623939100
transform 1 0 49680 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_535
timestamp 1623939100
transform 1 0 50324 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input236
timestamp 1623939100
transform 1 0 51336 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input237
timestamp 1623939100
transform 1 0 51980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input238
timestamp 1623939100
transform 1 0 52624 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_542
timestamp 1623939100
transform 1 0 50968 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_549
timestamp 1623939100
transform 1 0 51612 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_556
timestamp 1623939100
transform 1 0 52256 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1623939100
transform 1 0 53544 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input241
timestamp 1623939100
transform 1 0 54004 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input242
timestamp 1623939100
transform 1 0 54648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_563
timestamp 1623939100
transform 1 0 52900 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_569
timestamp 1623939100
transform 1 0 53452 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_571
timestamp 1623939100
transform 1 0 53636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_578
timestamp 1623939100
transform 1 0 54280 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input244
timestamp 1623939100
transform 1 0 55292 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input245
timestamp 1623939100
transform 1 0 55936 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input246
timestamp 1623939100
transform 1 0 56580 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_585
timestamp 1623939100
transform 1 0 54924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_592
timestamp 1623939100
transform 1 0 55568 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_599
timestamp 1623939100
transform 1 0 56212 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input247
timestamp 1623939100
transform 1 0 57224 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input248
timestamp 1623939100
transform 1 0 57868 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_606
timestamp 1623939100
transform 1 0 56856 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_613
timestamp 1623939100
transform 1 0 57500 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_620
timestamp 1623939100
transform 1 0 58144 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1623939100
transform 1 0 58788 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input251
timestamp 1623939100
transform 1 0 59248 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input252
timestamp 1623939100
transform 1 0 59892 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_626
timestamp 1623939100
transform 1 0 58696 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_628
timestamp 1623939100
transform 1 0 58880 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_635
timestamp 1623939100
transform 1 0 59524 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_642
timestamp 1623939100
transform 1 0 60168 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input253
timestamp 1623939100
transform 1 0 60536 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input254
timestamp 1623939100
transform 1 0 61180 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input255
timestamp 1623939100
transform 1 0 61824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_649
timestamp 1623939100
transform 1 0 60812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_656
timestamp 1623939100
transform 1 0 61456 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_663
timestamp 1623939100
transform 1 0 62100 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1623939100
transform 1 0 64032 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input256
timestamp 1623939100
transform 1 0 62468 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input257
timestamp 1623939100
transform 1 0 63112 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_670
timestamp 1623939100
transform 1 0 62744 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_677
timestamp 1623939100
transform 1 0 63388 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_683
timestamp 1623939100
transform 1 0 63940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_685
timestamp 1623939100
transform 1 0 64124 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input258
timestamp 1623939100
transform 1 0 64492 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input259
timestamp 1623939100
transform 1 0 65136 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input262
timestamp 1623939100
transform 1 0 65780 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_692
timestamp 1623939100
transform 1 0 64768 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_699
timestamp 1623939100
transform 1 0 65412 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_706
timestamp 1623939100
transform 1 0 66056 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input263
timestamp 1623939100
transform 1 0 66424 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input265
timestamp 1623939100
transform 1 0 67068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input266
timestamp 1623939100
transform 1 0 67712 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_713
timestamp 1623939100
transform 1 0 66700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_720
timestamp 1623939100
transform 1 0 67344 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_727
timestamp 1623939100
transform 1 0 67988 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1623939100
transform 1 0 69276 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input267
timestamp 1623939100
transform 1 0 68356 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input269
timestamp 1623939100
transform 1 0 69736 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_734
timestamp 1623939100
transform 1 0 68632 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_740
timestamp 1623939100
transform 1 0 69184 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_742
timestamp 1623939100
transform 1 0 69368 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_749
timestamp 1623939100
transform 1 0 70012 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input270
timestamp 1623939100
transform 1 0 70380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input271
timestamp 1623939100
transform 1 0 71024 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input274
timestamp 1623939100
transform 1 0 71668 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_756
timestamp 1623939100
transform 1 0 70656 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_763
timestamp 1623939100
transform 1 0 71300 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_770
timestamp 1623939100
transform 1 0 71944 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input275
timestamp 1623939100
transform 1 0 72312 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input276
timestamp 1623939100
transform 1 0 72956 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input277
timestamp 1623939100
transform 1 0 73600 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_777
timestamp 1623939100
transform 1 0 72588 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_784
timestamp 1623939100
transform 1 0 73232 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_791
timestamp 1623939100
transform 1 0 73876 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1623939100
transform 1 0 74520 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input279
timestamp 1623939100
transform 1 0 74980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input280
timestamp 1623939100
transform 1 0 75624 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_797
timestamp 1623939100
transform 1 0 74428 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_799
timestamp 1623939100
transform 1 0 74612 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_806
timestamp 1623939100
transform 1 0 75256 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input157
timestamp 1623939100
transform 1 0 77096 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input281
timestamp 1623939100
transform 1 0 76268 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_813
timestamp 1623939100
transform 1 0 75900 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_820
timestamp 1623939100
transform 1 0 76544 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_829
timestamp 1623939100
transform 1 0 77372 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input159
timestamp 1623939100
transform 1 0 78292 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input160
timestamp 1623939100
transform 1 0 78936 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_837
timestamp 1623939100
transform 1 0 78108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_842
timestamp 1623939100
transform 1 0 78568 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_849
timestamp 1623939100
transform 1 0 79212 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1623939100
transform 1 0 79764 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input163
timestamp 1623939100
transform 1 0 80776 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input164
timestamp 1623939100
transform 1 0 81420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_856
timestamp 1623939100
transform 1 0 79856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_864
timestamp 1623939100
transform 1 0 80592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_869
timestamp 1623939100
transform 1 0 81052 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input165
timestamp 1623939100
transform 1 0 82064 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input291
timestamp 1623939100
transform 1 0 82708 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_876
timestamp 1623939100
transform 1 0 81696 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_883
timestamp 1623939100
transform 1 0 82340 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_890
timestamp 1623939100
transform 1 0 82984 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1623939100
transform 1 0 85008 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input169
timestamp 1623939100
transform 1 0 83628 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input170
timestamp 1623939100
transform 1 0 84272 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_896
timestamp 1623939100
transform 1 0 83536 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_900
timestamp 1623939100
transform 1 0 83904 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_907
timestamp 1623939100
transform 1 0 84548 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_911
timestamp 1623939100
transform 1 0 84916 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_913
timestamp 1623939100
transform 1 0 85100 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _584_
timestamp 1623939100
transform 1 0 86664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input171
timestamp 1623939100
transform 1 0 85468 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_920
timestamp 1623939100
transform 1 0 85744 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_928
timestamp 1623939100
transform 1 0 86480 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_933
timestamp 1623939100
transform 1 0 86940 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _771_
timestamp 1623939100
transform 1 0 87860 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_3_941
timestamp 1623939100
transform 1 0 87676 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_4  _530_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 91172 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1623939100
transform 1 0 90252 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1623939100
transform 1 0 90988 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_962
timestamp 1623939100
transform 1 0 89608 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_968
timestamp 1623939100
transform 1 0 90160 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_970
timestamp 1623939100
transform 1 0 90344 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_976
timestamp 1623939100
transform 1 0 90896 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1623939100
transform 1 0 93012 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_995
timestamp 1623939100
transform 1 0 92644 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1623939100
transform 1 0 93656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1623939100
transform 1 0 94300 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1002
timestamp 1623939100
transform 1 0 93288 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1009
timestamp 1623939100
transform 1 0 93932 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1016
timestamp 1623939100
transform 1 0 94576 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1623939100
transform 1 0 95496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1623939100
transform 1 0 95956 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_292
timestamp 1623939100
transform 1 0 96876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1024
timestamp 1623939100
transform 1 0 95312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1027
timestamp 1623939100
transform 1 0 95588 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1034
timestamp 1623939100
transform 1 0 96232 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1040
timestamp 1623939100
transform 1 0 96784 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1623939100
transform -1 0 98808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output475
timestamp 1623939100
transform 1 0 97796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output477
timestamp 1623939100
transform 1 0 97060 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_288
timestamp 1623939100
transform 1 0 97612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1047
timestamp 1623939100
transform 1 0 97428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1055
timestamp 1623939100
transform 1 0 98164 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1623939100
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input366
timestamp 1623939100
transform 1 0 1748 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output576
timestamp 1623939100
transform -1 0 3036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_377
timestamp 1623939100
transform -1 0 2668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1623939100
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1623939100
transform 1 0 2300 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1623939100
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1623939100
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1623939100
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1623939100
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1623939100
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1623939100
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1623939100
transform 1 0 3864 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_21
timestamp 1623939100
transform 1 0 3036 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _711_
timestamp 1623939100
transform 1 0 4968 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1623939100
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output604
timestamp 1623939100
transform -1 0 7452 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output606
timestamp 1623939100
transform 1 0 7820 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1623939100
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1623939100
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_388
timestamp 1623939100
transform -1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_77
timestamp 1623939100
transform 1 0 8188 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1623939100
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input299
timestamp 1623939100
transform 1 0 9476 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input302
timestamp 1623939100
transform 1 0 10580 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1623939100
transform 1 0 8924 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1623939100
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_94
timestamp 1623939100
transform 1 0 9752 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_102
timestamp 1623939100
transform 1 0 10488 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input303
timestamp 1623939100
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input304
timestamp 1623939100
transform 1 0 11868 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input305
timestamp 1623939100
transform 1 0 12512 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_106
timestamp 1623939100
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_113
timestamp 1623939100
transform 1 0 11500 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_120
timestamp 1623939100
transform 1 0 12144 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1623939100
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_127
timestamp 1623939100
transform 1 0 12788 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_139
timestamp 1623939100
transform 1 0 13892 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1623939100
transform 1 0 14352 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input309
timestamp 1623939100
transform 1 0 14720 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input310
timestamp 1623939100
transform 1 0 15364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input312
timestamp 1623939100
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_151
timestamp 1623939100
transform 1 0 14996 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_158
timestamp 1623939100
transform 1 0 15640 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_162
timestamp 1623939100
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_166
timestamp 1623939100
transform 1 0 16376 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input314
timestamp 1623939100
transform 1 0 17296 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input315
timestamp 1623939100
transform 1 0 17940 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_174
timestamp 1623939100
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1623939100
transform 1 0 17572 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1623939100
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1623939100
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input316
timestamp 1623939100
transform 1 0 18584 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input318
timestamp 1623939100
transform 1 0 19964 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_193
timestamp 1623939100
transform 1 0 18860 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_199
timestamp 1623939100
transform 1 0 19412 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1623939100
transform 1 0 19596 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_208
timestamp 1623939100
transform 1 0 20240 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input167
timestamp 1623939100
transform 1 0 21988 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input321
timestamp 1623939100
transform 1 0 20976 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_219
timestamp 1623939100
transform 1 0 21252 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input206
timestamp 1623939100
transform 1 0 22632 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input217
timestamp 1623939100
transform 1 0 23276 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1623939100
transform 1 0 22264 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1623939100
transform 1 0 22908 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_244
timestamp 1623939100
transform 1 0 23552 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _348_
timestamp 1623939100
transform 1 0 25668 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1623939100
transform 1 0 24748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_256
timestamp 1623939100
transform 1 0 24656 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_258
timestamp 1623939100
transform 1 0 24840 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_266
timestamp 1623939100
transform 1 0 25576 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1623939100
transform 1 0 27508 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_283
timestamp 1623939100
transform 1 0 27140 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_290
timestamp 1623939100
transform 1 0 27784 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _649_
timestamp 1623939100
transform 1 0 28428 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input294
timestamp 1623939100
transform 1 0 29072 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_296
timestamp 1623939100
transform 1 0 28336 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_300
timestamp 1623939100
transform 1 0 28704 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_307
timestamp 1623939100
transform 1 0 29348 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1623939100
transform 1 0 29992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_313
timestamp 1623939100
transform 1 0 29900 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_315
timestamp 1623939100
transform 1 0 30084 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_327
timestamp 1623939100
transform 1 0 31188 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _556_
timestamp 1623939100
transform 1 0 32936 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_214
timestamp 1623939100
transform 1 0 32752 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_339
timestamp 1623939100
transform 1 0 32292 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_343
timestamp 1623939100
transform 1 0 32660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_349
timestamp 1623939100
transform 1 0 33212 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1623939100
transform 1 0 35236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input207
timestamp 1623939100
transform 1 0 34224 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_357
timestamp 1623939100
transform 1 0 33948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_363
timestamp 1623939100
transform 1 0 34500 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_372
timestamp 1623939100
transform 1 0 35328 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _745_
timestamp 1623939100
transform 1 0 37352 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  input210
timestamp 1623939100
transform 1 0 36064 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input211
timestamp 1623939100
transform 1 0 36708 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_78
timestamp 1623939100
transform 1 0 37168 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_383
timestamp 1623939100
transform 1 0 36340 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_390
timestamp 1623939100
transform 1 0 36984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_413
timestamp 1623939100
transform 1 0 39100 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1623939100
transform 1 0 40480 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input213
timestamp 1623939100
transform 1 0 39468 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input218
timestamp 1623939100
transform 1 0 40940 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_420
timestamp 1623939100
transform 1 0 39744 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_429
timestamp 1623939100
transform 1 0 40572 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_436
timestamp 1623939100
transform 1 0 41216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _591_
timestamp 1623939100
transform 1 0 42596 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input220
timestamp 1623939100
transform 1 0 41584 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_443
timestamp 1623939100
transform 1 0 41860 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_454
timestamp 1623939100
transform 1 0 42872 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input224
timestamp 1623939100
transform 1 0 43976 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input225
timestamp 1623939100
transform 1 0 44620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_469
timestamp 1623939100
transform 1 0 44252 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_476
timestamp 1623939100
transform 1 0 44896 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1623939100
transform 1 0 45724 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input227
timestamp 1623939100
transform 1 0 46184 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input230
timestamp 1623939100
transform 1 0 47012 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_484
timestamp 1623939100
transform 1 0 45632 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_486
timestamp 1623939100
transform 1 0 45816 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_493
timestamp 1623939100
transform 1 0 46460 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input231
timestamp 1623939100
transform 1 0 47656 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_502
timestamp 1623939100
transform 1 0 47288 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_509
timestamp 1623939100
transform 1 0 47932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_521
timestamp 1623939100
transform 1 0 49036 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_533
timestamp 1623939100
transform 1 0 50140 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_541
timestamp 1623939100
transform 1 0 50876 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1623939100
transform 1 0 50968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input240
timestamp 1623939100
transform 1 0 52532 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_543
timestamp 1623939100
transform 1 0 51060 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_555
timestamp 1623939100
transform 1 0 52164 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_562
timestamp 1623939100
transform 1 0 52808 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _548_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform -1 0 53912 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  input243
timestamp 1623939100
transform 1 0 54280 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_178
timestamp 1623939100
transform -1 0 53452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_179
timestamp 1623939100
transform -1 0 54096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_566
timestamp 1623939100
transform 1 0 53176 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_576
timestamp 1623939100
transform 1 0 54096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_581
timestamp 1623939100
transform 1 0 54556 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1623939100
transform 1 0 56212 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_593
timestamp 1623939100
transform 1 0 55660 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_600
timestamp 1623939100
transform 1 0 56304 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_612
timestamp 1623939100
transform 1 0 57408 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_624
timestamp 1623939100
transform 1 0 58512 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_636
timestamp 1623939100
transform 1 0 59616 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _474_
timestamp 1623939100
transform 1 0 61916 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1623939100
transform 1 0 61456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_648
timestamp 1623939100
transform 1 0 60720 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_657
timestamp 1623939100
transform 1 0 61548 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _634_
timestamp 1623939100
transform 1 0 63296 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _748_
timestamp 1623939100
transform 1 0 63940 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_4_670
timestamp 1623939100
transform 1 0 62744 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_679
timestamp 1623939100
transform 1 0 63572 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input264
timestamp 1623939100
transform 1 0 66056 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_702
timestamp 1623939100
transform 1 0 65688 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1623939100
transform 1 0 66700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_709
timestamp 1623939100
transform 1 0 66332 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_714
timestamp 1623939100
transform 1 0 66792 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_726
timestamp 1623939100
transform 1 0 67896 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input268
timestamp 1623939100
transform 1 0 68356 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_730
timestamp 1623939100
transform 1 0 68264 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_734
timestamp 1623939100
transform 1 0 68632 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_746
timestamp 1623939100
transform 1 0 69736 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1623939100
transform 1 0 71944 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input273
timestamp 1623939100
transform 1 0 70748 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_754
timestamp 1623939100
transform 1 0 70472 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_760
timestamp 1623939100
transform 1 0 71024 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_768
timestamp 1623939100
transform 1 0 71760 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input278
timestamp 1623939100
transform 1 0 73784 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_771
timestamp 1623939100
transform 1 0 72036 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_783
timestamp 1623939100
transform 1 0 73140 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_789
timestamp 1623939100
transform 1 0 73692 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_793
timestamp 1623939100
transform 1 0 74060 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_805
timestamp 1623939100
transform 1 0 75164 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_2  _358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 77648 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1623939100
transform 1 0 77188 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input282
timestamp 1623939100
transform 1 0 76268 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_820
timestamp 1623939100
transform 1 0 76544 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_826
timestamp 1623939100
transform 1 0 77096 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_828
timestamp 1623939100
transform 1 0 77280 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input286
timestamp 1623939100
transform 1 0 78660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input287
timestamp 1623939100
transform 1 0 79304 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_839
timestamp 1623939100
transform 1 0 78292 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_846
timestamp 1623939100
transform 1 0 78936 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_853
timestamp 1623939100
transform 1 0 79580 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input288
timestamp 1623939100
transform 1 0 79948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input289
timestamp 1623939100
transform 1 0 80592 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input290
timestamp 1623939100
transform 1 0 81236 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_860
timestamp 1623939100
transform 1 0 80224 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_867
timestamp 1623939100
transform 1 0 80868 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_874
timestamp 1623939100
transform 1 0 81512 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1623939100
transform 1 0 82432 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input292
timestamp 1623939100
transform 1 0 82892 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_882
timestamp 1623939100
transform 1 0 82248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_885
timestamp 1623939100
transform 1 0 82524 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_892
timestamp 1623939100
transform 1 0 83168 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input172
timestamp 1623939100
transform 1 0 85376 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input293
timestamp 1623939100
transform 1 0 83536 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_899
timestamp 1623939100
transform 1 0 83812 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_911
timestamp 1623939100
transform 1 0 84916 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_915
timestamp 1623939100
transform 1 0 85284 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _692_
timestamp 1623939100
transform 1 0 86848 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input173
timestamp 1623939100
transform 1 0 86020 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_919
timestamp 1623939100
transform 1 0 85652 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_926
timestamp 1623939100
transform 1 0 86296 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_935
timestamp 1623939100
transform 1 0 87124 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1623939100
transform 1 0 87676 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input174
timestamp 1623939100
transform 1 0 88136 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input176
timestamp 1623939100
transform 1 0 88780 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_942
timestamp 1623939100
transform 1 0 87768 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_949
timestamp 1623939100
transform 1 0 88412 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_956
timestamp 1623939100
transform 1 0 89056 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input179
timestamp 1623939100
transform 1 0 89424 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input180
timestamp 1623939100
transform 1 0 90068 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input181
timestamp 1623939100
transform 1 0 90712 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_963
timestamp 1623939100
transform 1 0 89700 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_970
timestamp 1623939100
transform 1 0 90344 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_977
timestamp 1623939100
transform 1 0 90988 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1623939100
transform 1 0 92920 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input182
timestamp 1623939100
transform 1 0 91356 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input183
timestamp 1623939100
transform 1 0 92000 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_984
timestamp 1623939100
transform 1 0 91632 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_991
timestamp 1623939100
transform 1 0 92276 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_997
timestamp 1623939100
transform 1 0 92828 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_999
timestamp 1623939100
transform 1 0 93012 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input185
timestamp 1623939100
transform 1 0 93380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input186
timestamp 1623939100
transform 1 0 94024 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input187
timestamp 1623939100
transform 1 0 94668 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1006
timestamp 1623939100
transform 1 0 93656 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1013
timestamp 1623939100
transform 1 0 94300 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1020
timestamp 1623939100
transform 1 0 94944 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1623939100
transform 1 0 95956 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1623939100
transform 1 0 96600 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input188
timestamp 1623939100
transform 1 0 95312 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1027
timestamp 1623939100
transform 1 0 95588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1034
timestamp 1623939100
transform 1 0 96232 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1041
timestamp 1623939100
transform 1 0 96876 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1623939100
transform -1 0 98808 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1623939100
transform 1 0 98164 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1623939100
transform 1 0 97244 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1048
timestamp 1623939100
transform 1 0 97520 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1054
timestamp 1623939100
transform 1 0 98072 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1056
timestamp 1623939100
transform 1 0 98256 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _672_
timestamp 1623939100
transform 1 0 2484 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1623939100
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output575
timestamp 1623939100
transform 1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_258
timestamp 1623939100
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_259
timestamp 1623939100
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1623939100
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1623939100
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_20
timestamp 1623939100
transform 1 0 2944 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output587
timestamp 1623939100
transform 1 0 3220 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output601
timestamp 1623939100
transform 1 0 4232 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_27
timestamp 1623939100
transform 1 0 3588 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_33
timestamp 1623939100
transform 1 0 4140 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_38
timestamp 1623939100
transform 1 0 4600 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1623939100
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output603
timestamp 1623939100
transform 1 0 5520 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output605
timestamp 1623939100
transform -1 0 7176 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_389
timestamp 1623939100
transform -1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_46
timestamp 1623939100
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1623939100
transform 1 0 5888 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1623939100
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_58
timestamp 1623939100
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_6  _470_
timestamp 1623939100
transform 1 0 7912 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_66
timestamp 1623939100
transform 1 0 7176 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 1623939100
transform 1 0 8740 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input328
timestamp 1623939100
transform 1 0 9108 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_90
timestamp 1623939100
transform 1 0 9384 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_102
timestamp 1623939100
transform 1 0 10488 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _626_
timestamp 1623939100
transform 1 0 12328 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1623939100
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1623939100
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1623939100
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1623939100
transform 1 0 12604 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1623939100
transform 1 0 13708 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1623939100
transform 1 0 14812 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_161
timestamp 1623939100
transform 1 0 15916 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1623939100
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1623939100
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_172
timestamp 1623939100
transform 1 0 16928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1623939100
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1623939100
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1623939100
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1623939100
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_220
timestamp 1623939100
transform 1 0 21344 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_229
timestamp 1623939100
transform 1 0 22172 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _712_
timestamp 1623939100
transform 1 0 22908 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  input250
timestamp 1623939100
transform 1 0 25024 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input261
timestamp 1623939100
transform 1 0 25668 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_256
timestamp 1623939100
transform 1 0 24656 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_263
timestamp 1623939100
transform 1 0 25300 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_270
timestamp 1623939100
transform 1 0 25944 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1623939100
transform 1 0 27324 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input272
timestamp 1623939100
transform 1 0 26312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input283
timestamp 1623939100
transform 1 0 27784 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_277
timestamp 1623939100
transform 1 0 26588 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_286
timestamp 1623939100
transform 1 0 27416 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1623939100
transform 1 0 28060 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1623939100
transform 1 0 29164 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1623939100
transform 1 0 30268 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_329
timestamp 1623939100
transform 1 0 31372 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1623939100
transform 1 0 32568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_341
timestamp 1623939100
transform 1 0 32476 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_343
timestamp 1623939100
transform 1 0 32660 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 33764 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_5_362
timestamp 1623939100
transform 1 0 34408 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_374
timestamp 1623939100
transform 1 0 35512 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _346_
timestamp 1623939100
transform 1 0 36432 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_141
timestamp 1623939100
transform 1 0 36248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_390
timestamp 1623939100
transform 1 0 36984 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _589_
timestamp 1623939100
transform 1 0 38548 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1623939100
transform 1 0 37812 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input214
timestamp 1623939100
transform 1 0 39192 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_398
timestamp 1623939100
transform 1 0 37720 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_400
timestamp 1623939100
transform 1 0 37904 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1623939100
transform 1 0 38456 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_410
timestamp 1623939100
transform 1 0 38824 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1623939100
transform 1 0 39468 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1623939100
transform 1 0 40572 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1623939100
transform 1 0 43056 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_441
timestamp 1623939100
transform 1 0 41676 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_453
timestamp 1623939100
transform 1 0 42780 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_457
timestamp 1623939100
transform 1 0 43148 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _512_
timestamp 1623939100
transform 1 0 44804 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_469
timestamp 1623939100
transform 1 0 44252 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_484
timestamp 1623939100
transform 1 0 45632 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_496
timestamp 1623939100
transform 1 0 46736 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1623939100
transform 1 0 48300 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_508
timestamp 1623939100
transform 1 0 47840 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_512
timestamp 1623939100
transform 1 0 48208 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_514
timestamp 1623939100
transform 1 0 48392 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_526
timestamp 1623939100
transform 1 0 49496 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_538
timestamp 1623939100
transform 1 0 50600 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_550
timestamp 1623939100
transform 1 0 51704 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_562
timestamp 1623939100
transform 1 0 52808 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1623939100
transform 1 0 53544 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_571
timestamp 1623939100
transform 1 0 53636 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_583
timestamp 1623939100
transform 1 0 54740 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_595
timestamp 1623939100
transform 1 0 55844 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_607
timestamp 1623939100
transform 1 0 56948 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_619
timestamp 1623939100
transform 1 0 58052 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1623939100
transform 1 0 58788 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_628
timestamp 1623939100
transform 1 0 58880 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_640
timestamp 1623939100
transform 1 0 59984 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_652
timestamp 1623939100
transform 1 0 61088 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_664
timestamp 1623939100
transform 1 0 62192 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1623939100
transform 1 0 64032 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_676
timestamp 1623939100
transform 1 0 63296 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_685
timestamp 1623939100
transform 1 0 64124 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _304_
timestamp 1623939100
transform 1 0 64676 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_5_698
timestamp 1623939100
transform 1 0 65320 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_710
timestamp 1623939100
transform 1 0 66424 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_722
timestamp 1623939100
transform 1 0 67528 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1623939100
transform 1 0 69276 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_734
timestamp 1623939100
transform 1 0 68632 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_740
timestamp 1623939100
transform 1 0 69184 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_742
timestamp 1623939100
transform 1 0 69368 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_754
timestamp 1623939100
transform 1 0 70472 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_766
timestamp 1623939100
transform 1 0 71576 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_778
timestamp 1623939100
transform 1 0 72680 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_790
timestamp 1623939100
transform 1 0 73784 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1623939100
transform 1 0 74520 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_799
timestamp 1623939100
transform 1 0 74612 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_811
timestamp 1623939100
transform 1 0 75716 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input284
timestamp 1623939100
transform 1 0 76912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input285
timestamp 1623939100
transform 1 0 77556 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_823
timestamp 1623939100
transform 1 0 76820 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_827
timestamp 1623939100
transform 1 0 77188 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_834
timestamp 1623939100
transform 1 0 77832 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_846
timestamp 1623939100
transform 1 0 78936 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_854
timestamp 1623939100
transform 1 0 79672 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1623939100
transform 1 0 79764 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_856
timestamp 1623939100
transform 1 0 79856 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_868
timestamp 1623939100
transform 1 0 80960 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 82248 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_201
timestamp 1623939100
transform 1 0 82064 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_889
timestamp 1623939100
transform 1 0 82892 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1623939100
transform 1 0 85008 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_901
timestamp 1623939100
transform 1 0 83996 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_909
timestamp 1623939100
transform 1 0 84732 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_913
timestamp 1623939100
transform 1 0 85100 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _706_
timestamp 1623939100
transform -1 0 87676 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1623939100
transform -1 0 85928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_919
timestamp 1623939100
transform 1 0 85652 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input175
timestamp 1623939100
transform 1 0 88044 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input177
timestamp 1623939100
transform 1 0 88688 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_941
timestamp 1623939100
transform 1 0 87676 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_948
timestamp 1623939100
transform 1 0 88320 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_955
timestamp 1623939100
transform 1 0 88964 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _497_
timestamp 1623939100
transform 1 0 90712 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1623939100
transform 1 0 90252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1623939100
transform 1 0 90528 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1623939100
transform 1 0 90344 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1623939100
transform 1 0 90068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input184
timestamp 1623939100
transform 1 0 92920 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1623939100
transform 1 0 92184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1623939100
transform 1 0 92368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1623939100
transform 1 0 92552 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1623939100
transform 1 0 92736 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input191
timestamp 1623939100
transform 1 0 94852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input197
timestamp 1623939100
transform 1 0 94208 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1001
timestamp 1623939100
transform 1 0 93196 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1009
timestamp 1623939100
transform 1 0 93932 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1015
timestamp 1623939100
transform 1 0 94484 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1623939100
transform 1 0 95496 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input190
timestamp 1623939100
transform 1 0 95956 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1022
timestamp 1623939100
transform 1 0 95128 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1027
timestamp 1623939100
transform 1 0 95588 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1034
timestamp 1623939100
transform 1 0 96232 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1623939100
transform -1 0 98808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1623939100
transform 1 0 97796 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1623939100
transform 1 0 97152 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1042
timestamp 1623939100
transform 1 0 96968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1047
timestamp 1623939100
transform 1 0 97428 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1054
timestamp 1623939100
transform 1 0 98072 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1058
timestamp 1623939100
transform 1 0 98440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1623939100
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1623939100
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input362
timestamp 1623939100
transform 1 0 2392 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1623939100
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_11
timestamp 1623939100
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1623939100
transform 1 0 2668 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1623939100
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1623939100
transform 1 0 2484 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp 1623939100
transform 1 0 3588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_23
timestamp 1623939100
transform 1 0 3220 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_30
timestamp 1623939100
transform 1 0 3864 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_28
timestamp 1623939100
transform 1 0 3680 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1623939100
transform 1 0 3312 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input364
timestamp 1623939100
transform 1 0 3312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input363
timestamp 1623939100
transform 1 0 3036 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1623939100
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_37
timestamp 1623939100
transform 1 0 4508 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input365
timestamp 1623939100
transform 1 0 4324 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _603_
timestamp 1623939100
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _575_
timestamp 1623939100
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1623939100
transform 1 0 4600 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1623939100
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1623939100
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_56
timestamp 1623939100
transform 1 0 6256 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1623939100
transform 1 0 5704 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_56
timestamp 1623939100
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1623939100
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _465_
timestamp 1623939100
transform 1 0 7636 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input327
timestamp 1623939100
transform 1 0 6992 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_191
timestamp 1623939100
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_202
timestamp 1623939100
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_67
timestamp 1623939100
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_82
timestamp 1623939100
transform 1 0 8648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1623939100
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1623939100
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1623939100
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1623939100
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1623939100
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1623939100
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1623939100
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1623939100
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1623939100
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1623939100
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1623939100
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1623939100
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_135
timestamp 1623939100
transform 1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1623939100
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1623939100
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_139
timestamp 1623939100
transform 1 0 13892 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 15088 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_194
timestamp 1623939100
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_156
timestamp 1623939100
transform 1 0 15456 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_147
timestamp 1623939100
transform 1 0 14628 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_161
timestamp 1623939100
transform 1 0 15916 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1623939100
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_168
timestamp 1623939100
transform 1 0 16560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_180
timestamp 1623939100
transform 1 0 17664 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1623939100
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1623939100
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1623939100
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1623939100
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_192
timestamp 1623939100
transform 1 0 18768 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1623939100
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1623939100
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1623939100
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform -1 0 21436 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1623939100
transform 1 0 22080 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_176
timestamp 1623939100
transform -1 0 20608 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_213
timestamp 1623939100
transform 1 0 20700 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_225
timestamp 1623939100
transform 1 0 21804 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_221
timestamp 1623939100
transform 1 0 21436 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_227
timestamp 1623939100
transform 1 0 21988 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_229
timestamp 1623939100
transform 1 0 22172 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_237
timestamp 1623939100
transform 1 0 22908 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_249
timestamp 1623939100
transform 1 0 24012 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_241
timestamp 1623939100
transform 1 0 23276 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1623939100
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_258
timestamp 1623939100
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_270
timestamp 1623939100
transform 1 0 25944 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_253
timestamp 1623939100
transform 1 0 24380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_265
timestamp 1623939100
transform 1 0 25484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _774_
timestamp 1623939100
transform 1 0 26220 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1623939100
transform 1 0 27324 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_277
timestamp 1623939100
transform 1 0 26588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_286
timestamp 1623939100
transform 1 0 27416 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_292
timestamp 1623939100
transform 1 0 27968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_304
timestamp 1623939100
transform 1 0 29072 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_312
timestamp 1623939100
transform 1 0 29808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_298
timestamp 1623939100
transform 1 0 28520 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_310
timestamp 1623939100
transform 1 0 29624 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1623939100
transform 1 0 29992 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_315
timestamp 1623939100
transform 1 0 30084 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_327
timestamp 1623939100
transform 1 0 31188 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_322
timestamp 1623939100
transform 1 0 30728 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _487_
timestamp 1623939100
transform 1 0 33028 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1623939100
transform 1 0 32568 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_339
timestamp 1623939100
transform 1 0 32292 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_351
timestamp 1623939100
transform 1 0 33396 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_334
timestamp 1623939100
transform 1 0 31832 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_343
timestamp 1623939100
transform 1 0 32660 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _622_
timestamp 1623939100
transform 1 0 34224 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1623939100
transform 1 0 35236 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_363
timestamp 1623939100
transform 1 0 34500 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_372
timestamp 1623939100
transform 1 0 35328 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_356
timestamp 1623939100
transform 1 0 33856 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_363
timestamp 1623939100
transform 1 0 34500 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_375
timestamp 1623939100
transform 1 0 35604 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_384
timestamp 1623939100
transform 1 0 36432 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_387
timestamp 1623939100
transform 1 0 36708 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1623939100
transform 1 0 37812 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_396
timestamp 1623939100
transform 1 0 37536 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_408
timestamp 1623939100
transform 1 0 38640 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_400
timestamp 1623939100
transform 1 0 37904 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_412
timestamp 1623939100
transform 1 0 39008 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1623939100
transform 1 0 40480 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_420
timestamp 1623939100
transform 1 0 39744 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_429
timestamp 1623939100
transform 1 0 40572 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_424
timestamp 1623939100
transform 1 0 40112 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_436
timestamp 1623939100
transform 1 0 41216 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1623939100
transform 1 0 43056 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_441
timestamp 1623939100
transform 1 0 41676 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_453
timestamp 1623939100
transform 1 0 42780 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_448
timestamp 1623939100
transform 1 0 42320 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_457
timestamp 1623939100
transform 1 0 43148 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_465
timestamp 1623939100
transform 1 0 43884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_477
timestamp 1623939100
transform 1 0 44988 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_469
timestamp 1623939100
transform 1 0 44252 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1623939100
transform 1 0 45724 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_486
timestamp 1623939100
transform 1 0 45816 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_498
timestamp 1623939100
transform 1 0 46920 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_481
timestamp 1623939100
transform 1 0 45356 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_493
timestamp 1623939100
transform 1 0 46460 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1623939100
transform 1 0 48300 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_510
timestamp 1623939100
transform 1 0 48024 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1623939100
transform 1 0 47564 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_514
timestamp 1623939100
transform 1 0 48392 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_522
timestamp 1623939100
transform 1 0 49128 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_534
timestamp 1623939100
transform 1 0 50232 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_526
timestamp 1623939100
transform 1 0 49496 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_538
timestamp 1623939100
transform 1 0 50600 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _731_
timestamp 1623939100
transform -1 0 53084 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1623939100
transform 1 0 50968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_58
timestamp 1623939100
transform -1 0 51336 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_543
timestamp 1623939100
transform 1 0 51060 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_555
timestamp 1623939100
transform 1 0 52164 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1623939100
transform 1 0 53544 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_567
timestamp 1623939100
transform 1 0 53268 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_579
timestamp 1623939100
transform 1 0 54372 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_565
timestamp 1623939100
transform 1 0 53084 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_569
timestamp 1623939100
transform 1 0 53452 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_571
timestamp 1623939100
transform 1 0 53636 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_583
timestamp 1623939100
transform 1 0 54740 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1623939100
transform 1 0 56212 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_591
timestamp 1623939100
transform 1 0 55476 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_600
timestamp 1623939100
transform 1 0 56304 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_595
timestamp 1623939100
transform 1 0 55844 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_612
timestamp 1623939100
transform 1 0 57408 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_624
timestamp 1623939100
transform 1 0 58512 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_607
timestamp 1623939100
transform 1 0 56948 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_619
timestamp 1623939100
transform 1 0 58052 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1623939100
transform 1 0 58788 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_636
timestamp 1623939100
transform 1 0 59616 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_628
timestamp 1623939100
transform 1 0 58880 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_640
timestamp 1623939100
transform 1 0 59984 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1623939100
transform 1 0 61456 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_648
timestamp 1623939100
transform 1 0 60720 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_657
timestamp 1623939100
transform 1 0 61548 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_652
timestamp 1623939100
transform 1 0 61088 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_664
timestamp 1623939100
transform 1 0 62192 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1623939100
transform 1 0 64032 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_669
timestamp 1623939100
transform 1 0 62652 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_681
timestamp 1623939100
transform 1 0 63756 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_676
timestamp 1623939100
transform 1 0 63296 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_685
timestamp 1623939100
transform 1 0 64124 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_693
timestamp 1623939100
transform 1 0 64860 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_705
timestamp 1623939100
transform 1 0 65964 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_697
timestamp 1623939100
transform 1 0 65228 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1623939100
transform 1 0 66700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_714
timestamp 1623939100
transform 1 0 66792 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_726
timestamp 1623939100
transform 1 0 67896 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_709
timestamp 1623939100
transform 1 0 66332 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_721
timestamp 1623939100
transform 1 0 67436 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1623939100
transform 1 0 69276 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_738
timestamp 1623939100
transform 1 0 69000 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_750
timestamp 1623939100
transform 1 0 70104 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_733
timestamp 1623939100
transform 1 0 68540 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_742
timestamp 1623939100
transform 1 0 69368 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1623939100
transform 1 0 71944 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_762
timestamp 1623939100
transform 1 0 71208 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_754
timestamp 1623939100
transform 1 0 70472 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_766
timestamp 1623939100
transform 1 0 71576 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_4  _424_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 73784 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_6_771
timestamp 1623939100
transform 1 0 72036 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_783
timestamp 1623939100
transform 1 0 73140 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_789
timestamp 1623939100
transform 1 0 73692 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_778
timestamp 1623939100
transform 1 0 72680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_790
timestamp 1623939100
transform 1 0 73784 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1623939100
transform 1 0 74520 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_795
timestamp 1623939100
transform 1 0 74244 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_807
timestamp 1623939100
transform 1 0 75348 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_799
timestamp 1623939100
transform 1 0 74612 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_811
timestamp 1623939100
transform 1 0 75716 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1623939100
transform 1 0 77188 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_819
timestamp 1623939100
transform 1 0 76452 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_828
timestamp 1623939100
transform 1 0 77280 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_823
timestamp 1623939100
transform 1 0 76820 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_840
timestamp 1623939100
transform 1 0 78384 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_852
timestamp 1623939100
transform 1 0 79488 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_835
timestamp 1623939100
transform 1 0 77924 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_847
timestamp 1623939100
transform 1 0 79028 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _551_
timestamp 1623939100
transform 1 0 81512 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1623939100
transform 1 0 79764 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_864
timestamp 1623939100
transform 1 0 80592 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_856
timestamp 1623939100
transform 1 0 79856 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_868
timestamp 1623939100
transform 1 0 80960 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1623939100
transform 1 0 82432 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_876
timestamp 1623939100
transform 1 0 81696 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_885
timestamp 1623939100
transform 1 0 82524 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_881
timestamp 1623939100
transform 1 0 82156 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_893
timestamp 1623939100
transform 1 0 83260 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1623939100
transform 1 0 85008 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_897
timestamp 1623939100
transform 1 0 83628 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_909
timestamp 1623939100
transform 1 0 84732 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_905
timestamp 1623939100
transform 1 0 84364 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_911
timestamp 1623939100
transform 1 0 84916 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_913
timestamp 1623939100
transform 1 0 85100 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_8  _437_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 85928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_921
timestamp 1623939100
transform 1 0 85836 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_933
timestamp 1623939100
transform 1 0 86940 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_921
timestamp 1623939100
transform 1 0 85836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_934
timestamp 1623939100
transform 1 0 87032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1623939100
transform 1 0 87676 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_942
timestamp 1623939100
transform 1 0 87768 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_954
timestamp 1623939100
transform 1 0 88872 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_946
timestamp 1623939100
transform 1 0 88136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_958
timestamp 1623939100
transform 1 0 89240 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1623939100
transform 1 0 90252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_966
timestamp 1623939100
transform 1 0 89976 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_978
timestamp 1623939100
transform 1 0 91080 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_966
timestamp 1623939100
transform 1 0 89976 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_970
timestamp 1623939100
transform 1 0 90344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1623939100
transform 1 0 92920 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_990
timestamp 1623939100
transform 1 0 92184 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_999
timestamp 1623939100
transform 1 0 93012 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_982
timestamp 1623939100
transform 1 0 91448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_994
timestamp 1623939100
transform 1 0 92552 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_197
timestamp 1623939100
transform 1 0 95036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1011
timestamp 1623939100
transform 1 0 94116 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_1019
timestamp 1623939100
transform 1 0 94852 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1006
timestamp 1623939100
transform 1 0 93656 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1018
timestamp 1623939100
transform 1 0 94760 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1027
timestamp 1623939100
transform 1 0 95588 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1623939100
transform 1 0 95496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _494_
timestamp 1623939100
transform 1 0 95220 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1037
timestamp 1623939100
transform 1 0 96508 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1031
timestamp 1623939100
transform 1 0 95956 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_1039
timestamp 1623939100
transform 1 0 96692 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1032
timestamp 1623939100
transform 1 0 96048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_217
timestamp 1623939100
transform -1 0 96232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input192
timestamp 1623939100
transform 1 0 96416 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _557_
timestamp 1623939100
transform -1 0 96508 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1041
timestamp 1623939100
transform 1 0 96876 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1045
timestamp 1623939100
transform 1 0 97244 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1047
timestamp 1623939100
transform 1 0 97428 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input193
timestamp 1623939100
transform 1 0 96968 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1623939100
transform 1 0 97520 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1052
timestamp 1623939100
transform 1 0 97888 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1051
timestamp 1623939100
transform 1 0 97796 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input194
timestamp 1623939100
transform 1 0 97612 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1623939100
transform 1 0 98164 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1058
timestamp 1623939100
transform 1 0 98440 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_1056
timestamp 1623939100
transform 1 0 98256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1623939100
transform -1 0 98808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1623939100
transform -1 0 98808 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1623939100
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1623939100
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_15
timestamp 1623939100
transform 1 0 2484 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_4  _461_
timestamp 1623939100
transform -1 0 5704 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1623939100
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_60
timestamp 1623939100
transform -1 0 4232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_62
timestamp 1623939100
transform -1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_65
timestamp 1623939100
transform -1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_67
timestamp 1623939100
transform -1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1623939100
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_61
timestamp 1623939100
transform -1 0 5888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_63
timestamp 1623939100
transform -1 0 6072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_64
timestamp 1623939100
transform -1 0 6256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_66
timestamp 1623939100
transform -1 0 6440 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_192
timestamp 1623939100
transform -1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_60
timestamp 1623939100
transform 1 0 6624 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_72
timestamp 1623939100
transform 1 0 7728 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1623939100
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1623939100
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1623939100
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1623939100
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1623939100
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1623939100
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1623939100
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1623939100
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1623939100
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_156
timestamp 1623939100
transform 1 0 15456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_168
timestamp 1623939100
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_180
timestamp 1623939100
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1623939100
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_192
timestamp 1623939100
transform 1 0 18768 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1623939100
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_213
timestamp 1623939100
transform 1 0 20700 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_225
timestamp 1623939100
transform 1 0 21804 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_237
timestamp 1623939100
transform 1 0 22908 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_249
timestamp 1623939100
transform 1 0 24012 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1623939100
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_258
timestamp 1623939100
transform 1 0 24840 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_270
timestamp 1623939100
transform 1 0 25944 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_282
timestamp 1623939100
transform 1 0 27048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_294
timestamp 1623939100
transform 1 0 28152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_306
timestamp 1623939100
transform 1 0 29256 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1623939100
transform 1 0 29992 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_315
timestamp 1623939100
transform 1 0 30084 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_327
timestamp 1623939100
transform 1 0 31188 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_339
timestamp 1623939100
transform 1 0 32292 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_351
timestamp 1623939100
transform 1 0 33396 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1623939100
transform 1 0 35236 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_363
timestamp 1623939100
transform 1 0 34500 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_372
timestamp 1623939100
transform 1 0 35328 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_384
timestamp 1623939100
transform 1 0 36432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_396
timestamp 1623939100
transform 1 0 37536 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_408
timestamp 1623939100
transform 1 0 38640 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1623939100
transform 1 0 40480 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_420
timestamp 1623939100
transform 1 0 39744 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_429
timestamp 1623939100
transform 1 0 40572 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _654_
timestamp 1623939100
transform 1 0 43148 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_441
timestamp 1623939100
transform 1 0 41676 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_453
timestamp 1623939100
transform 1 0 42780 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_460
timestamp 1623939100
transform 1 0 43424 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_472
timestamp 1623939100
transform 1 0 44528 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1623939100
transform 1 0 45724 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_484
timestamp 1623939100
transform 1 0 45632 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_486
timestamp 1623939100
transform 1 0 45816 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_498
timestamp 1623939100
transform 1 0 46920 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_510
timestamp 1623939100
transform 1 0 48024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_522
timestamp 1623939100
transform 1 0 49128 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_534
timestamp 1623939100
transform 1 0 50232 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1623939100
transform 1 0 50968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_543
timestamp 1623939100
transform 1 0 51060 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_555
timestamp 1623939100
transform 1 0 52164 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_567
timestamp 1623939100
transform 1 0 53268 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_579
timestamp 1623939100
transform 1 0 54372 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1623939100
transform 1 0 56212 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_591
timestamp 1623939100
transform 1 0 55476 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_600
timestamp 1623939100
transform 1 0 56304 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_612
timestamp 1623939100
transform 1 0 57408 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_624
timestamp 1623939100
transform 1 0 58512 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_636
timestamp 1623939100
transform 1 0 59616 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _790_
timestamp 1623939100
transform 1 0 61916 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1623939100
transform 1 0 61456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_648
timestamp 1623939100
transform 1 0 60720 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_657
timestamp 1623939100
transform 1 0 61548 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_680
timestamp 1623939100
transform 1 0 63664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_692
timestamp 1623939100
transform 1 0 64768 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_704
timestamp 1623939100
transform 1 0 65872 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1623939100
transform 1 0 66700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_712
timestamp 1623939100
transform 1 0 66608 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_714
timestamp 1623939100
transform 1 0 66792 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_726
timestamp 1623939100
transform 1 0 67896 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_738
timestamp 1623939100
transform 1 0 69000 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_750
timestamp 1623939100
transform 1 0 70104 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1623939100
transform 1 0 71944 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_762
timestamp 1623939100
transform 1 0 71208 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _550_
timestamp 1623939100
transform 1 0 72404 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_771
timestamp 1623939100
transform 1 0 72036 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_781
timestamp 1623939100
transform 1 0 72956 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_793
timestamp 1623939100
transform 1 0 74060 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_805
timestamp 1623939100
transform 1 0 75164 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1623939100
transform 1 0 77188 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_817
timestamp 1623939100
transform 1 0 76268 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_825
timestamp 1623939100
transform 1 0 77004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_828
timestamp 1623939100
transform 1 0 77280 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_840
timestamp 1623939100
transform 1 0 78384 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_852
timestamp 1623939100
transform 1 0 79488 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_864
timestamp 1623939100
transform 1 0 80592 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1623939100
transform 1 0 82432 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_876
timestamp 1623939100
transform 1 0 81696 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_885
timestamp 1623939100
transform 1 0 82524 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_897
timestamp 1623939100
transform 1 0 83628 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_909
timestamp 1623939100
transform 1 0 84732 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_921
timestamp 1623939100
transform 1 0 85836 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_933
timestamp 1623939100
transform 1 0 86940 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1623939100
transform 1 0 87676 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_942
timestamp 1623939100
transform 1 0 87768 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_954
timestamp 1623939100
transform 1 0 88872 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_966
timestamp 1623939100
transform 1 0 89976 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_978
timestamp 1623939100
transform 1 0 91080 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1623939100
transform 1 0 92920 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_990
timestamp 1623939100
transform 1 0 92184 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_999
timestamp 1623939100
transform 1 0 93012 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1011
timestamp 1623939100
transform 1 0 94116 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1023
timestamp 1623939100
transform 1 0 95220 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1035
timestamp 1623939100
transform 1 0 96324 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1623939100
transform -1 0 98808 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1623939100
transform 1 0 98164 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input195
timestamp 1623939100
transform 1 0 97520 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1047
timestamp 1623939100
transform 1 0 97428 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1051
timestamp 1623939100
transform 1 0 97796 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_1056
timestamp 1623939100
transform 1 0 98256 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1623939100
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1623939100
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1623939100
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1623939100
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1623939100
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1623939100
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1623939100
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1623939100
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1623939100
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1623939100
transform 1 0 8648 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_4  _490_
timestamp 1623939100
transform 1 0 9108 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_86
timestamp 1623939100
transform 1 0 9016 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1623939100
transform 1 0 10580 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _564_
timestamp 1623939100
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1623939100
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_240
timestamp 1623939100
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_111
timestamp 1623939100
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_115
timestamp 1623939100
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_122
timestamp 1623939100
transform 1 0 12328 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_134
timestamp 1623939100
transform 1 0 13432 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_146
timestamp 1623939100
transform 1 0 14536 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_158
timestamp 1623939100
transform 1 0 15640 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1623939100
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_170
timestamp 1623939100
transform 1 0 16744 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1623939100
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1623939100
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1623939100
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1623939100
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1623939100
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_220
timestamp 1623939100
transform 1 0 21344 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_229
timestamp 1623939100
transform 1 0 22172 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_241
timestamp 1623939100
transform 1 0 23276 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _472_
timestamp 1623939100
transform -1 0 25852 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_164
timestamp 1623939100
transform -1 0 25024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_200
timestamp 1623939100
transform -1 0 26036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_253
timestamp 1623939100
transform 1 0 24380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_257
timestamp 1623939100
transform 1 0 24748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1623939100
transform 1 0 27324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_271
timestamp 1623939100
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1623939100
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_286
timestamp 1623939100
transform 1 0 27416 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_298
timestamp 1623939100
transform 1 0 28520 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_310
timestamp 1623939100
transform 1 0 29624 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_322
timestamp 1623939100
transform 1 0 30728 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1623939100
transform 1 0 32568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_334
timestamp 1623939100
transform 1 0 31832 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_343
timestamp 1623939100
transform 1 0 32660 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_355
timestamp 1623939100
transform 1 0 33764 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1623939100
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1623939100
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_391
timestamp 1623939100
transform 1 0 37076 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _659_
timestamp 1623939100
transform 1 0 38364 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1623939100
transform 1 0 37812 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_400
timestamp 1623939100
transform 1 0 37904 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_404
timestamp 1623939100
transform 1 0 38272 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_408
timestamp 1623939100
transform 1 0 38640 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_420
timestamp 1623939100
transform 1 0 39744 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_432
timestamp 1623939100
transform 1 0 40848 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1623939100
transform 1 0 43056 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_444
timestamp 1623939100
transform 1 0 41952 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_457
timestamp 1623939100
transform 1 0 43148 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_469
timestamp 1623939100
transform 1 0 44252 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_481
timestamp 1623939100
transform 1 0 45356 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_493
timestamp 1623939100
transform 1 0 46460 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1623939100
transform 1 0 48300 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1623939100
transform 1 0 47564 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_514
timestamp 1623939100
transform 1 0 48392 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_4  _327_
timestamp 1623939100
transform 1 0 49220 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_522
timestamp 1623939100
transform 1 0 49128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_539
timestamp 1623939100
transform 1 0 50692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_551
timestamp 1623939100
transform 1 0 51796 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1623939100
transform 1 0 53544 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_563
timestamp 1623939100
transform 1 0 52900 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_569
timestamp 1623939100
transform 1 0 53452 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_571
timestamp 1623939100
transform 1 0 53636 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_583
timestamp 1623939100
transform 1 0 54740 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_595
timestamp 1623939100
transform 1 0 55844 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_607
timestamp 1623939100
transform 1 0 56948 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_619
timestamp 1623939100
transform 1 0 58052 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1623939100
transform 1 0 58788 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_628
timestamp 1623939100
transform 1 0 58880 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_640
timestamp 1623939100
transform 1 0 59984 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_652
timestamp 1623939100
transform 1 0 61088 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_664
timestamp 1623939100
transform 1 0 62192 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1623939100
transform 1 0 64032 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_676
timestamp 1623939100
transform 1 0 63296 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_685
timestamp 1623939100
transform 1 0 64124 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_697
timestamp 1623939100
transform 1 0 65228 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_709
timestamp 1623939100
transform 1 0 66332 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_721
timestamp 1623939100
transform 1 0 67436 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _559_
timestamp 1623939100
transform 1 0 69736 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1623939100
transform 1 0 69276 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_219
timestamp 1623939100
transform 1 0 69552 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_733
timestamp 1623939100
transform 1 0 68540 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_742
timestamp 1623939100
transform 1 0 69368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_749
timestamp 1623939100
transform 1 0 70012 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_761
timestamp 1623939100
transform 1 0 71116 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_773
timestamp 1623939100
transform 1 0 72220 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_785
timestamp 1623939100
transform 1 0 73324 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1623939100
transform 1 0 74520 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_797
timestamp 1623939100
transform 1 0 74428 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_799
timestamp 1623939100
transform 1 0 74612 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_811
timestamp 1623939100
transform 1 0 75716 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_823
timestamp 1623939100
transform 1 0 76820 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_835
timestamp 1623939100
transform 1 0 77924 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_847
timestamp 1623939100
transform 1 0 79028 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1623939100
transform 1 0 79764 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_856
timestamp 1623939100
transform 1 0 79856 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_868
timestamp 1623939100
transform 1 0 80960 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_880
timestamp 1623939100
transform 1 0 82064 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_892
timestamp 1623939100
transform 1 0 83168 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1623939100
transform 1 0 85008 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_904
timestamp 1623939100
transform 1 0 84272 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_913
timestamp 1623939100
transform 1 0 85100 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _317_
timestamp 1623939100
transform 1 0 86848 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_925
timestamp 1623939100
transform 1 0 86204 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_931
timestamp 1623939100
transform 1 0 86756 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_938
timestamp 1623939100
transform 1 0 87400 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_950
timestamp 1623939100
transform 1 0 88504 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1623939100
transform 1 0 90252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_962
timestamp 1623939100
transform 1 0 89608 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_968
timestamp 1623939100
transform 1 0 90160 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_970
timestamp 1623939100
transform 1 0 90344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_982
timestamp 1623939100
transform 1 0 91448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_994
timestamp 1623939100
transform 1 0 92552 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1006
timestamp 1623939100
transform 1 0 93656 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1018
timestamp 1623939100
transform 1 0 94760 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1623939100
transform 1 0 95496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1027
timestamp 1623939100
transform 1 0 95588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1039
timestamp 1623939100
transform 1 0 96692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1623939100
transform -1 0 98808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input196
timestamp 1623939100
transform 1 0 97888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1051
timestamp 1623939100
transform 1 0 97796 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1055
timestamp 1623939100
transform 1 0 98164 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_4  _488_
timestamp 1623939100
transform 1 0 1380 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1623939100
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1623939100
transform 1 0 2852 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1623939100
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1623939100
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1623939100
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1623939100
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1623939100
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1623939100
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1623939100
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _393_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 9752 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1623939100
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_246
timestamp 1623939100
transform 1 0 9568 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1623939100
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1623939100
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_108
timestamp 1623939100
transform 1 0 11040 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_120
timestamp 1623939100
transform 1 0 12144 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1623939100
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_132
timestamp 1623939100
transform 1 0 13248 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_140
timestamp 1623939100
transform 1 0 13984 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1623939100
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_156
timestamp 1623939100
transform 1 0 15456 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_168
timestamp 1623939100
transform 1 0 16560 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1623939100
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1623939100
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_192
timestamp 1623939100
transform 1 0 18768 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1623939100
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_213
timestamp 1623939100
transform 1 0 20700 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_225
timestamp 1623939100
transform 1 0 21804 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_237
timestamp 1623939100
transform 1 0 22908 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_249
timestamp 1623939100
transform 1 0 24012 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1623939100
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_258
timestamp 1623939100
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_270
timestamp 1623939100
transform 1 0 25944 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_282
timestamp 1623939100
transform 1 0 27048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_294
timestamp 1623939100
transform 1 0 28152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_306
timestamp 1623939100
transform 1 0 29256 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1623939100
transform 1 0 29992 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_315
timestamp 1623939100
transform 1 0 30084 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_327
timestamp 1623939100
transform 1 0 31188 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _703_
timestamp 1623939100
transform 1 0 31924 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_10_354
timestamp 1623939100
transform 1 0 33672 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1623939100
transform 1 0 35236 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_366
timestamp 1623939100
transform 1 0 34776 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_370
timestamp 1623939100
transform 1 0 35144 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_372
timestamp 1623939100
transform 1 0 35328 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _519_
timestamp 1623939100
transform 1 0 37260 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_384
timestamp 1623939100
transform 1 0 36432 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_392
timestamp 1623939100
transform 1 0 37168 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _420_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 39100 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_409
timestamp 1623939100
transform 1 0 38732 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1623939100
transform 1 0 40480 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_421
timestamp 1623939100
transform 1 0 39836 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_427
timestamp 1623939100
transform 1 0 40388 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_429
timestamp 1623939100
transform 1 0 40572 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_441
timestamp 1623939100
transform 1 0 41676 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_453
timestamp 1623939100
transform 1 0 42780 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_465
timestamp 1623939100
transform 1 0 43884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_477
timestamp 1623939100
transform 1 0 44988 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1623939100
transform 1 0 45724 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_486
timestamp 1623939100
transform 1 0 45816 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_498
timestamp 1623939100
transform 1 0 46920 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_510
timestamp 1623939100
transform 1 0 48024 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_522
timestamp 1623939100
transform 1 0 49128 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_534
timestamp 1623939100
transform 1 0 50232 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1623939100
transform 1 0 50968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_543
timestamp 1623939100
transform 1 0 51060 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_555
timestamp 1623939100
transform 1 0 52164 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_567
timestamp 1623939100
transform 1 0 53268 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_579
timestamp 1623939100
transform 1 0 54372 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1623939100
transform 1 0 56212 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_591
timestamp 1623939100
transform 1 0 55476 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_600
timestamp 1623939100
transform 1 0 56304 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_612
timestamp 1623939100
transform 1 0 57408 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_624
timestamp 1623939100
transform 1 0 58512 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_636
timestamp 1623939100
transform 1 0 59616 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1623939100
transform 1 0 61456 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_648
timestamp 1623939100
transform 1 0 60720 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_657
timestamp 1623939100
transform 1 0 61548 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_669
timestamp 1623939100
transform 1 0 62652 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_681
timestamp 1623939100
transform 1 0 63756 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_693
timestamp 1623939100
transform 1 0 64860 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_705
timestamp 1623939100
transform 1 0 65964 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1623939100
transform 1 0 66700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_714
timestamp 1623939100
transform 1 0 66792 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_726
timestamp 1623939100
transform 1 0 67896 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_738
timestamp 1623939100
transform 1 0 69000 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_750
timestamp 1623939100
transform 1 0 70104 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1623939100
transform 1 0 71944 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_762
timestamp 1623939100
transform 1 0 71208 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_771
timestamp 1623939100
transform 1 0 72036 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_783
timestamp 1623939100
transform 1 0 73140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_795
timestamp 1623939100
transform 1 0 74244 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_807
timestamp 1623939100
transform 1 0 75348 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1623939100
transform 1 0 77188 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_819
timestamp 1623939100
transform 1 0 76452 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_828
timestamp 1623939100
transform 1 0 77280 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_840
timestamp 1623939100
transform 1 0 78384 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_852
timestamp 1623939100
transform 1 0 79488 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_864
timestamp 1623939100
transform 1 0 80592 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1623939100
transform 1 0 82432 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_876
timestamp 1623939100
transform 1 0 81696 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_885
timestamp 1623939100
transform 1 0 82524 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_897
timestamp 1623939100
transform 1 0 83628 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_909
timestamp 1623939100
transform 1 0 84732 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_921
timestamp 1623939100
transform 1 0 85836 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_933
timestamp 1623939100
transform 1 0 86940 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1623939100
transform 1 0 87676 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_942
timestamp 1623939100
transform 1 0 87768 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_954
timestamp 1623939100
transform 1 0 88872 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_966
timestamp 1623939100
transform 1 0 89976 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_978
timestamp 1623939100
transform 1 0 91080 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1623939100
transform 1 0 92920 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_990
timestamp 1623939100
transform 1 0 92184 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_999
timestamp 1623939100
transform 1 0 93012 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _301_
timestamp 1623939100
transform 1 0 94392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1011
timestamp 1623939100
transform 1 0 94116 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1023
timestamp 1623939100
transform 1 0 95220 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1035
timestamp 1623939100
transform 1 0 96324 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1623939100
transform -1 0 98808 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1623939100
transform 1 0 98164 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1047
timestamp 1623939100
transform 1 0 97428 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_1056
timestamp 1623939100
transform 1 0 98256 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1623939100
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1623939100
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1623939100
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1623939100
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1623939100
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1623939100
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1623939100
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1623939100
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1623939100
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_82
timestamp 1623939100
transform 1 0 8648 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_94
timestamp 1623939100
transform 1 0 9752 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1623939100
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_106
timestamp 1623939100
transform 1 0 10856 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1623939100
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1623939100
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1623939100
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_151
timestamp 1623939100
transform 1 0 14996 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_163
timestamp 1623939100
transform 1 0 16100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1623939100
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1623939100
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1623939100
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _373_
timestamp 1623939100
transform 1 0 19780 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_196
timestamp 1623939100
transform 1 0 19136 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_202
timestamp 1623939100
transform 1 0 19688 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1623939100
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_212
timestamp 1623939100
transform 1 0 20608 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_224
timestamp 1623939100
transform 1 0 21712 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_229
timestamp 1623939100
transform 1 0 22172 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _432_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 23000 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_237
timestamp 1623939100
transform 1 0 22908 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_246
timestamp 1623939100
transform 1 0 23736 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_258
timestamp 1623939100
transform 1 0 24840 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_270
timestamp 1623939100
transform 1 0 25944 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1623939100
transform 1 0 27324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_282
timestamp 1623939100
transform 1 0 27048 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_286
timestamp 1623939100
transform 1 0 27416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_298
timestamp 1623939100
transform 1 0 28520 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_310
timestamp 1623939100
transform 1 0 29624 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_322
timestamp 1623939100
transform 1 0 30728 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _427_
timestamp 1623939100
transform 1 0 33672 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1623939100
transform 1 0 32568 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_334
timestamp 1623939100
transform 1 0 31832 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_343
timestamp 1623939100
transform 1 0 32660 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_351
timestamp 1623939100
transform 1 0 33396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _321_
timestamp 1623939100
transform 1 0 35144 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_11_366
timestamp 1623939100
transform 1 0 34776 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_377
timestamp 1623939100
transform 1 0 35788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_389
timestamp 1623939100
transform 1 0 36892 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _434_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 38824 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1623939100
transform 1 0 37812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_397
timestamp 1623939100
transform 1 0 37628 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_400
timestamp 1623939100
transform 1 0 37904 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_408
timestamp 1623939100
transform 1 0 38640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_419
timestamp 1623939100
transform 1 0 39652 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_431
timestamp 1623939100
transform 1 0 40756 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1623939100
transform 1 0 43056 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_443
timestamp 1623939100
transform 1 0 41860 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_455
timestamp 1623939100
transform 1 0 42964 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_457
timestamp 1623939100
transform 1 0 43148 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_469
timestamp 1623939100
transform 1 0 44252 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_481
timestamp 1623939100
transform 1 0 45356 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_493
timestamp 1623939100
transform 1 0 46460 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1623939100
transform 1 0 48300 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1623939100
transform 1 0 47564 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_514
timestamp 1623939100
transform 1 0 48392 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_520
timestamp 1623939100
transform 1 0 48944 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_2  _401_
timestamp 1623939100
transform 1 0 50416 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__conb_1  _612_
timestamp 1623939100
transform 1 0 49036 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_524
timestamp 1623939100
transform 1 0 49312 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_543
timestamp 1623939100
transform 1 0 51060 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_555
timestamp 1623939100
transform 1 0 52164 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _604_
timestamp 1623939100
transform 1 0 54096 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1623939100
transform 1 0 53544 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_567
timestamp 1623939100
transform 1 0 53268 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_571
timestamp 1623939100
transform 1 0 53636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_575
timestamp 1623939100
transform 1 0 54004 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_579
timestamp 1623939100
transform 1 0 54372 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _632_
timestamp 1623939100
transform 1 0 56396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_591
timestamp 1623939100
transform 1 0 55476 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_599
timestamp 1623939100
transform 1 0 56212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_604
timestamp 1623939100
transform 1 0 56672 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_616
timestamp 1623939100
transform 1 0 57776 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_624
timestamp 1623939100
transform 1 0 58512 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1623939100
transform 1 0 58788 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_628
timestamp 1623939100
transform 1 0 58880 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_640
timestamp 1623939100
transform 1 0 59984 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _496_
timestamp 1623939100
transform 1 0 61180 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_652
timestamp 1623939100
transform 1 0 61088 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_662
timestamp 1623939100
transform 1 0 62008 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1623939100
transform 1 0 64032 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_674
timestamp 1623939100
transform 1 0 63112 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_682
timestamp 1623939100
transform 1 0 63848 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_685
timestamp 1623939100
transform 1 0 64124 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _336_
timestamp 1623939100
transform 1 0 65872 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_697
timestamp 1623939100
transform 1 0 65228 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_703
timestamp 1623939100
transform 1 0 65780 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _374_
timestamp 1623939100
transform 1 0 67344 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_713
timestamp 1623939100
transform 1 0 66700 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_719
timestamp 1623939100
transform 1 0 67252 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_729
timestamp 1623939100
transform 1 0 68172 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1623939100
transform 1 0 69276 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_742
timestamp 1623939100
transform 1 0 69368 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_754
timestamp 1623939100
transform 1 0 70472 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_766
timestamp 1623939100
transform 1 0 71576 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_778
timestamp 1623939100
transform 1 0 72680 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_790
timestamp 1623939100
transform 1 0 73784 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1623939100
transform 1 0 74520 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_799
timestamp 1623939100
transform 1 0 74612 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_811
timestamp 1623939100
transform 1 0 75716 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_823
timestamp 1623939100
transform 1 0 76820 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_835
timestamp 1623939100
transform 1 0 77924 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_847
timestamp 1623939100
transform 1 0 79028 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1623939100
transform 1 0 79764 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_856
timestamp 1623939100
transform 1 0 79856 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_868
timestamp 1623939100
transform 1 0 80960 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_880
timestamp 1623939100
transform 1 0 82064 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_892
timestamp 1623939100
transform 1 0 83168 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1623939100
transform 1 0 85008 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_904
timestamp 1623939100
transform 1 0 84272 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_913
timestamp 1623939100
transform 1 0 85100 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_925
timestamp 1623939100
transform 1 0 86204 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_937
timestamp 1623939100
transform 1 0 87308 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_949
timestamp 1623939100
transform 1 0 88412 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1623939100
transform 1 0 90252 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_961
timestamp 1623939100
transform 1 0 89516 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_970
timestamp 1623939100
transform 1 0 90344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_982
timestamp 1623939100
transform 1 0 91448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_994
timestamp 1623939100
transform 1 0 92552 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _538_
timestamp 1623939100
transform 1 0 94300 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_378
timestamp 1623939100
transform 1 0 94116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1006
timestamp 1623939100
transform 1 0 93656 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1010
timestamp 1623939100
transform 1 0 94024 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1623939100
transform 1 0 95496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_385
timestamp 1623939100
transform 1 0 95128 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1024
timestamp 1623939100
transform 1 0 95312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1027
timestamp 1623939100
transform 1 0 95588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1039
timestamp 1623939100
transform 1 0 96692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1623939100
transform -1 0 98808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1051
timestamp 1623939100
transform 1 0 97796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1623939100
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1623939100
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1623939100
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _532_
timestamp 1623939100
transform 1 0 4692 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1623939100
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1623939100
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_30
timestamp 1623939100
transform 1 0 3864 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_38
timestamp 1623939100
transform 1 0 4600 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_55
timestamp 1623939100
transform 1 0 6164 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_67
timestamp 1623939100
transform 1 0 7268 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_79
timestamp 1623939100
transform 1 0 8372 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1623939100
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1623939100
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_87
timestamp 1623939100
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_99
timestamp 1623939100
transform 1 0 10212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _460_
timestamp 1623939100
transform 1 0 11592 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_162
timestamp 1623939100
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_204
timestamp 1623939100
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_111
timestamp 1623939100
transform 1 0 11316 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_125
timestamp 1623939100
transform 1 0 12604 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1623939100
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_137
timestamp 1623939100
transform 1 0 13708 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1623939100
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_2  _325_
timestamp 1623939100
transform 1 0 16192 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_156
timestamp 1623939100
transform 1 0 15456 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_171
timestamp 1623939100
transform 1 0 16836 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_183
timestamp 1623939100
transform 1 0 17940 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1623939100
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_195
timestamp 1623939100
transform 1 0 19044 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_199
timestamp 1623939100
transform 1 0 19412 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1623939100
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _776_
timestamp 1623939100
transform 1 0 20792 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1623939100
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1623939100
transform 1 0 22540 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_245
timestamp 1623939100
transform 1 0 23644 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1623939100
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_258
timestamp 1623939100
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_270
timestamp 1623939100
transform 1 0 25944 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_282
timestamp 1623939100
transform 1 0 27048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_294
timestamp 1623939100
transform 1 0 28152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_306
timestamp 1623939100
transform 1 0 29256 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1623939100
transform 1 0 29992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_315
timestamp 1623939100
transform 1 0 30084 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_327
timestamp 1623939100
transform 1 0 31188 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_339
timestamp 1623939100
transform 1 0 32292 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_351
timestamp 1623939100
transform 1 0 33396 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1623939100
transform 1 0 35236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_363
timestamp 1623939100
transform 1 0 34500 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_372
timestamp 1623939100
transform 1 0 35328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _383_
timestamp 1623939100
transform 1 0 36892 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_384
timestamp 1623939100
transform 1 0 36432 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_388
timestamp 1623939100
transform 1 0 36800 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _727_
timestamp 1623939100
transform 1 0 38088 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_12_398
timestamp 1623939100
transform 1 0 37720 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1623939100
transform 1 0 40480 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_421
timestamp 1623939100
transform 1 0 39836 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_427
timestamp 1623939100
transform 1 0 40388 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_429
timestamp 1623939100
transform 1 0 40572 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_441
timestamp 1623939100
transform 1 0 41676 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_453
timestamp 1623939100
transform 1 0 42780 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_465
timestamp 1623939100
transform 1 0 43884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_477
timestamp 1623939100
transform 1 0 44988 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1623939100
transform 1 0 45724 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_486
timestamp 1623939100
transform 1 0 45816 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_498
timestamp 1623939100
transform 1 0 46920 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_510
timestamp 1623939100
transform 1 0 48024 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_522
timestamp 1623939100
transform 1 0 49128 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_534
timestamp 1623939100
transform 1 0 50232 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1623939100
transform 1 0 50968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_543
timestamp 1623939100
transform 1 0 51060 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_555
timestamp 1623939100
transform 1 0 52164 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_567
timestamp 1623939100
transform 1 0 53268 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_579
timestamp 1623939100
transform 1 0 54372 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1623939100
transform 1 0 56212 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_591
timestamp 1623939100
transform 1 0 55476 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_600
timestamp 1623939100
transform 1 0 56304 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_612
timestamp 1623939100
transform 1 0 57408 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_624
timestamp 1623939100
transform 1 0 58512 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_636
timestamp 1623939100
transform 1 0 59616 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1623939100
transform 1 0 61456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_648
timestamp 1623939100
transform 1 0 60720 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_657
timestamp 1623939100
transform 1 0 61548 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _715_
timestamp 1623939100
transform 1 0 62744 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_12_669
timestamp 1623939100
transform 1 0 62652 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_689
timestamp 1623939100
transform 1 0 64492 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_701
timestamp 1623939100
transform 1 0 65596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1623939100
transform 1 0 66700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_714
timestamp 1623939100
transform 1 0 66792 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_726
timestamp 1623939100
transform 1 0 67896 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_738
timestamp 1623939100
transform 1 0 69000 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_750
timestamp 1623939100
transform 1 0 70104 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1623939100
transform 1 0 71944 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_762
timestamp 1623939100
transform 1 0 71208 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _283_
timestamp 1623939100
transform 1 0 73784 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_771
timestamp 1623939100
transform 1 0 72036 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_783
timestamp 1623939100
transform 1 0 73140 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_789
timestamp 1623939100
transform 1 0 73692 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_799
timestamp 1623939100
transform 1 0 74612 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_811
timestamp 1623939100
transform 1 0 75716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1623939100
transform 1 0 77188 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_823
timestamp 1623939100
transform 1 0 76820 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_828
timestamp 1623939100
transform 1 0 77280 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_840
timestamp 1623939100
transform 1 0 78384 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_852
timestamp 1623939100
transform 1 0 79488 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_864
timestamp 1623939100
transform 1 0 80592 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1623939100
transform 1 0 82432 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_876
timestamp 1623939100
transform 1 0 81696 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_885
timestamp 1623939100
transform 1 0 82524 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_897
timestamp 1623939100
transform 1 0 83628 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_909
timestamp 1623939100
transform 1 0 84732 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_921
timestamp 1623939100
transform 1 0 85836 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_933
timestamp 1623939100
transform 1 0 86940 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _318_
timestamp 1623939100
transform 1 0 88320 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1623939100
transform 1 0 87676 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_942
timestamp 1623939100
transform 1 0 87768 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_962
timestamp 1623939100
transform 1 0 89608 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_974
timestamp 1623939100
transform 1 0 90712 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1623939100
transform 1 0 92920 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_986
timestamp 1623939100
transform 1 0 91816 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_999
timestamp 1623939100
transform 1 0 93012 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _467_
timestamp 1623939100
transform 1 0 95036 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1011
timestamp 1623939100
transform 1 0 94116 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_1019
timestamp 1623939100
transform 1 0 94852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1030
timestamp 1623939100
transform 1 0 95864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1623939100
transform -1 0 98808 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1623939100
transform 1 0 98164 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1042
timestamp 1623939100
transform 1 0 96968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1054
timestamp 1623939100
transform 1 0 98072 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_1056
timestamp 1623939100
transform 1 0 98256 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1623939100
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1623939100
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1623939100
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_15
timestamp 1623939100
transform 1 0 2484 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1623939100
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1623939100
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _331_
timestamp 1623939100
transform 1 0 4232 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _396_
timestamp 1623939100
transform 1 0 3128 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1623939100
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_21
timestamp 1623939100
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_29
timestamp 1623939100
transform 1 0 3772 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_41
timestamp 1623939100
transform 1 0 4876 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1623939100
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_30
timestamp 1623939100
transform 1 0 3864 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _294_
timestamp 1623939100
transform 1 0 6440 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1623939100
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_53
timestamp 1623939100
transform 1 0 5980 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1623939100
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_43
timestamp 1623939100
transform 1 0 5060 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_55
timestamp 1623939100
transform 1 0 6164 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1623939100
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1623939100
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_70
timestamp 1623939100
transform 1 0 7544 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_82
timestamp 1623939100
transform 1 0 8648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _764_
timestamp 1623939100
transform -1 0 11224 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1623939100
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_115
timestamp 1623939100
transform -1 0 9476 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1623939100
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_87
timestamp 1623939100
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _364_
timestamp 1623939100
transform 1 0 12420 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1623939100
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_106
timestamp 1623939100
transform 1 0 10856 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_115
timestamp 1623939100
transform 1 0 11684 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_110
timestamp 1623939100
transform 1 0 11224 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_122
timestamp 1623939100
transform 1 0 12328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1623939100
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_130
timestamp 1623939100
transform 1 0 13064 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_142
timestamp 1623939100
transform 1 0 14168 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_134
timestamp 1623939100
transform 1 0 13432 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1623939100
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1623939100
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1623939100
transform 1 0 15272 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_166
timestamp 1623939100
transform 1 0 16376 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1623939100
transform 1 0 15456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1623939100
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_170
timestamp 1623939100
transform 1 0 16744 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1623939100
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_184
timestamp 1623939100
transform 1 0 18032 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_168
timestamp 1623939100
transform 1 0 16560 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1623939100
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _388_
timestamp 1623939100
transform -1 0 19780 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _628_
timestamp 1623939100
transform 1 0 20148 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1623939100
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_148
timestamp 1623939100
transform -1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_203
timestamp 1623939100
transform 1 0 19780 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_192
timestamp 1623939100
transform 1 0 18768 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1623939100
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1623939100
transform 1 0 22080 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_210
timestamp 1623939100
transform 1 0 20424 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_222
timestamp 1623939100
transform 1 0 21528 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_229
timestamp 1623939100
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_213
timestamp 1623939100
transform 1 0 20700 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_225
timestamp 1623939100
transform 1 0 21804 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_241
timestamp 1623939100
transform 1 0 23276 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_237
timestamp 1623939100
transform 1 0 22908 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_249
timestamp 1623939100
transform 1 0 24012 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _772_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 25852 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1623939100
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_253
timestamp 1623939100
transform 1 0 24380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_265
timestamp 1623939100
transform 1 0 25484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1623939100
transform 1 0 24840 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_266
timestamp 1623939100
transform 1 0 25576 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1623939100
transform 1 0 27324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_277
timestamp 1623939100
transform 1 0 26588 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_286
timestamp 1623939100
transform 1 0 27416 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_286
timestamp 1623939100
transform 1 0 27416 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__inv_4  _279_
timestamp 1623939100
transform 1 0 27968 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_13_298
timestamp 1623939100
transform 1 0 28520 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_310
timestamp 1623939100
transform 1 0 29624 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_297
timestamp 1623939100
transform 1 0 28428 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_309
timestamp 1623939100
transform 1 0 29532 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1623939100
transform 1 0 29992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_322
timestamp 1623939100
transform 1 0 30728 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_313
timestamp 1623939100
transform 1 0 29900 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_315
timestamp 1623939100
transform 1 0 30084 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_327
timestamp 1623939100
transform 1 0 31188 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1623939100
transform 1 0 32568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_334
timestamp 1623939100
transform 1 0 31832 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_343
timestamp 1623939100
transform 1 0 32660 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_339
timestamp 1623939100
transform 1 0 32292 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_351
timestamp 1623939100
transform 1 0 33396 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_4  _549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 35512 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1623939100
transform 1 0 35236 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_355
timestamp 1623939100
transform 1 0 33764 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_367
timestamp 1623939100
transform 1 0 34868 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_373
timestamp 1623939100
transform 1 0 35420 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_363
timestamp 1623939100
transform 1 0 34500 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_372
timestamp 1623939100
transform 1 0 35328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_391
timestamp 1623939100
transform 1 0 37076 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_384
timestamp 1623939100
transform 1 0 36432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _791_
timestamp 1623939100
transform 1 0 38088 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1623939100
transform 1 0 37812 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_400
timestamp 1623939100
transform 1 0 37904 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_412
timestamp 1623939100
transform 1 0 39008 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_396
timestamp 1623939100
transform 1 0 37536 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1623939100
transform 1 0 40480 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_424
timestamp 1623939100
transform 1 0 40112 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_436
timestamp 1623939100
transform 1 0 41216 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_421
timestamp 1623939100
transform 1 0 39836 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_427
timestamp 1623939100
transform 1 0 40388 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_429
timestamp 1623939100
transform 1 0 40572 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1623939100
transform 1 0 43056 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_448
timestamp 1623939100
transform 1 0 42320 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_457
timestamp 1623939100
transform 1 0 43148 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_441
timestamp 1623939100
transform 1 0 41676 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_453
timestamp 1623939100
transform 1 0 42780 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_469
timestamp 1623939100
transform 1 0 44252 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_465
timestamp 1623939100
transform 1 0 43884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_477
timestamp 1623939100
transform 1 0 44988 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1623939100
transform 1 0 45724 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_481
timestamp 1623939100
transform 1 0 45356 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_493
timestamp 1623939100
transform 1 0 46460 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_486
timestamp 1623939100
transform 1 0 45816 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_498
timestamp 1623939100
transform 1 0 46920 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1623939100
transform 1 0 48300 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1623939100
transform 1 0 47564 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_514
timestamp 1623939100
transform 1 0 48392 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_510
timestamp 1623939100
transform 1 0 48024 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _380_
timestamp 1623939100
transform 1 0 50876 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_203
timestamp 1623939100
transform 1 0 50692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_526
timestamp 1623939100
transform 1 0 49496 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_538
timestamp 1623939100
transform 1 0 50600 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_522
timestamp 1623939100
transform 1 0 49128 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_534
timestamp 1623939100
transform 1 0 50232 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _565_
timestamp 1623939100
transform 1 0 52256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _665_
timestamp 1623939100
transform 1 0 52072 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1623939100
transform 1 0 50968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_547
timestamp 1623939100
transform 1 0 51428 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_553
timestamp 1623939100
transform 1 0 51980 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_557
timestamp 1623939100
transform 1 0 52348 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_543
timestamp 1623939100
transform 1 0 51060 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_555
timestamp 1623939100
transform 1 0 52164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_559
timestamp 1623939100
transform 1 0 52532 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _376_
timestamp 1623939100
transform 1 0 54004 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1623939100
transform 1 0 53544 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_569
timestamp 1623939100
transform 1 0 53452 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_571
timestamp 1623939100
transform 1 0 53636 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_581
timestamp 1623939100
transform 1 0 54556 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_571
timestamp 1623939100
transform 1 0 53636 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_583
timestamp 1623939100
transform 1 0 54740 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1623939100
transform 1 0 56212 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_593
timestamp 1623939100
transform 1 0 55660 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_595
timestamp 1623939100
transform 1 0 55844 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_600
timestamp 1623939100
transform 1 0 56304 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _454_
timestamp 1623939100
transform 1 0 57592 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_605
timestamp 1623939100
transform 1 0 56764 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1623939100
transform 1 0 57868 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_625
timestamp 1623939100
transform 1 0 58604 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_612
timestamp 1623939100
transform 1 0 57408 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_623
timestamp 1623939100
transform 1 0 58420 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _690_
timestamp 1623939100
transform 1 0 59340 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1623939100
transform 1 0 58788 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_628
timestamp 1623939100
transform 1 0 58880 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_640
timestamp 1623939100
transform 1 0 59984 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_631
timestamp 1623939100
transform 1 0 59156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_636
timestamp 1623939100
transform 1 0 59616 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1623939100
transform 1 0 61456 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_652
timestamp 1623939100
transform 1 0 61088 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_664
timestamp 1623939100
transform 1 0 62192 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_648
timestamp 1623939100
transform 1 0 60720 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_657
timestamp 1623939100
transform 1 0 61548 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1623939100
transform 1 0 64032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_676
timestamp 1623939100
transform 1 0 63296 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_685
timestamp 1623939100
transform 1 0 64124 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_669
timestamp 1623939100
transform 1 0 62652 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_681
timestamp 1623939100
transform 1 0 63756 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_697
timestamp 1623939100
transform 1 0 65228 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_693
timestamp 1623939100
transform 1 0 64860 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_705
timestamp 1623939100
transform 1 0 65964 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _670_
timestamp 1623939100
transform 1 0 67160 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1623939100
transform 1 0 66700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_709
timestamp 1623939100
transform 1 0 66332 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_717
timestamp 1623939100
transform 1 0 67068 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_721
timestamp 1623939100
transform 1 0 67436 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_714
timestamp 1623939100
transform 1 0 66792 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_726
timestamp 1623939100
transform 1 0 67896 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1623939100
transform 1 0 69276 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_733
timestamp 1623939100
transform 1 0 68540 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_742
timestamp 1623939100
transform 1 0 69368 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_738
timestamp 1623939100
transform 1 0 69000 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_750
timestamp 1623939100
transform 1 0 70104 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1623939100
transform 1 0 71944 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_754
timestamp 1623939100
transform 1 0 70472 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_766
timestamp 1623939100
transform 1 0 71576 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_762
timestamp 1623939100
transform 1 0 71208 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_778
timestamp 1623939100
transform 1 0 72680 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_790
timestamp 1623939100
transform 1 0 73784 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_771
timestamp 1623939100
transform 1 0 72036 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_783
timestamp 1623939100
transform 1 0 73140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1623939100
transform 1 0 74520 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_799
timestamp 1623939100
transform 1 0 74612 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_811
timestamp 1623939100
transform 1 0 75716 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_795
timestamp 1623939100
transform 1 0 74244 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_807
timestamp 1623939100
transform 1 0 75348 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1623939100
transform 1 0 77188 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_823
timestamp 1623939100
transform 1 0 76820 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_819
timestamp 1623939100
transform 1 0 76452 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_828
timestamp 1623939100
transform 1 0 77280 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_835
timestamp 1623939100
transform 1 0 77924 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_847
timestamp 1623939100
transform 1 0 79028 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_840
timestamp 1623939100
transform 1 0 78384 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_852
timestamp 1623939100
transform 1 0 79488 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _293_
timestamp 1623939100
transform 1 0 81052 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1623939100
transform 1 0 79764 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_856
timestamp 1623939100
transform 1 0 79856 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_868
timestamp 1623939100
transform 1 0 80960 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_864
timestamp 1623939100
transform 1 0 80592 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_868
timestamp 1623939100
transform 1 0 80960 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1623939100
transform 1 0 82432 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_880
timestamp 1623939100
transform 1 0 82064 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_892
timestamp 1623939100
transform 1 0 83168 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_878
timestamp 1623939100
transform 1 0 81880 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_885
timestamp 1623939100
transform 1 0 82524 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1623939100
transform 1 0 85008 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_904
timestamp 1623939100
transform 1 0 84272 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_913
timestamp 1623939100
transform 1 0 85100 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_897
timestamp 1623939100
transform 1 0 83628 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_909
timestamp 1623939100
transform 1 0 84732 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_925
timestamp 1623939100
transform 1 0 86204 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_937
timestamp 1623939100
transform 1 0 87308 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_921
timestamp 1623939100
transform 1 0 85836 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_933
timestamp 1623939100
transform 1 0 86940 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1623939100
transform 1 0 87676 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_949
timestamp 1623939100
transform 1 0 88412 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_942
timestamp 1623939100
transform 1 0 87768 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_954
timestamp 1623939100
transform 1 0 88872 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _425_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 90712 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1623939100
transform 1 0 90252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_961
timestamp 1623939100
transform 1 0 89516 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_970
timestamp 1623939100
transform 1 0 90344 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_966
timestamp 1623939100
transform 1 0 89976 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_978
timestamp 1623939100
transform 1 0 91080 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1623939100
transform 1 0 92920 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_983
timestamp 1623939100
transform 1 0 91540 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_995
timestamp 1623939100
transform 1 0 92644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_990
timestamp 1623939100
transform 1 0 92184 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_999
timestamp 1623939100
transform 1 0 93012 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1007
timestamp 1623939100
transform 1 0 93748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1019
timestamp 1623939100
transform 1 0 94852 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1011
timestamp 1623939100
transform 1 0 94116 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _586_
timestamp 1623939100
transform 1 0 95680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1623939100
transform 1 0 95496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1025
timestamp 1623939100
transform 1 0 95404 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1027
timestamp 1623939100
transform 1 0 95588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1039
timestamp 1623939100
transform 1 0 96692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1023
timestamp 1623939100
transform 1 0 95220 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1027
timestamp 1623939100
transform 1 0 95588 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1031
timestamp 1623939100
transform 1 0 95956 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1623939100
transform -1 0 98808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1623939100
transform -1 0 98808 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1623939100
transform 1 0 98164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1051
timestamp 1623939100
transform 1 0 97796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1043
timestamp 1623939100
transform 1 0 97060 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_1056
timestamp 1623939100
transform 1 0 98256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1623939100
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1623939100
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1623939100
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1623939100
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1623939100
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1623939100
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1623939100
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1623939100
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1623939100
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1623939100
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1623939100
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1623939100
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_106
timestamp 1623939100
transform 1 0 10856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1623939100
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_127
timestamp 1623939100
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1623939100
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1623939100
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_163
timestamp 1623939100
transform 1 0 16100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1623939100
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1623939100
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1623939100
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1623939100
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1623939100
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1623939100
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_220
timestamp 1623939100
transform 1 0 21344 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_229
timestamp 1623939100
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_241
timestamp 1623939100
transform 1 0 23276 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_253
timestamp 1623939100
transform 1 0 24380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_265
timestamp 1623939100
transform 1 0 25484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1623939100
transform 1 0 27324 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_277
timestamp 1623939100
transform 1 0 26588 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_286
timestamp 1623939100
transform 1 0 27416 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _598_
timestamp 1623939100
transform 1 0 28152 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_297
timestamp 1623939100
transform 1 0 28428 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_309
timestamp 1623939100
transform 1 0 29532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_321
timestamp 1623939100
transform 1 0 30636 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_333
timestamp 1623939100
transform 1 0 31740 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1623939100
transform 1 0 32568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_341
timestamp 1623939100
transform 1 0 32476 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_343
timestamp 1623939100
transform 1 0 32660 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_355
timestamp 1623939100
transform 1 0 33764 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_367
timestamp 1623939100
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1623939100
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_391
timestamp 1623939100
transform 1 0 37076 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1623939100
transform 1 0 37812 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_400
timestamp 1623939100
transform 1 0 37904 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_412
timestamp 1623939100
transform 1 0 39008 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_424
timestamp 1623939100
transform 1 0 40112 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_436
timestamp 1623939100
transform 1 0 41216 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1623939100
transform 1 0 43056 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_448
timestamp 1623939100
transform 1 0 42320 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_457
timestamp 1623939100
transform 1 0 43148 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _356_
timestamp 1623939100
transform 1 0 44160 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_465
timestamp 1623939100
transform 1 0 43884 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_477
timestamp 1623939100
transform 1 0 44988 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_489
timestamp 1623939100
transform 1 0 46092 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1623939100
transform 1 0 48300 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_501
timestamp 1623939100
transform 1 0 47196 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_514
timestamp 1623939100
transform 1 0 48392 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_526
timestamp 1623939100
transform 1 0 49496 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_538
timestamp 1623939100
transform 1 0 50600 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_550
timestamp 1623939100
transform 1 0 51704 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_562
timestamp 1623939100
transform 1 0 52808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1623939100
transform 1 0 53544 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_571
timestamp 1623939100
transform 1 0 53636 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_583
timestamp 1623939100
transform 1 0 54740 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_595
timestamp 1623939100
transform 1 0 55844 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_607
timestamp 1623939100
transform 1 0 56948 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_619
timestamp 1623939100
transform 1 0 58052 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1623939100
transform 1 0 58788 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_628
timestamp 1623939100
transform 1 0 58880 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_640
timestamp 1623939100
transform 1 0 59984 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _783_
timestamp 1623939100
transform 1 0 61824 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_118
timestamp 1623939100
transform 1 0 61640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_652
timestamp 1623939100
transform 1 0 61088 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1623939100
transform 1 0 64032 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_679
timestamp 1623939100
transform 1 0 63572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_683
timestamp 1623939100
transform 1 0 63940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_685
timestamp 1623939100
transform 1 0 64124 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_8  _426_
timestamp 1623939100
transform 1 0 65228 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _583_
timestamp 1623939100
transform 1 0 67068 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_710
timestamp 1623939100
transform 1 0 66424 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_716
timestamp 1623939100
transform 1 0 66976 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_720
timestamp 1623939100
transform 1 0 67344 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _647_
timestamp 1623939100
transform 1 0 68540 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1623939100
transform 1 0 69276 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_732
timestamp 1623939100
transform 1 0 68448 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_736
timestamp 1623939100
transform 1 0 68816 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_740
timestamp 1623939100
transform 1 0 69184 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_742
timestamp 1623939100
transform 1 0 69368 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_754
timestamp 1623939100
transform 1 0 70472 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_766
timestamp 1623939100
transform 1 0 71576 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_778
timestamp 1623939100
transform 1 0 72680 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_790
timestamp 1623939100
transform 1 0 73784 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1623939100
transform 1 0 74520 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_799
timestamp 1623939100
transform 1 0 74612 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_811
timestamp 1623939100
transform 1 0 75716 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_823
timestamp 1623939100
transform 1 0 76820 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_835
timestamp 1623939100
transform 1 0 77924 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_847
timestamp 1623939100
transform 1 0 79028 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1623939100
transform 1 0 79764 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_856
timestamp 1623939100
transform 1 0 79856 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_868
timestamp 1623939100
transform 1 0 80960 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_880
timestamp 1623939100
transform 1 0 82064 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_892
timestamp 1623939100
transform 1 0 83168 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1623939100
transform 1 0 85008 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_904
timestamp 1623939100
transform 1 0 84272 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_913
timestamp 1623939100
transform 1 0 85100 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_925
timestamp 1623939100
transform 1 0 86204 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_937
timestamp 1623939100
transform 1 0 87308 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_949
timestamp 1623939100
transform 1 0 88412 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _400_
timestamp 1623939100
transform 1 0 90988 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1623939100
transform 1 0 90252 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_961
timestamp 1623939100
transform 1 0 89516 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_970
timestamp 1623939100
transform 1 0 90344 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_976
timestamp 1623939100
transform 1 0 90896 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_983
timestamp 1623939100
transform 1 0 91540 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_995
timestamp 1623939100
transform 1 0 92644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1007
timestamp 1623939100
transform 1 0 93748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1019
timestamp 1623939100
transform 1 0 94852 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1623939100
transform 1 0 95496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1025
timestamp 1623939100
transform 1 0 95404 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1027
timestamp 1623939100
transform 1 0 95588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1039
timestamp 1623939100
transform 1 0 96692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1623939100
transform -1 0 98808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1051
timestamp 1623939100
transform 1 0 97796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1623939100
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1623939100
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1623939100
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1623939100
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1623939100
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1623939100
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _751_
timestamp 1623939100
transform 1 0 6440 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1623939100
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_54
timestamp 1623939100
transform 1 0 6072 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_77
timestamp 1623939100
transform 1 0 8188 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1623939100
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1623939100
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1623939100
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1623939100
transform 1 0 10212 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _340_
timestamp 1623939100
transform -1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_138
timestamp 1623939100
transform -1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_142
timestamp 1623939100
transform -1 0 12236 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_111
timestamp 1623939100
transform 1 0 11316 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1623939100
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_139
timestamp 1623939100
transform -1 0 13432 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_134
timestamp 1623939100
transform 1 0 13432 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1623939100
transform 1 0 14168 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1623939100
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_156
timestamp 1623939100
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_168
timestamp 1623939100
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_180
timestamp 1623939100
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1623939100
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_192
timestamp 1623939100
transform 1 0 18768 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1623939100
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _645_
timestamp 1623939100
transform 1 0 21528 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_347
timestamp 1623939100
transform 1 0 21344 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_213
timestamp 1623939100
transform 1 0 20700 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1623939100
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_225
timestamp 1623939100
transform 1 0 21804 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_237
timestamp 1623939100
transform 1 0 22908 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_249
timestamp 1623939100
transform 1 0 24012 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1623939100
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 25208 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_258
timestamp 1623939100
transform 1 0 24840 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1623939100
transform 1 0 25484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _736_
timestamp 1623939100
transform 1 0 26680 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_16_277
timestamp 1623939100
transform 1 0 26588 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_297
timestamp 1623939100
transform 1 0 28428 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_309
timestamp 1623939100
transform 1 0 29532 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1623939100
transform 1 0 29992 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_313
timestamp 1623939100
transform 1 0 29900 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_315
timestamp 1623939100
transform 1 0 30084 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_327
timestamp 1623939100
transform 1 0 31188 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_339
timestamp 1623939100
transform 1 0 32292 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_351
timestamp 1623939100
transform 1 0 33396 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1623939100
transform 1 0 35236 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_363
timestamp 1623939100
transform 1 0 34500 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_372
timestamp 1623939100
transform 1 0 35328 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_384
timestamp 1623939100
transform 1 0 36432 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _524_
timestamp 1623939100
transform 1 0 38180 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _640_
timestamp 1623939100
transform 1 0 37536 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_399
timestamp 1623939100
transform 1 0 37812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1623939100
transform 1 0 40480 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_419
timestamp 1623939100
transform 1 0 39652 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_427
timestamp 1623939100
transform 1 0 40388 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_429
timestamp 1623939100
transform 1 0 40572 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _600_
timestamp 1623939100
transform 1 0 42412 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_441
timestamp 1623939100
transform 1 0 41676 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_452
timestamp 1623939100
transform 1 0 42688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_464
timestamp 1623939100
transform 1 0 43792 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_476
timestamp 1623939100
transform 1 0 44896 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1623939100
transform 1 0 45724 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_484
timestamp 1623939100
transform 1 0 45632 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_486
timestamp 1623939100
transform 1 0 45816 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_498
timestamp 1623939100
transform 1 0 46920 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_510
timestamp 1623939100
transform 1 0 48024 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_522
timestamp 1623939100
transform 1 0 49128 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_534
timestamp 1623939100
transform 1 0 50232 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1623939100
transform 1 0 50968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_543
timestamp 1623939100
transform 1 0 51060 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_555
timestamp 1623939100
transform 1 0 52164 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_567
timestamp 1623939100
transform 1 0 53268 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_579
timestamp 1623939100
transform 1 0 54372 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1623939100
transform 1 0 56212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_591
timestamp 1623939100
transform 1 0 55476 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_600
timestamp 1623939100
transform 1 0 56304 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_612
timestamp 1623939100
transform 1 0 57408 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_624
timestamp 1623939100
transform 1 0 58512 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_636
timestamp 1623939100
transform 1 0 59616 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1623939100
transform 1 0 61456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_648
timestamp 1623939100
transform 1 0 60720 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_657
timestamp 1623939100
transform 1 0 61548 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_669
timestamp 1623939100
transform 1 0 62652 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_681
timestamp 1623939100
transform 1 0 63756 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_693
timestamp 1623939100
transform 1 0 64860 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_705
timestamp 1623939100
transform 1 0 65964 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  _509_
timestamp 1623939100
transform 1 0 67160 0 -1 11424
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1623939100
transform 1 0 66700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_714
timestamp 1623939100
transform 1 0 66792 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_729
timestamp 1623939100
transform 1 0 68172 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _287_
timestamp 1623939100
transform 1 0 69092 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_737
timestamp 1623939100
transform 1 0 68908 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_745
timestamp 1623939100
transform 1 0 69644 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1623939100
transform 1 0 71944 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_757
timestamp 1623939100
transform 1 0 70748 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_769
timestamp 1623939100
transform 1 0 71852 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_771
timestamp 1623939100
transform 1 0 72036 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_783
timestamp 1623939100
transform 1 0 73140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_795
timestamp 1623939100
transform 1 0 74244 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_807
timestamp 1623939100
transform 1 0 75348 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1623939100
transform 1 0 77188 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_819
timestamp 1623939100
transform 1 0 76452 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_828
timestamp 1623939100
transform 1 0 77280 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_840
timestamp 1623939100
transform 1 0 78384 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_852
timestamp 1623939100
transform 1 0 79488 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_864
timestamp 1623939100
transform 1 0 80592 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1623939100
transform 1 0 82432 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_876
timestamp 1623939100
transform 1 0 81696 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_885
timestamp 1623939100
transform 1 0 82524 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_897
timestamp 1623939100
transform 1 0 83628 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_909
timestamp 1623939100
transform 1 0 84732 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_921
timestamp 1623939100
transform 1 0 85836 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_933
timestamp 1623939100
transform 1 0 86940 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1623939100
transform 1 0 87676 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_942
timestamp 1623939100
transform 1 0 87768 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_954
timestamp 1623939100
transform 1 0 88872 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_966
timestamp 1623939100
transform 1 0 89976 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_978
timestamp 1623939100
transform 1 0 91080 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1623939100
transform 1 0 92920 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_990
timestamp 1623939100
transform 1 0 92184 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_999
timestamp 1623939100
transform 1 0 93012 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1011
timestamp 1623939100
transform 1 0 94116 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _511_
timestamp 1623939100
transform 1 0 96324 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_193
timestamp 1623939100
transform 1 0 96140 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1023
timestamp 1623939100
transform 1 0 95220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1031
timestamp 1623939100
transform 1 0 95956 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1623939100
transform -1 0 98808 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1623939100
transform 1 0 98164 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1051
timestamp 1623939100
transform 1 0 97796 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_1056
timestamp 1623939100
transform 1 0 98256 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1623939100
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1623939100
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1623939100
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1623939100
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1623939100
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _767_
timestamp 1623939100
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1623939100
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1623939100
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_58
timestamp 1623939100
transform 1 0 6440 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1623939100
transform 1 0 8556 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _671_
timestamp 1623939100
transform 1 0 10120 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1623939100
transform 1 0 9660 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_97
timestamp 1623939100
transform 1 0 10028 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_101
timestamp 1623939100
transform 1 0 10396 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _446_
timestamp 1623939100
transform 1 0 12604 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1623939100
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1623939100
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_115
timestamp 1623939100
transform 1 0 11684 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1623939100
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1623939100
transform 1 0 13708 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_wb_clk_i
timestamp 1623939100
transform 1 0 14996 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_149
timestamp 1623939100
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_154
timestamp 1623939100
transform 1 0 15272 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_166
timestamp 1623939100
transform 1 0 16376 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1623939100
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_170
timestamp 1623939100
transform 1 0 16744 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1623939100
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1623939100
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1623939100
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1623939100
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1623939100
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_220
timestamp 1623939100
transform 1 0 21344 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1623939100
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_241
timestamp 1623939100
transform 1 0 23276 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_253
timestamp 1623939100
transform 1 0 24380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_265
timestamp 1623939100
transform 1 0 25484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  _526_
timestamp 1623939100
transform 1 0 27784 0 1 11424
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1623939100
transform 1 0 27324 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_277
timestamp 1623939100
transform 1 0 26588 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_286
timestamp 1623939100
transform 1 0 27416 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_301
timestamp 1623939100
transform 1 0 28796 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_313
timestamp 1623939100
transform 1 0 29900 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_325
timestamp 1623939100
transform 1 0 31004 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1623939100
transform 1 0 32568 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1623939100
transform 1 0 32108 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_341
timestamp 1623939100
transform 1 0 32476 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_343
timestamp 1623939100
transform 1 0 32660 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_wb_clk_i
timestamp 1623939100
transform 1 0 34868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_355
timestamp 1623939100
transform 1 0 33764 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_370
timestamp 1623939100
transform 1 0 35144 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_382
timestamp 1623939100
transform 1 0 36248 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_394
timestamp 1623939100
transform 1 0 37352 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _469_
timestamp 1623939100
transform 1 0 38364 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1623939100
transform 1 0 37812 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_163
timestamp 1623939100
transform 1 0 38180 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_398
timestamp 1623939100
transform 1 0 37720 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_400
timestamp 1623939100
transform 1 0 37904 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_414
timestamp 1623939100
transform 1 0 39192 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_426
timestamp 1623939100
transform 1 0 40296 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1623939100
transform 1 0 43056 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_438
timestamp 1623939100
transform 1 0 41400 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_450
timestamp 1623939100
transform 1 0 42504 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_457
timestamp 1623939100
transform 1 0 43148 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_469
timestamp 1623939100
transform 1 0 44252 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_481
timestamp 1623939100
transform 1 0 45356 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_493
timestamp 1623939100
transform 1 0 46460 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1623939100
transform 1 0 48300 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1623939100
transform 1 0 47564 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_514
timestamp 1623939100
transform 1 0 48392 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_526
timestamp 1623939100
transform 1 0 49496 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_538
timestamp 1623939100
transform 1 0 50600 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_550
timestamp 1623939100
transform 1 0 51704 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_562
timestamp 1623939100
transform 1 0 52808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1623939100
transform 1 0 53544 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_571
timestamp 1623939100
transform 1 0 53636 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_583
timestamp 1623939100
transform 1 0 54740 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_595
timestamp 1623939100
transform 1 0 55844 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_607
timestamp 1623939100
transform 1 0 56948 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_619
timestamp 1623939100
transform 1 0 58052 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1623939100
transform 1 0 58788 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_628
timestamp 1623939100
transform 1 0 58880 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_640
timestamp 1623939100
transform 1 0 59984 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_652
timestamp 1623939100
transform 1 0 61088 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_664
timestamp 1623939100
transform 1 0 62192 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1623939100
transform 1 0 64032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_676
timestamp 1623939100
transform 1 0 63296 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_685
timestamp 1623939100
transform 1 0 64124 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_697
timestamp 1623939100
transform 1 0 65228 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_709
timestamp 1623939100
transform 1 0 66332 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_721
timestamp 1623939100
transform 1 0 67436 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1623939100
transform 1 0 69276 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_733
timestamp 1623939100
transform 1 0 68540 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_742
timestamp 1623939100
transform 1 0 69368 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_754
timestamp 1623939100
transform 1 0 70472 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_766
timestamp 1623939100
transform 1 0 71576 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_778
timestamp 1623939100
transform 1 0 72680 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_790
timestamp 1623939100
transform 1 0 73784 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _384_
timestamp 1623939100
transform 1 0 74980 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1623939100
transform 1 0 74520 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_799
timestamp 1623939100
transform 1 0 74612 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_812
timestamp 1623939100
transform 1 0 75808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_824
timestamp 1623939100
transform 1 0 76912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_836
timestamp 1623939100
transform 1 0 78016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_848
timestamp 1623939100
transform 1 0 79120 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_854
timestamp 1623939100
transform 1 0 79672 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1623939100
transform 1 0 79764 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_856
timestamp 1623939100
transform 1 0 79856 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_868
timestamp 1623939100
transform 1 0 80960 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_880
timestamp 1623939100
transform 1 0 82064 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_892
timestamp 1623939100
transform 1 0 83168 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1623939100
transform 1 0 85008 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_904
timestamp 1623939100
transform 1 0 84272 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_913
timestamp 1623939100
transform 1 0 85100 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_wb_clk_i
timestamp 1623939100
transform 1 0 85468 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_920
timestamp 1623939100
transform 1 0 85744 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_932
timestamp 1623939100
transform 1 0 86848 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_944
timestamp 1623939100
transform 1 0 87952 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_956
timestamp 1623939100
transform 1 0 89056 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _576_
timestamp 1623939100
transform 1 0 90804 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1623939100
transform 1 0 90252 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_968
timestamp 1623939100
transform 1 0 90160 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_970
timestamp 1623939100
transform 1 0 90344 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_974
timestamp 1623939100
transform 1 0 90712 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_978
timestamp 1623939100
transform 1 0 91080 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_990
timestamp 1623939100
transform 1 0 92184 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1002
timestamp 1623939100
transform 1 0 93288 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1014
timestamp 1623939100
transform 1 0 94392 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1623939100
transform 1 0 95496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1027
timestamp 1623939100
transform 1 0 95588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1039
timestamp 1623939100
transform 1 0 96692 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _633_
timestamp 1623939100
transform 1 0 97428 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1623939100
transform -1 0 98808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1050
timestamp 1623939100
transform 1 0 97704 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1058
timestamp 1623939100
transform 1 0 98440 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1623939100
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1623939100
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1623939100
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _601_
timestamp 1623939100
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1623939100
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1623939100
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_30
timestamp 1623939100
transform 1 0 3864 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_37
timestamp 1623939100
transform 1 0 4508 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_49
timestamp 1623939100
transform 1 0 5612 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_61
timestamp 1623939100
transform 1 0 6716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_73
timestamp 1623939100
transform 1 0 7820 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _695_
timestamp 1623939100
transform 1 0 10672 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1623939100
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_291
timestamp 1623939100
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1623939100
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1623939100
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_99
timestamp 1623939100
transform 1 0 10212 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_107
timestamp 1623939100
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_119
timestamp 1623939100
transform 1 0 12052 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1623939100
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_131
timestamp 1623939100
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1623939100
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_156
timestamp 1623939100
transform 1 0 15456 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _280_
timestamp 1623939100
transform 1 0 17572 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_168
timestamp 1623939100
transform 1 0 16560 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_176
timestamp 1623939100
transform 1 0 17296 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1623939100
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_188
timestamp 1623939100
transform 1 0 18400 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1623939100
transform 1 0 19596 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_213
timestamp 1623939100
transform 1 0 20700 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_225
timestamp 1623939100
transform 1 0 21804 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_237
timestamp 1623939100
transform 1 0 22908 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_249
timestamp 1623939100
transform 1 0 24012 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1623939100
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_258
timestamp 1623939100
transform 1 0 24840 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_270
timestamp 1623939100
transform 1 0 25944 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_282
timestamp 1623939100
transform 1 0 27048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_294
timestamp 1623939100
transform 1 0 28152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_306
timestamp 1623939100
transform 1 0 29256 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1623939100
transform 1 0 29992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_315
timestamp 1623939100
transform 1 0 30084 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_327
timestamp 1623939100
transform 1 0 31188 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_339
timestamp 1623939100
transform 1 0 32292 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_351
timestamp 1623939100
transform 1 0 33396 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1623939100
transform 1 0 35236 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_363
timestamp 1623939100
transform 1 0 34500 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_372
timestamp 1623939100
transform 1 0 35328 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_384
timestamp 1623939100
transform 1 0 36432 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_396
timestamp 1623939100
transform 1 0 37536 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_408
timestamp 1623939100
transform 1 0 38640 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1623939100
transform 1 0 40480 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_420
timestamp 1623939100
transform 1 0 39744 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_429
timestamp 1623939100
transform 1 0 40572 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _326_
timestamp 1623939100
transform 1 0 42504 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_18_441
timestamp 1623939100
transform 1 0 41676 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_449
timestamp 1623939100
transform 1 0 42412 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1623939100
transform 1 0 43148 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_469
timestamp 1623939100
transform 1 0 44252 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _733_
timestamp 1623939100
transform 1 0 46184 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1623939100
transform 1 0 45724 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_481
timestamp 1623939100
transform 1 0 45356 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_486
timestamp 1623939100
transform 1 0 45816 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_509
timestamp 1623939100
transform 1 0 47932 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_521
timestamp 1623939100
transform 1 0 49036 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_533
timestamp 1623939100
transform 1 0 50140 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_541
timestamp 1623939100
transform 1 0 50876 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1623939100
transform 1 0 50968 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_543
timestamp 1623939100
transform 1 0 51060 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_555
timestamp 1623939100
transform 1 0 52164 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_567
timestamp 1623939100
transform 1 0 53268 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_579
timestamp 1623939100
transform 1 0 54372 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1623939100
transform 1 0 56212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_591
timestamp 1623939100
transform 1 0 55476 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_600
timestamp 1623939100
transform 1 0 56304 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _491_
timestamp 1623939100
transform 1 0 58420 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _581_
timestamp 1623939100
transform 1 0 57500 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_612
timestamp 1623939100
transform 1 0 57408 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_616
timestamp 1623939100
transform 1 0 57776 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_622
timestamp 1623939100
transform 1 0 58328 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_639
timestamp 1623939100
transform 1 0 59892 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _463_
timestamp 1623939100
transform 1 0 62192 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1623939100
transform 1 0 61456 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_651
timestamp 1623939100
transform 1 0 60996 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_655
timestamp 1623939100
transform 1 0 61364 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_657
timestamp 1623939100
transform 1 0 61548 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_663
timestamp 1623939100
transform 1 0 62100 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_670
timestamp 1623939100
transform 1 0 62744 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_682
timestamp 1623939100
transform 1 0 63848 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _602_
timestamp 1623939100
transform 1 0 65136 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_wb_clk_i
timestamp 1623939100
transform 1 0 65780 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_694
timestamp 1623939100
transform 1 0 64952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_699
timestamp 1623939100
transform 1 0 65412 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_706
timestamp 1623939100
transform 1 0 66056 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _691_
timestamp 1623939100
transform 1 0 67160 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1623939100
transform 1 0 66700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_712
timestamp 1623939100
transform 1 0 66608 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_714
timestamp 1623939100
transform 1 0 66792 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_721
timestamp 1623939100
transform 1 0 67436 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_733
timestamp 1623939100
transform 1 0 68540 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_745
timestamp 1623939100
transform 1 0 69644 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1623939100
transform 1 0 71944 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_757
timestamp 1623939100
transform 1 0 70748 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_769
timestamp 1623939100
transform 1 0 71852 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _570_
timestamp 1623939100
transform 1 0 72404 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_771
timestamp 1623939100
transform 1 0 72036 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_778
timestamp 1623939100
transform 1 0 72680 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_790
timestamp 1623939100
transform 1 0 73784 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_802
timestamp 1623939100
transform 1 0 74888 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1623939100
transform 1 0 77188 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_814
timestamp 1623939100
transform 1 0 75992 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_826
timestamp 1623939100
transform 1 0 77096 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_828
timestamp 1623939100
transform 1 0 77280 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_840
timestamp 1623939100
transform 1 0 78384 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_852
timestamp 1623939100
transform 1 0 79488 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_864
timestamp 1623939100
transform 1 0 80592 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1623939100
transform 1 0 82432 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_876
timestamp 1623939100
transform 1 0 81696 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_885
timestamp 1623939100
transform 1 0 82524 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_897
timestamp 1623939100
transform 1 0 83628 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_909
timestamp 1623939100
transform 1 0 84732 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_921
timestamp 1623939100
transform 1 0 85836 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_933
timestamp 1623939100
transform 1 0 86940 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1623939100
transform 1 0 87676 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_942
timestamp 1623939100
transform 1 0 87768 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_954
timestamp 1623939100
transform 1 0 88872 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_966
timestamp 1623939100
transform 1 0 89976 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_978
timestamp 1623939100
transform 1 0 91080 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1623939100
transform 1 0 92920 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_990
timestamp 1623939100
transform 1 0 92184 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_999
timestamp 1623939100
transform 1 0 93012 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1011
timestamp 1623939100
transform 1 0 94116 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1023
timestamp 1623939100
transform 1 0 95220 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1035
timestamp 1623939100
transform 1 0 96324 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1623939100
transform -1 0 98808 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1623939100
transform 1 0 98164 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1047
timestamp 1623939100
transform 1 0 97428 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_1056
timestamp 1623939100
transform 1 0 98256 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1623939100
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1623939100
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1623939100
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1623939100
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1623939100
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1623939100
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1623939100
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1623939100
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1623939100
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1623939100
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1623939100
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1623939100
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1623939100
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1623939100
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1623939100
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1623939100
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _713_
timestamp 1623939100
transform 1 0 7636 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_19_70
timestamp 1623939100
transform 1 0 7544 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_66
timestamp 1623939100
transform 1 0 7176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1623939100
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1623939100
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_90
timestamp 1623939100
transform 1 0 9384 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_102
timestamp 1623939100
transform 1 0 10488 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1623939100
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1623939100
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1623939100
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_232
timestamp 1623939100
transform -1 0 12696 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_115
timestamp 1623939100
transform 1 0 11684 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_123
timestamp 1623939100
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1623939100
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1623939100
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _498_
timestamp 1623939100
transform -1 0 13524 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1623939100
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1623939100
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1623939100
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1623939100
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1623939100
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1623939100
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1623939100
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1623939100
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1623939100
transform 1 0 16928 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1623939100
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1623939100
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_180
timestamp 1623939100
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1623939100
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1623939100
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1623939100
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_192
timestamp 1623939100
transform 1 0 18768 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1623939100
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1623939100
transform 1 0 22080 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_220
timestamp 1623939100
transform 1 0 21344 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_229
timestamp 1623939100
transform 1 0 22172 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_213
timestamp 1623939100
transform 1 0 20700 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_225
timestamp 1623939100
transform 1 0 21804 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _289_
timestamp 1623939100
transform -1 0 23092 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_131
timestamp 1623939100
transform -1 0 22540 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_239
timestamp 1623939100
transform 1 0 23092 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_237
timestamp 1623939100
transform 1 0 22908 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_249
timestamp 1623939100
transform 1 0 24012 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1623939100
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_251
timestamp 1623939100
transform 1 0 24196 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_263
timestamp 1623939100
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_258
timestamp 1623939100
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_270
timestamp 1623939100
transform 1 0 25944 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _377_
timestamp 1623939100
transform 1 0 26864 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1623939100
transform 1 0 27324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_275
timestamp 1623939100
transform 1 0 26404 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_283
timestamp 1623939100
transform 1 0 27140 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_286
timestamp 1623939100
transform 1 0 27416 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_278
timestamp 1623939100
transform 1 0 26680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_287
timestamp 1623939100
transform 1 0 27508 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_298
timestamp 1623939100
transform 1 0 28520 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_310
timestamp 1623939100
transform 1 0 29624 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_299
timestamp 1623939100
transform 1 0 28612 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_311
timestamp 1623939100
transform 1 0 29716 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1623939100
transform 1 0 29992 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_322
timestamp 1623939100
transform 1 0 30728 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_315
timestamp 1623939100
transform 1 0 30084 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_327
timestamp 1623939100
transform 1 0 31188 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1623939100
transform 1 0 32568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_334
timestamp 1623939100
transform 1 0 31832 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_343
timestamp 1623939100
transform 1 0 32660 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_339
timestamp 1623939100
transform 1 0 32292 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_351
timestamp 1623939100
transform 1 0 33396 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1623939100
transform 1 0 35236 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_355
timestamp 1623939100
transform 1 0 33764 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_367
timestamp 1623939100
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_363
timestamp 1623939100
transform 1 0 34500 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_372
timestamp 1623939100
transform 1 0 35328 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_379
timestamp 1623939100
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_391
timestamp 1623939100
transform 1 0 37076 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_384
timestamp 1623939100
transform 1 0 36432 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1623939100
transform 1 0 37812 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_400
timestamp 1623939100
transform 1 0 37904 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_412
timestamp 1623939100
transform 1 0 39008 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_396
timestamp 1623939100
transform 1 0 37536 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_408
timestamp 1623939100
transform 1 0 38640 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1623939100
transform 1 0 40480 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_424
timestamp 1623939100
transform 1 0 40112 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_436
timestamp 1623939100
transform 1 0 41216 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_420
timestamp 1623939100
transform 1 0 39744 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_429
timestamp 1623939100
transform 1 0 40572 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1623939100
transform 1 0 43056 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_448
timestamp 1623939100
transform 1 0 42320 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_457
timestamp 1623939100
transform 1 0 43148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_441
timestamp 1623939100
transform 1 0 41676 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_453
timestamp 1623939100
transform 1 0 42780 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _740_
timestamp 1623939100
transform 1 0 43516 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_59
timestamp 1623939100
transform 1 0 43332 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_465
timestamp 1623939100
transform 1 0 43884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_477
timestamp 1623939100
transform 1 0 44988 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1623939100
transform 1 0 45724 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_480
timestamp 1623939100
transform 1 0 45264 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_492
timestamp 1623939100
transform 1 0 46368 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_486
timestamp 1623939100
transform 1 0 45816 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_498
timestamp 1623939100
transform 1 0 46920 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1623939100
transform 1 0 48300 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_504
timestamp 1623939100
transform 1 0 47472 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_512
timestamp 1623939100
transform 1 0 48208 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_514
timestamp 1623939100
transform 1 0 48392 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_510
timestamp 1623939100
transform 1 0 48024 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_526
timestamp 1623939100
transform 1 0 49496 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_538
timestamp 1623939100
transform 1 0 50600 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_522
timestamp 1623939100
transform 1 0 49128 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_534
timestamp 1623939100
transform 1 0 50232 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _686_
timestamp 1623939100
transform 1 0 51888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1623939100
transform 1 0 50968 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_550
timestamp 1623939100
transform 1 0 51704 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_562
timestamp 1623939100
transform 1 0 52808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_543
timestamp 1623939100
transform 1 0 51060 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_551
timestamp 1623939100
transform 1 0 51796 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_555
timestamp 1623939100
transform 1 0 52164 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1623939100
transform 1 0 53544 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_571
timestamp 1623939100
transform 1 0 53636 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_583
timestamp 1623939100
transform 1 0 54740 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_567
timestamp 1623939100
transform 1 0 53268 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_579
timestamp 1623939100
transform 1 0 54372 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1623939100
transform 1 0 56212 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_595
timestamp 1623939100
transform 1 0 55844 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_591
timestamp 1623939100
transform 1 0 55476 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_600
timestamp 1623939100
transform 1 0 56304 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_607
timestamp 1623939100
transform 1 0 56948 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_619
timestamp 1623939100
transform 1 0 58052 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_612
timestamp 1623939100
transform 1 0 57408 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_624
timestamp 1623939100
transform 1 0 58512 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1623939100
transform 1 0 58788 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_628
timestamp 1623939100
transform 1 0 58880 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_640
timestamp 1623939100
transform 1 0 59984 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_636
timestamp 1623939100
transform 1 0 59616 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1623939100
transform 1 0 61456 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_652
timestamp 1623939100
transform 1 0 61088 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_664
timestamp 1623939100
transform 1 0 62192 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_648
timestamp 1623939100
transform 1 0 60720 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_657
timestamp 1623939100
transform 1 0 61548 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1623939100
transform 1 0 64032 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_676
timestamp 1623939100
transform 1 0 63296 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_685
timestamp 1623939100
transform 1 0 64124 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_669
timestamp 1623939100
transform 1 0 62652 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_681
timestamp 1623939100
transform 1 0 63756 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_697
timestamp 1623939100
transform 1 0 65228 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_693
timestamp 1623939100
transform 1 0 64860 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_705
timestamp 1623939100
transform 1 0 65964 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _504_
timestamp 1623939100
transform 1 0 66332 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1623939100
transform 1 0 66700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_718
timestamp 1623939100
transform 1 0 67160 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_714
timestamp 1623939100
transform 1 0 66792 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_726
timestamp 1623939100
transform 1 0 67896 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1623939100
transform 1 0 69276 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_730
timestamp 1623939100
transform 1 0 68264 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_738
timestamp 1623939100
transform 1 0 69000 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_742
timestamp 1623939100
transform 1 0 69368 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_738
timestamp 1623939100
transform 1 0 69000 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_750
timestamp 1623939100
transform 1 0 70104 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _697_
timestamp 1623939100
transform 1 0 71300 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1623939100
transform 1 0 71944 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_754
timestamp 1623939100
transform 1 0 70472 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_762
timestamp 1623939100
transform 1 0 71208 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_762
timestamp 1623939100
transform 1 0 71208 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _365_
timestamp 1623939100
transform 1 0 72680 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_782
timestamp 1623939100
transform 1 0 73048 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_771
timestamp 1623939100
transform 1 0 72036 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_777
timestamp 1623939100
transform 1 0 72588 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_787
timestamp 1623939100
transform 1 0 73508 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1623939100
transform 1 0 74520 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1623939100
transform 1 0 75440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_794
timestamp 1623939100
transform 1 0 74152 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_799
timestamp 1623939100
transform 1 0 74612 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_807
timestamp 1623939100
transform 1 0 75348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_811
timestamp 1623939100
transform 1 0 75716 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_799
timestamp 1623939100
transform 1 0 74612 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_811
timestamp 1623939100
transform 1 0 75716 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1623939100
transform 1 0 77188 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_823
timestamp 1623939100
transform 1 0 76820 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_823
timestamp 1623939100
transform 1 0 76820 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_828
timestamp 1623939100
transform 1 0 77280 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_835
timestamp 1623939100
transform 1 0 77924 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_847
timestamp 1623939100
transform 1 0 79028 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_840
timestamp 1623939100
transform 1 0 78384 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_852
timestamp 1623939100
transform 1 0 79488 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _582_
timestamp 1623939100
transform 1 0 81420 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1623939100
transform 1 0 79764 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_856
timestamp 1623939100
transform 1 0 79856 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_868
timestamp 1623939100
transform 1 0 80960 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_864
timestamp 1623939100
transform 1 0 80592 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_872
timestamp 1623939100
transform 1 0 81328 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _501_
timestamp 1623939100
transform 1 0 82892 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1623939100
transform 1 0 82432 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_880
timestamp 1623939100
transform 1 0 82064 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_892
timestamp 1623939100
transform 1 0 83168 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_876
timestamp 1623939100
transform 1 0 81696 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_885
timestamp 1623939100
transform 1 0 82524 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1623939100
transform 1 0 85008 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_173
timestamp 1623939100
transform 1 0 85284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_904
timestamp 1623939100
transform 1 0 84272 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_913
timestamp 1623939100
transform 1 0 85100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_898
timestamp 1623939100
transform 1 0 83720 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_910
timestamp 1623939100
transform 1 0 84824 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _527_
timestamp 1623939100
transform 1 0 85468 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_174
timestamp 1623939100
transform 1 0 86296 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_928
timestamp 1623939100
transform 1 0 86480 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_922
timestamp 1623939100
transform 1 0 85928 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_934
timestamp 1623939100
transform 1 0 87032 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1623939100
transform 1 0 87676 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_940
timestamp 1623939100
transform 1 0 87584 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_952
timestamp 1623939100
transform 1 0 88688 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_940
timestamp 1623939100
transform 1 0 87584 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_942
timestamp 1623939100
transform 1 0 87768 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_954
timestamp 1623939100
transform 1 0 88872 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1623939100
transform 1 0 90252 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_964
timestamp 1623939100
transform 1 0 89792 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_968
timestamp 1623939100
transform 1 0 90160 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_970
timestamp 1623939100
transform 1 0 90344 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_966
timestamp 1623939100
transform 1 0 89976 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_978
timestamp 1623939100
transform 1 0 91080 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1623939100
transform 1 0 92920 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_982
timestamp 1623939100
transform 1 0 91448 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_994
timestamp 1623939100
transform 1 0 92552 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_990
timestamp 1623939100
transform 1 0 92184 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_999
timestamp 1623939100
transform 1 0 93012 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _643_
timestamp 1623939100
transform 1 0 95036 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1006
timestamp 1623939100
transform 1 0 93656 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1018
timestamp 1623939100
transform 1 0 94760 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1011
timestamp 1623939100
transform 1 0 94116 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_1019
timestamp 1623939100
transform 1 0 94852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _641_
timestamp 1623939100
transform 1 0 96324 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1623939100
transform 1 0 95496 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1027
timestamp 1623939100
transform 1 0 95588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1038
timestamp 1623939100
transform 1 0 96600 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1024
timestamp 1623939100
transform 1 0 95312 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1036
timestamp 1623939100
transform 1 0 96416 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1623939100
transform -1 0 98808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1623939100
transform -1 0 98808 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1623939100
transform 1 0 98164 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1050
timestamp 1623939100
transform 1 0 97704 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1058
timestamp 1623939100
transform 1 0 98440 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1048
timestamp 1623939100
transform 1 0 97520 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1054
timestamp 1623939100
transform 1 0 98072 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_1056
timestamp 1623939100
transform 1 0 98256 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1623939100
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1623939100
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1623939100
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1623939100
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1623939100
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1623939100
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1623939100
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1623939100
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1623939100
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_82
timestamp 1623939100
transform 1 0 8648 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _312_
timestamp 1623939100
transform 1 0 9660 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_90
timestamp 1623939100
transform 1 0 9384 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_102
timestamp 1623939100
transform 1 0 10488 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1623939100
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1623939100
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1623939100
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1623939100
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1623939100
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1623939100
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1623939100
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_172
timestamp 1623939100
transform 1 0 16928 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1623939100
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1623939100
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1623939100
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1623939100
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_220
timestamp 1623939100
transform 1 0 21344 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_229
timestamp 1623939100
transform 1 0 22172 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_241
timestamp 1623939100
transform 1 0 23276 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_253
timestamp 1623939100
transform 1 0 24380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_265
timestamp 1623939100
transform 1 0 25484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1623939100
transform 1 0 27324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_277
timestamp 1623939100
transform 1 0 26588 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_286
timestamp 1623939100
transform 1 0 27416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_298
timestamp 1623939100
transform 1 0 28520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_310
timestamp 1623939100
transform 1 0 29624 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_322
timestamp 1623939100
transform 1 0 30728 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1623939100
transform 1 0 32568 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_334
timestamp 1623939100
transform 1 0 31832 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_343
timestamp 1623939100
transform 1 0 32660 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_355
timestamp 1623939100
transform 1 0 33764 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_367
timestamp 1623939100
transform 1 0 34868 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1623939100
transform 1 0 35972 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_391
timestamp 1623939100
transform 1 0 37076 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1623939100
transform 1 0 37812 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_400
timestamp 1623939100
transform 1 0 37904 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_412
timestamp 1623939100
transform 1 0 39008 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _563_
timestamp 1623939100
transform 1 0 40664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_424
timestamp 1623939100
transform 1 0 40112 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_433
timestamp 1623939100
transform 1 0 40940 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1623939100
transform 1 0 43056 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_445
timestamp 1623939100
transform 1 0 42044 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_453
timestamp 1623939100
transform 1 0 42780 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_457
timestamp 1623939100
transform 1 0 43148 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _334_
timestamp 1623939100
transform 1 0 43516 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_469
timestamp 1623939100
transform 1 0 44252 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_481
timestamp 1623939100
transform 1 0 45356 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_493
timestamp 1623939100
transform 1 0 46460 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1623939100
transform 1 0 48300 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1623939100
transform 1 0 47564 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_514
timestamp 1623939100
transform 1 0 48392 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _678_
timestamp 1623939100
transform 1 0 49312 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_522
timestamp 1623939100
transform 1 0 49128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_527
timestamp 1623939100
transform 1 0 49588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_539
timestamp 1623939100
transform 1 0 50692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_551
timestamp 1623939100
transform 1 0 51796 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1623939100
transform 1 0 53544 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_563
timestamp 1623939100
transform 1 0 52900 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_569
timestamp 1623939100
transform 1 0 53452 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_571
timestamp 1623939100
transform 1 0 53636 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_583
timestamp 1623939100
transform 1 0 54740 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_4  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 55292 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_605
timestamp 1623939100
transform 1 0 56764 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1623939100
transform 1 0 57868 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_625
timestamp 1623939100
transform 1 0 58604 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1623939100
transform 1 0 58788 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_628
timestamp 1623939100
transform 1 0 58880 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_640
timestamp 1623939100
transform 1 0 59984 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_652
timestamp 1623939100
transform 1 0 61088 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_664
timestamp 1623939100
transform 1 0 62192 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1623939100
transform 1 0 64032 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_676
timestamp 1623939100
transform 1 0 63296 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_685
timestamp 1623939100
transform 1 0 64124 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_2  _410_
timestamp 1623939100
transform -1 0 66792 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_223
timestamp 1623939100
transform -1 0 66148 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_697
timestamp 1623939100
transform 1 0 65228 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_714
timestamp 1623939100
transform 1 0 66792 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_726
timestamp 1623939100
transform 1 0 67896 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _651_
timestamp 1623939100
transform 1 0 69736 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1623939100
transform 1 0 69276 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_738
timestamp 1623939100
transform 1 0 69000 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_742
timestamp 1623939100
transform 1 0 69368 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_749
timestamp 1623939100
transform 1 0 70012 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_761
timestamp 1623939100
transform 1 0 71116 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _521_
timestamp 1623939100
transform 1 0 72680 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_773
timestamp 1623939100
transform 1 0 72220 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_777
timestamp 1623939100
transform 1 0 72588 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1623939100
transform 1 0 74520 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_794
timestamp 1623939100
transform 1 0 74152 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_799
timestamp 1623939100
transform 1 0 74612 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_811
timestamp 1623939100
transform 1 0 75716 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_823
timestamp 1623939100
transform 1 0 76820 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_835
timestamp 1623939100
transform 1 0 77924 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_847
timestamp 1623939100
transform 1 0 79028 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1623939100
transform 1 0 79764 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_856
timestamp 1623939100
transform 1 0 79856 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_868
timestamp 1623939100
transform 1 0 80960 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  _442_
timestamp 1623939100
transform 1 0 81972 0 1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_21_876
timestamp 1623939100
transform 1 0 81696 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_890
timestamp 1623939100
transform 1 0 82984 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1623939100
transform 1 0 85008 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_902
timestamp 1623939100
transform 1 0 84088 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_910
timestamp 1623939100
transform 1 0 84824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_913
timestamp 1623939100
transform 1 0 85100 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_925
timestamp 1623939100
transform 1 0 86204 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_937
timestamp 1623939100
transform 1 0 87308 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_949
timestamp 1623939100
transform 1 0 88412 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1623939100
transform 1 0 90252 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_961
timestamp 1623939100
transform 1 0 89516 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_970
timestamp 1623939100
transform 1 0 90344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_982
timestamp 1623939100
transform 1 0 91448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_994
timestamp 1623939100
transform 1 0 92552 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1006
timestamp 1623939100
transform 1 0 93656 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_1018
timestamp 1623939100
transform 1 0 94760 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_4  _447_
timestamp 1623939100
transform 1 0 96600 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1623939100
transform 1 0 95496 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_195
timestamp 1623939100
transform 1 0 96416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_1027
timestamp 1623939100
transform 1 0 95588 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1035
timestamp 1623939100
transform 1 0 96324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1623939100
transform -1 0 98808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_1054
timestamp 1623939100
transform 1 0 98072 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1058
timestamp 1623939100
transform 1 0 98440 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1623939100
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1623939100
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1623939100
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1623939100
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1623939100
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1623939100
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _779_
timestamp 1623939100
transform 1 0 5060 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_22_42
timestamp 1623939100
transform 1 0 4968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_62
timestamp 1623939100
transform 1 0 6808 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_74
timestamp 1623939100
transform 1 0 7912 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1623939100
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1623939100
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1623939100
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1623939100
transform 1 0 10304 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1623939100
transform 1 0 10120 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_87
timestamp 1623939100
transform 1 0 9108 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_95
timestamp 1623939100
transform 1 0 9844 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _723_
timestamp 1623939100
transform 1 0 10856 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1623939100
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1623939100
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1623939100
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1623939100
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_131
timestamp 1623939100
transform 1 0 13156 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1623939100
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1623939100
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1623939100
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1623939100
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1623939100
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_192
timestamp 1623939100
transform 1 0 18768 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1623939100
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_213
timestamp 1623939100
transform 1 0 20700 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_225
timestamp 1623939100
transform 1 0 21804 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_237
timestamp 1623939100
transform 1 0 22908 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_249
timestamp 1623939100
transform 1 0 24012 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1623939100
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_258
timestamp 1623939100
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_270
timestamp 1623939100
transform 1 0 25944 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_282
timestamp 1623939100
transform 1 0 27048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_294
timestamp 1623939100
transform 1 0 28152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_306
timestamp 1623939100
transform 1 0 29256 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _760_
timestamp 1623939100
transform 1 0 30452 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1623939100
transform 1 0 29992 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_315
timestamp 1623939100
transform 1 0 30084 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_338
timestamp 1623939100
transform 1 0 32200 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_350
timestamp 1623939100
transform 1 0 33304 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1623939100
transform 1 0 35236 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_362
timestamp 1623939100
transform 1 0 34408 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_370
timestamp 1623939100
transform 1 0 35144 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_372
timestamp 1623939100
transform 1 0 35328 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_384
timestamp 1623939100
transform 1 0 36432 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_396
timestamp 1623939100
transform 1 0 37536 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_408
timestamp 1623939100
transform 1 0 38640 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _707_
timestamp 1623939100
transform -1 0 42504 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1623939100
transform 1 0 40480 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1623939100
transform -1 0 40940 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_420
timestamp 1623939100
transform 1 0 39744 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_429
timestamp 1623939100
transform 1 0 40572 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_450
timestamp 1623939100
transform 1 0 42504 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_462
timestamp 1623939100
transform 1 0 43608 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_474
timestamp 1623939100
transform 1 0 44712 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1623939100
transform 1 0 45724 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_482
timestamp 1623939100
transform 1 0 45448 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_486
timestamp 1623939100
transform 1 0 45816 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_498
timestamp 1623939100
transform 1 0 46920 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_510
timestamp 1623939100
transform 1 0 48024 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_522
timestamp 1623939100
transform 1 0 49128 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_534
timestamp 1623939100
transform 1 0 50232 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1623939100
transform 1 0 50968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_543
timestamp 1623939100
transform 1 0 51060 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_555
timestamp 1623939100
transform 1 0 52164 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_567
timestamp 1623939100
transform 1 0 53268 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_579
timestamp 1623939100
transform 1 0 54372 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1623939100
transform 1 0 56212 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_591
timestamp 1623939100
transform 1 0 55476 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_600
timestamp 1623939100
transform 1 0 56304 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_612
timestamp 1623939100
transform 1 0 57408 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_624
timestamp 1623939100
transform 1 0 58512 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _456_
timestamp 1623939100
transform 1 0 59616 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_645
timestamp 1623939100
transform 1 0 60444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1623939100
transform 1 0 61456 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_653
timestamp 1623939100
transform 1 0 61180 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_657
timestamp 1623939100
transform 1 0 61548 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_669
timestamp 1623939100
transform 1 0 62652 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_681
timestamp 1623939100
transform 1 0 63756 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_693
timestamp 1623939100
transform 1 0 64860 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_705
timestamp 1623939100
transform 1 0 65964 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1623939100
transform 1 0 66700 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_714
timestamp 1623939100
transform 1 0 66792 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_726
timestamp 1623939100
transform 1 0 67896 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_738
timestamp 1623939100
transform 1 0 69000 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_750
timestamp 1623939100
transform 1 0 70104 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _347_
timestamp 1623939100
transform 1 0 70196 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1623939100
transform 1 0 71944 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_759
timestamp 1623939100
transform 1 0 70932 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_767
timestamp 1623939100
transform 1 0 71668 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_771
timestamp 1623939100
transform 1 0 72036 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_783
timestamp 1623939100
transform 1 0 73140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_795
timestamp 1623939100
transform 1 0 74244 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_807
timestamp 1623939100
transform 1 0 75348 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1623939100
transform 1 0 77188 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_819
timestamp 1623939100
transform 1 0 76452 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_828
timestamp 1623939100
transform 1 0 77280 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_840
timestamp 1623939100
transform 1 0 78384 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_852
timestamp 1623939100
transform 1 0 79488 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_864
timestamp 1623939100
transform 1 0 80592 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1623939100
transform 1 0 82432 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_876
timestamp 1623939100
transform 1 0 81696 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_885
timestamp 1623939100
transform 1 0 82524 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_897
timestamp 1623939100
transform 1 0 83628 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_909
timestamp 1623939100
transform 1 0 84732 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_921
timestamp 1623939100
transform 1 0 85836 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_933
timestamp 1623939100
transform 1 0 86940 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1623939100
transform 1 0 87676 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_942
timestamp 1623939100
transform 1 0 87768 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_954
timestamp 1623939100
transform 1 0 88872 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_966
timestamp 1623939100
transform 1 0 89976 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_978
timestamp 1623939100
transform 1 0 91080 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1623939100
transform 1 0 92920 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_990
timestamp 1623939100
transform 1 0 92184 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_999
timestamp 1623939100
transform 1 0 93012 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1011
timestamp 1623939100
transform 1 0 94116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_4  _417_
timestamp 1623939100
transform 1 0 96508 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1023
timestamp 1623939100
transform 1 0 95220 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_1035
timestamp 1623939100
transform 1 0 96324 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1623939100
transform -1 0 98808 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1623939100
transform 1 0 98164 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_1051
timestamp 1623939100
transform 1 0 97796 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_1056
timestamp 1623939100
transform 1 0 98256 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1623939100
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1623939100
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1623939100
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1623939100
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1623939100
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1623939100
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1623939100
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_58
timestamp 1623939100
transform 1 0 6440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_70
timestamp 1623939100
transform 1 0 7544 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_82
timestamp 1623939100
transform 1 0 8648 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _621_
timestamp 1623939100
transform 1 0 9476 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_323
timestamp 1623939100
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_88
timestamp 1623939100
transform 1 0 9200 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1623939100
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _560_
timestamp 1623939100
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1623939100
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1623939100
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1623939100
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_122
timestamp 1623939100
transform 1 0 12328 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_134
timestamp 1623939100
transform 1 0 13432 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_146
timestamp 1623939100
transform 1 0 14536 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_158
timestamp 1623939100
transform 1 0 15640 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _362_
timestamp 1623939100
transform 1 0 18308 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1623939100
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_170
timestamp 1623939100
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1623939100
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_184
timestamp 1623939100
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _378_
timestamp 1623939100
transform 1 0 19504 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_379
timestamp 1623939100
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1623939100
transform 1 0 19136 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1623939100
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_209
timestamp 1623939100
transform 1 0 20332 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_221
timestamp 1623939100
transform 1 0 21436 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_227
timestamp 1623939100
transform 1 0 21988 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_229
timestamp 1623939100
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_241
timestamp 1623939100
transform 1 0 23276 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_253
timestamp 1623939100
transform 1 0 24380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_265
timestamp 1623939100
transform 1 0 25484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1623939100
transform 1 0 27324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_277
timestamp 1623939100
transform 1 0 26588 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_286
timestamp 1623939100
transform 1 0 27416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_298
timestamp 1623939100
transform 1 0 28520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_310
timestamp 1623939100
transform 1 0 29624 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_322
timestamp 1623939100
transform 1 0 30728 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_8  _292_
timestamp 1623939100
transform 1 0 33028 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1623939100
transform 1 0 32568 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_334
timestamp 1623939100
transform 1 0 31832 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_343
timestamp 1623939100
transform 1 0 32660 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _477_
timestamp 1623939100
transform 1 0 35512 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_360
timestamp 1623939100
transform 1 0 34224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_372
timestamp 1623939100
transform 1 0 35328 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_383
timestamp 1623939100
transform 1 0 36340 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_395
timestamp 1623939100
transform 1 0 37444 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1623939100
transform 1 0 37812 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_400
timestamp 1623939100
transform 1 0 37904 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_412
timestamp 1623939100
transform 1 0 39008 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_424
timestamp 1623939100
transform 1 0 40112 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_436
timestamp 1623939100
transform 1 0 41216 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1623939100
transform 1 0 43056 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_448
timestamp 1623939100
transform 1 0 42320 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_457
timestamp 1623939100
transform 1 0 43148 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_469
timestamp 1623939100
transform 1 0 44252 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_481
timestamp 1623939100
transform 1 0 45356 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_493
timestamp 1623939100
transform 1 0 46460 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1623939100
transform 1 0 48300 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1623939100
transform 1 0 47564 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_514
timestamp 1623939100
transform 1 0 48392 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_526
timestamp 1623939100
transform 1 0 49496 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_538
timestamp 1623939100
transform 1 0 50600 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _679_
timestamp 1623939100
transform 1 0 52348 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_550
timestamp 1623939100
transform 1 0 51704 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_556
timestamp 1623939100
transform 1 0 52256 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_560
timestamp 1623939100
transform 1 0 52624 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1623939100
transform 1 0 53544 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_568
timestamp 1623939100
transform 1 0 53360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_571
timestamp 1623939100
transform 1 0 53636 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_583
timestamp 1623939100
transform 1 0 54740 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_595
timestamp 1623939100
transform 1 0 55844 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_607
timestamp 1623939100
transform 1 0 56948 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_619
timestamp 1623939100
transform 1 0 58052 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _352_
timestamp 1623939100
transform 1 0 60352 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1623939100
transform 1 0 58788 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_628
timestamp 1623939100
transform 1 0 58880 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_640
timestamp 1623939100
transform 1 0 59984 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_653
timestamp 1623939100
transform 1 0 61180 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_665
timestamp 1623939100
transform 1 0 62284 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1623939100
transform 1 0 64032 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_677
timestamp 1623939100
transform 1 0 63388 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_683
timestamp 1623939100
transform 1 0 63940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_685
timestamp 1623939100
transform 1 0 64124 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_697
timestamp 1623939100
transform 1 0 65228 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_709
timestamp 1623939100
transform 1 0 66332 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_721
timestamp 1623939100
transform 1 0 67436 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _766_
timestamp 1623939100
transform 1 0 70012 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1623939100
transform 1 0 69276 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_116
timestamp 1623939100
transform 1 0 69828 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_733
timestamp 1623939100
transform 1 0 68540 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_742
timestamp 1623939100
transform 1 0 69368 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_746
timestamp 1623939100
transform 1 0 69736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_768
timestamp 1623939100
transform 1 0 71760 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _381_
timestamp 1623939100
transform 1 0 72680 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_776
timestamp 1623939100
transform 1 0 72496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_787
timestamp 1623939100
transform 1 0 73508 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1623939100
transform 1 0 74520 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_795
timestamp 1623939100
transform 1 0 74244 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_799
timestamp 1623939100
transform 1 0 74612 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_811
timestamp 1623939100
transform 1 0 75716 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_823
timestamp 1623939100
transform 1 0 76820 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_835
timestamp 1623939100
transform 1 0 77924 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_847
timestamp 1623939100
transform 1 0 79028 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1623939100
transform 1 0 79764 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_856
timestamp 1623939100
transform 1 0 79856 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_868
timestamp 1623939100
transform 1 0 80960 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_880
timestamp 1623939100
transform 1 0 82064 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_892
timestamp 1623939100
transform 1 0 83168 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1623939100
transform 1 0 85008 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_904
timestamp 1623939100
transform 1 0 84272 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_913
timestamp 1623939100
transform 1 0 85100 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_925
timestamp 1623939100
transform 1 0 86204 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_937
timestamp 1623939100
transform 1 0 87308 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_949
timestamp 1623939100
transform 1 0 88412 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1623939100
transform 1 0 90252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_961
timestamp 1623939100
transform 1 0 89516 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_970
timestamp 1623939100
transform 1 0 90344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _750_
timestamp 1623939100
transform 1 0 92368 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_92
timestamp 1623939100
transform 1 0 92184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_982
timestamp 1623939100
transform 1 0 91448 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1011
timestamp 1623939100
transform 1 0 94116 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1623939100
transform 1 0 95496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_1023
timestamp 1623939100
transform 1 0 95220 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1027
timestamp 1623939100
transform 1 0 95588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1039
timestamp 1623939100
transform 1 0 96692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1623939100
transform -1 0 98808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_1051
timestamp 1623939100
transform 1 0 97796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1623939100
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1623939100
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1623939100
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1623939100
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1623939100
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1623939100
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1623939100
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1623939100
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1623939100
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1623939100
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1623939100
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1623939100
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1623939100
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1623939100
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1623939100
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1623939100
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1623939100
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1623939100
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1623939100
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _409_
timestamp 1623939100
transform -1 0 17940 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _438_
timestamp 1623939100
transform 1 0 18308 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_387
timestamp 1623939100
transform -1 0 17112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1623939100
transform 1 0 16560 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_183
timestamp 1623939100
transform 1 0 17940 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1623939100
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_196
timestamp 1623939100
transform 1 0 19136 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1623939100
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_213
timestamp 1623939100
transform 1 0 20700 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_225
timestamp 1623939100
transform 1 0 21804 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_237
timestamp 1623939100
transform 1 0 22908 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_249
timestamp 1623939100
transform 1 0 24012 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1623939100
transform 1 0 24748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_258
timestamp 1623939100
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_270
timestamp 1623939100
transform 1 0 25944 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_282
timestamp 1623939100
transform 1 0 27048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_294
timestamp 1623939100
transform 1 0 28152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_306
timestamp 1623939100
transform 1 0 29256 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1623939100
transform 1 0 29992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_315
timestamp 1623939100
transform 1 0 30084 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_327
timestamp 1623939100
transform 1 0 31188 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_339
timestamp 1623939100
transform 1 0 32292 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_351
timestamp 1623939100
transform 1 0 33396 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1623939100
transform 1 0 35236 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_363
timestamp 1623939100
transform 1 0 34500 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_372
timestamp 1623939100
transform 1 0 35328 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_384
timestamp 1623939100
transform 1 0 36432 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_396
timestamp 1623939100
transform 1 0 37536 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_408
timestamp 1623939100
transform 1 0 38640 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _411_
timestamp 1623939100
transform -1 0 41768 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1623939100
transform 1 0 40480 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_183
timestamp 1623939100
transform -1 0 41124 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_420
timestamp 1623939100
transform 1 0 39744 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_429
timestamp 1623939100
transform 1 0 40572 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_243
timestamp 1623939100
transform -1 0 41952 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_444
timestamp 1623939100
transform 1 0 41952 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_456
timestamp 1623939100
transform 1 0 43056 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_468
timestamp 1623939100
transform 1 0 44160 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1623939100
transform 1 0 45724 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_480
timestamp 1623939100
transform 1 0 45264 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_484
timestamp 1623939100
transform 1 0 45632 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_486
timestamp 1623939100
transform 1 0 45816 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_498
timestamp 1623939100
transform 1 0 46920 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _431_
timestamp 1623939100
transform 1 0 48760 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_510
timestamp 1623939100
transform 1 0 48024 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_527
timestamp 1623939100
transform 1 0 49588 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_539
timestamp 1623939100
transform 1 0 50692 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1623939100
transform 1 0 50968 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_543
timestamp 1623939100
transform 1 0 51060 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_555
timestamp 1623939100
transform 1 0 52164 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _322_
timestamp 1623939100
transform 1 0 54464 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__conb_1  _656_
timestamp 1623939100
transform 1 0 53820 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_137
timestamp 1623939100
transform 1 0 54280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_567
timestamp 1623939100
transform 1 0 53268 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_576
timestamp 1623939100
transform 1 0 54096 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1623939100
transform 1 0 56212 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_587
timestamp 1623939100
transform 1 0 55108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_600
timestamp 1623939100
transform 1 0 56304 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _323_
timestamp 1623939100
transform 1 0 58420 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_612
timestamp 1623939100
transform 1 0 57408 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_620
timestamp 1623939100
transform 1 0 58144 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_632
timestamp 1623939100
transform 1 0 59248 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_644
timestamp 1623939100
transform 1 0 60352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1623939100
transform 1 0 61456 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_657
timestamp 1623939100
transform 1 0 61548 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_669
timestamp 1623939100
transform 1 0 62652 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_681
timestamp 1623939100
transform 1 0 63756 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_693
timestamp 1623939100
transform 1 0 64860 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_705
timestamp 1623939100
transform 1 0 65964 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1623939100
transform 1 0 66700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_714
timestamp 1623939100
transform 1 0 66792 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_726
timestamp 1623939100
transform 1 0 67896 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _405_
timestamp 1623939100
transform 1 0 69000 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_747
timestamp 1623939100
transform 1 0 69828 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1623939100
transform 1 0 71944 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_759
timestamp 1623939100
transform 1 0 70932 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_767
timestamp 1623939100
transform 1 0 71668 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_771
timestamp 1623939100
transform 1 0 72036 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_783
timestamp 1623939100
transform 1 0 73140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_795
timestamp 1623939100
transform 1 0 74244 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_807
timestamp 1623939100
transform 1 0 75348 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1623939100
transform 1 0 77188 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_819
timestamp 1623939100
transform 1 0 76452 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_828
timestamp 1623939100
transform 1 0 77280 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_840
timestamp 1623939100
transform 1 0 78384 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_852
timestamp 1623939100
transform 1 0 79488 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_864
timestamp 1623939100
transform 1 0 80592 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 83444 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1623939100
transform 1 0 82432 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_876
timestamp 1623939100
transform 1 0 81696 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_885
timestamp 1623939100
transform 1 0 82524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_893
timestamp 1623939100
transform 1 0 83260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_907
timestamp 1623939100
transform 1 0 84548 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_919
timestamp 1623939100
transform 1 0 85652 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_931
timestamp 1623939100
transform 1 0 86756 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _337_
timestamp 1623939100
transform 1 0 89240 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1623939100
transform 1 0 87676 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_939
timestamp 1623939100
transform 1 0 87492 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_942
timestamp 1623939100
transform 1 0 87768 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_954
timestamp 1623939100
transform 1 0 88872 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_970
timestamp 1623939100
transform 1 0 90344 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1623939100
transform 1 0 92920 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_982
timestamp 1623939100
transform 1 0 91448 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_994
timestamp 1623939100
transform 1 0 92552 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_999
timestamp 1623939100
transform 1 0 93012 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1011
timestamp 1623939100
transform 1 0 94116 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1023
timestamp 1623939100
transform 1 0 95220 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1035
timestamp 1623939100
transform 1 0 96324 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1623939100
transform -1 0 98808 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1623939100
transform 1 0 98164 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_1047
timestamp 1623939100
transform 1 0 97428 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_1056
timestamp 1623939100
transform 1 0 98256 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1623939100
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1623939100
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1623939100
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1623939100
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1623939100
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _675_
timestamp 1623939100
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1623939100
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_266
timestamp 1623939100
transform 1 0 6624 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_51
timestamp 1623939100
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_58
timestamp 1623939100
transform 1 0 6440 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_65
timestamp 1623939100
transform 1 0 7084 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_77
timestamp 1623939100
transform 1 0 8188 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_89
timestamp 1623939100
transform 1 0 9292 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_101
timestamp 1623939100
transform 1 0 10396 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1623939100
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1623939100
transform 1 0 11500 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1623939100
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1623939100
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_139
timestamp 1623939100
transform 1 0 13892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_151
timestamp 1623939100
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_163
timestamp 1623939100
transform 1 0 16100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _319_
timestamp 1623939100
transform -1 0 18124 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1623939100
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_126
timestamp 1623939100
transform -1 0 17296 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1623939100
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_185
timestamp 1623939100
transform 1 0 18124 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_197
timestamp 1623939100
transform 1 0 19228 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1623939100
transform 1 0 22080 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_209
timestamp 1623939100
transform 1 0 20332 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_221
timestamp 1623939100
transform 1 0 21436 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_227
timestamp 1623939100
transform 1 0 21988 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_229
timestamp 1623939100
transform 1 0 22172 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_241
timestamp 1623939100
transform 1 0 23276 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _554_
timestamp 1623939100
transform 1 0 25668 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_253
timestamp 1623939100
transform 1 0 24380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_265
timestamp 1623939100
transform 1 0 25484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_270
timestamp 1623939100
transform 1 0 25944 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1623939100
transform 1 0 27324 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_282
timestamp 1623939100
transform 1 0 27048 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_286
timestamp 1623939100
transform 1 0 27416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_298
timestamp 1623939100
transform 1 0 28520 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_310
timestamp 1623939100
transform 1 0 29624 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _386_
timestamp 1623939100
transform -1 0 32200 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_228
timestamp 1623939100
transform -1 0 31556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_322
timestamp 1623939100
transform 1 0 30728 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_328
timestamp 1623939100
transform 1 0 31280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1623939100
transform 1 0 32568 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_338
timestamp 1623939100
transform 1 0 32200 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_343
timestamp 1623939100
transform 1 0 32660 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _562_
timestamp 1623939100
transform 1 0 33856 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_355
timestamp 1623939100
transform 1 0 33764 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_359
timestamp 1623939100
transform 1 0 34132 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_371
timestamp 1623939100
transform 1 0 35236 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_383
timestamp 1623939100
transform 1 0 36340 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_395
timestamp 1623939100
transform 1 0 37444 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1623939100
transform 1 0 37812 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_400
timestamp 1623939100
transform 1 0 37904 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_412
timestamp 1623939100
transform 1 0 39008 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_424
timestamp 1623939100
transform 1 0 40112 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_436
timestamp 1623939100
transform 1 0 41216 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1623939100
transform 1 0 43056 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_448
timestamp 1623939100
transform 1 0 42320 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_457
timestamp 1623939100
transform 1 0 43148 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_469
timestamp 1623939100
transform 1 0 44252 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_481
timestamp 1623939100
transform 1 0 45356 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_493
timestamp 1623939100
transform 1 0 46460 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1623939100
transform 1 0 48300 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1623939100
transform 1 0 47564 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_514
timestamp 1623939100
transform 1 0 48392 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_526
timestamp 1623939100
transform 1 0 49496 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_538
timestamp 1623939100
transform 1 0 50600 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_550
timestamp 1623939100
transform 1 0 51704 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_562
timestamp 1623939100
transform 1 0 52808 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1623939100
transform 1 0 53544 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_571
timestamp 1623939100
transform 1 0 53636 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_583
timestamp 1623939100
transform 1 0 54740 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _610_
timestamp 1623939100
transform 1 0 56120 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_595
timestamp 1623939100
transform 1 0 55844 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_601
timestamp 1623939100
transform 1 0 56396 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_613
timestamp 1623939100
transform 1 0 57500 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_625
timestamp 1623939100
transform 1 0 58604 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1623939100
transform 1 0 58788 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_628
timestamp 1623939100
transform 1 0 58880 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_640
timestamp 1623939100
transform 1 0 59984 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_652
timestamp 1623939100
transform 1 0 61088 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_664
timestamp 1623939100
transform 1 0 62192 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1623939100
transform 1 0 64032 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_676
timestamp 1623939100
transform 1 0 63296 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_685
timestamp 1623939100
transform 1 0 64124 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _629_
timestamp 1623939100
transform 1 0 65964 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_697
timestamp 1623939100
transform 1 0 65228 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_708
timestamp 1623939100
transform 1 0 66240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_720
timestamp 1623939100
transform 1 0 67344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1623939100
transform 1 0 69276 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_732
timestamp 1623939100
transform 1 0 68448 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_740
timestamp 1623939100
transform 1 0 69184 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_742
timestamp 1623939100
transform 1 0 69368 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _788_
timestamp 1623939100
transform 1 0 70840 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_25_754
timestamp 1623939100
transform 1 0 70472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_777
timestamp 1623939100
transform 1 0 72588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_789
timestamp 1623939100
transform 1 0 73692 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _770_
timestamp 1623939100
transform 1 0 75532 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1623939100
transform 1 0 74520 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_797
timestamp 1623939100
transform 1 0 74428 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_799
timestamp 1623939100
transform 1 0 74612 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_807
timestamp 1623939100
transform 1 0 75348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_828
timestamp 1623939100
transform 1 0 77280 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_840
timestamp 1623939100
transform 1 0 78384 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_852
timestamp 1623939100
transform 1 0 79488 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1623939100
transform 1 0 79764 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_856
timestamp 1623939100
transform 1 0 79856 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_868
timestamp 1623939100
transform 1 0 80960 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_880
timestamp 1623939100
transform 1 0 82064 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_892
timestamp 1623939100
transform 1 0 83168 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1623939100
transform 1 0 85008 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_904
timestamp 1623939100
transform 1 0 84272 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_913
timestamp 1623939100
transform 1 0 85100 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_925
timestamp 1623939100
transform 1 0 86204 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_937
timestamp 1623939100
transform 1 0 87308 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_949
timestamp 1623939100
transform 1 0 88412 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1623939100
transform 1 0 90252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_961
timestamp 1623939100
transform 1 0 89516 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_970
timestamp 1623939100
transform 1 0 90344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_982
timestamp 1623939100
transform 1 0 91448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_994
timestamp 1623939100
transform 1 0 92552 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1006
timestamp 1623939100
transform 1 0 93656 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_1018
timestamp 1623939100
transform 1 0 94760 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1623939100
transform 1 0 95496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1027
timestamp 1623939100
transform 1 0 95588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1039
timestamp 1623939100
transform 1 0 96692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1623939100
transform -1 0 98808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_1051
timestamp 1623939100
transform 1 0 97796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1623939100
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1623939100
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1623939100
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1623939100
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1623939100
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1623939100
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1623939100
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1623939100
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1623939100
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1623939100
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1623939100
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1623939100
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1623939100
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1623939100
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_51
timestamp 1623939100
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_58
timestamp 1623939100
transform 1 0 6440 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1623939100
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1623939100
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_70
timestamp 1623939100
transform 1 0 7544 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_82
timestamp 1623939100
transform 1 0 8648 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1623939100
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1623939100
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1623939100
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1623939100
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1623939100
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_111
timestamp 1623939100
transform 1 0 11316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1623939100
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_106
timestamp 1623939100
transform 1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_115
timestamp 1623939100
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _687_
timestamp 1623939100
transform 1 0 13616 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1623939100
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_280
timestamp 1623939100
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1623939100
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1623939100
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_127
timestamp 1623939100
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_133
timestamp 1623939100
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_139
timestamp 1623939100
transform 1 0 13892 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1623939100
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_151
timestamp 1623939100
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_163
timestamp 1623939100
transform 1 0 16100 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1623939100
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1623939100
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1623939100
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1623939100
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1623939100
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1623939100
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_192
timestamp 1623939100
transform 1 0 18768 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_201
timestamp 1623939100
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1623939100
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1623939100
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1623939100
transform 1 0 22080 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_213
timestamp 1623939100
transform 1 0 20700 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_225
timestamp 1623939100
transform 1 0 21804 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_220
timestamp 1623939100
transform 1 0 21344 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_229
timestamp 1623939100
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_237
timestamp 1623939100
transform 1 0 22908 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_249
timestamp 1623939100
transform 1 0 24012 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_241
timestamp 1623939100
transform 1 0 23276 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _734_
timestamp 1623939100
transform 1 0 25852 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1623939100
transform 1 0 24748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_258
timestamp 1623939100
transform 1 0 24840 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_266
timestamp 1623939100
transform 1 0 25576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_253
timestamp 1623939100
transform 1 0 24380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_265
timestamp 1623939100
transform 1 0 25484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1623939100
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_288
timestamp 1623939100
transform 1 0 27600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_277
timestamp 1623939100
transform 1 0 26588 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_286
timestamp 1623939100
transform 1 0 27416 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _357_
timestamp 1623939100
transform 1 0 27968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_304
timestamp 1623939100
transform 1 0 29072 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_312
timestamp 1623939100
transform 1 0 29808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_298
timestamp 1623939100
transform 1 0 28520 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_310
timestamp 1623939100
transform 1 0 29624 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1623939100
transform 1 0 29992 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_315
timestamp 1623939100
transform 1 0 30084 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_327
timestamp 1623939100
transform 1 0 31188 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1623939100
transform 1 0 30728 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1623939100
transform 1 0 32568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_339
timestamp 1623939100
transform 1 0 32292 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_351
timestamp 1623939100
transform 1 0 33396 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_334
timestamp 1623939100
transform 1 0 31832 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_343
timestamp 1623939100
transform 1 0 32660 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _466_
timestamp 1623939100
transform 1 0 34316 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1623939100
transform 1 0 35236 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_225
timestamp 1623939100
transform 1 0 34132 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_363
timestamp 1623939100
transform 1 0 34500 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_372
timestamp 1623939100
transform 1 0 35328 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_355
timestamp 1623939100
transform 1 0 33764 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_384
timestamp 1623939100
transform 1 0 36432 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_377
timestamp 1623939100
transform 1 0 35788 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_389
timestamp 1623939100
transform 1 0 36892 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1623939100
transform 1 0 37812 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_396
timestamp 1623939100
transform 1 0 37536 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_408
timestamp 1623939100
transform 1 0 38640 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_397
timestamp 1623939100
transform 1 0 37628 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_400
timestamp 1623939100
transform 1 0 37904 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_412
timestamp 1623939100
transform 1 0 39008 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _296_
timestamp 1623939100
transform 1 0 40940 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1623939100
transform 1 0 40480 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_420
timestamp 1623939100
transform 1 0 39744 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_429
timestamp 1623939100
transform 1 0 40572 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_424
timestamp 1623939100
transform 1 0 40112 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_436
timestamp 1623939100
transform 1 0 41216 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1623939100
transform 1 0 43056 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_442
timestamp 1623939100
transform 1 0 41768 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_454
timestamp 1623939100
transform 1 0 42872 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_448
timestamp 1623939100
transform 1 0 42320 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_457
timestamp 1623939100
transform 1 0 43148 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_466
timestamp 1623939100
transform 1 0 43976 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_478
timestamp 1623939100
transform 1 0 45080 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_469
timestamp 1623939100
transform 1 0 44252 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1623939100
transform 1 0 45724 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_484
timestamp 1623939100
transform 1 0 45632 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_486
timestamp 1623939100
transform 1 0 45816 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_498
timestamp 1623939100
transform 1 0 46920 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_481
timestamp 1623939100
transform 1 0 45356 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_493
timestamp 1623939100
transform 1 0 46460 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1623939100
transform 1 0 48300 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_510
timestamp 1623939100
transform 1 0 48024 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1623939100
transform 1 0 47564 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_514
timestamp 1623939100
transform 1 0 48392 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_522
timestamp 1623939100
transform 1 0 49128 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_534
timestamp 1623939100
transform 1 0 50232 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_526
timestamp 1623939100
transform 1 0 49496 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_538
timestamp 1623939100
transform 1 0 50600 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1623939100
transform 1 0 50968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_543
timestamp 1623939100
transform 1 0 51060 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_555
timestamp 1623939100
transform 1 0 52164 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_550
timestamp 1623939100
transform 1 0 51704 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_562
timestamp 1623939100
transform 1 0 52808 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1623939100
transform 1 0 53544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_567
timestamp 1623939100
transform 1 0 53268 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_579
timestamp 1623939100
transform 1 0 54372 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_571
timestamp 1623939100
transform 1 0 53636 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_583
timestamp 1623939100
transform 1 0 54740 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _320_
timestamp 1623939100
transform 1 0 56672 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1623939100
transform 1 0 56212 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_591
timestamp 1623939100
transform 1 0 55476 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_600
timestamp 1623939100
transform 1 0 56304 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_595
timestamp 1623939100
transform 1 0 55844 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1623939100
transform 1 0 57500 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_625
timestamp 1623939100
transform 1 0 58604 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_607
timestamp 1623939100
transform 1 0 56948 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_619
timestamp 1623939100
transform 1 0 58052 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1623939100
transform 1 0 58788 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_637
timestamp 1623939100
transform 1 0 59708 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_628
timestamp 1623939100
transform 1 0 58880 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_640
timestamp 1623939100
transform 1 0 59984 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1623939100
transform 1 0 61456 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_649
timestamp 1623939100
transform 1 0 60812 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_655
timestamp 1623939100
transform 1 0 61364 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_657
timestamp 1623939100
transform 1 0 61548 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_652
timestamp 1623939100
transform 1 0 61088 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_664
timestamp 1623939100
transform 1 0 62192 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1623939100
transform 1 0 64032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_669
timestamp 1623939100
transform 1 0 62652 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_681
timestamp 1623939100
transform 1 0 63756 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_676
timestamp 1623939100
transform 1 0 63296 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_685
timestamp 1623939100
transform 1 0 64124 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_693
timestamp 1623939100
transform 1 0 64860 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_705
timestamp 1623939100
transform 1 0 65964 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_697
timestamp 1623939100
transform 1 0 65228 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _720_
timestamp 1623939100
transform -1 0 69368 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1623939100
transform 1 0 66700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1623939100
transform -1 0 67804 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_714
timestamp 1623939100
transform 1 0 66792 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_722
timestamp 1623939100
transform 1 0 67528 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_709
timestamp 1623939100
transform 1 0 66332 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_721
timestamp 1623939100
transform 1 0 67436 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1623939100
transform 1 0 69276 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_742
timestamp 1623939100
transform 1 0 69368 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_733
timestamp 1623939100
transform 1 0 68540 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_742
timestamp 1623939100
transform 1 0 69368 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1623939100
transform 1 0 71944 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_754
timestamp 1623939100
transform 1 0 70472 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_766
timestamp 1623939100
transform 1 0 71576 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_754
timestamp 1623939100
transform 1 0 70472 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_766
timestamp 1623939100
transform 1 0 71576 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_771
timestamp 1623939100
transform 1 0 72036 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_783
timestamp 1623939100
transform 1 0 73140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_778
timestamp 1623939100
transform 1 0 72680 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_790
timestamp 1623939100
transform 1 0 73784 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1623939100
transform 1 0 74520 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_795
timestamp 1623939100
transform 1 0 74244 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_807
timestamp 1623939100
transform 1 0 75348 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_799
timestamp 1623939100
transform 1 0 74612 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_811
timestamp 1623939100
transform 1 0 75716 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1623939100
transform 1 0 77188 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_134
timestamp 1623939100
transform -1 0 77832 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_819
timestamp 1623939100
transform 1 0 76452 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_828
timestamp 1623939100
transform 1 0 77280 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_823
timestamp 1623939100
transform 1 0 76820 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_831
timestamp 1623939100
transform 1 0 77556 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _552_
timestamp 1623939100
transform -1 0 78660 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_386
timestamp 1623939100
transform -1 0 78844 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_840
timestamp 1623939100
transform 1 0 78384 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_852
timestamp 1623939100
transform 1 0 79488 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_845
timestamp 1623939100
transform 1 0 78844 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_853
timestamp 1623939100
transform 1 0 79580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1623939100
transform 1 0 79764 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_864
timestamp 1623939100
transform 1 0 80592 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_856
timestamp 1623939100
transform 1 0 79856 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_868
timestamp 1623939100
transform 1 0 80960 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1623939100
transform 1 0 82432 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_876
timestamp 1623939100
transform 1 0 81696 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_885
timestamp 1623939100
transform 1 0 82524 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_880
timestamp 1623939100
transform 1 0 82064 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_892
timestamp 1623939100
transform 1 0 83168 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _310_
timestamp 1623939100
transform 1 0 83996 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1623939100
transform 1 0 85008 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_897
timestamp 1623939100
transform 1 0 83628 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_910
timestamp 1623939100
transform 1 0 84824 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_904
timestamp 1623939100
transform 1 0 84272 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_913
timestamp 1623939100
transform 1 0 85100 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _611_
timestamp 1623939100
transform 1 0 87308 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_922
timestamp 1623939100
transform 1 0 85928 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_934
timestamp 1623939100
transform 1 0 87032 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_925
timestamp 1623939100
transform 1 0 86204 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1623939100
transform 1 0 87676 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_940
timestamp 1623939100
transform 1 0 87584 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_942
timestamp 1623939100
transform 1 0 87768 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_954
timestamp 1623939100
transform 1 0 88872 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_940
timestamp 1623939100
transform 1 0 87584 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_952
timestamp 1623939100
transform 1 0 88688 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1623939100
transform 1 0 90252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_966
timestamp 1623939100
transform 1 0 89976 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_978
timestamp 1623939100
transform 1 0 91080 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_964
timestamp 1623939100
transform 1 0 89792 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_968
timestamp 1623939100
transform 1 0 90160 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_970
timestamp 1623939100
transform 1 0 90344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1623939100
transform 1 0 92920 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_990
timestamp 1623939100
transform 1 0 92184 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_999
timestamp 1623939100
transform 1 0 93012 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_982
timestamp 1623939100
transform 1 0 91448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_994
timestamp 1623939100
transform 1 0 92552 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1000
timestamp 1623939100
transform 1 0 93104 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or4b_4  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 93564 0 1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__diode_2  ANTENNA_127
timestamp 1623939100
transform 1 0 93380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_128
timestamp 1623939100
transform 1 0 94576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_189
timestamp 1623939100
transform 1 0 93196 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1011
timestamp 1623939100
transform 1 0 94116 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_1018
timestamp 1623939100
transform 1 0 94760 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1623939100
transform 1 0 95496 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1023
timestamp 1623939100
transform 1 0 95220 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1035
timestamp 1623939100
transform 1 0 96324 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1027
timestamp 1623939100
transform 1 0 95588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1039
timestamp 1623939100
transform 1 0 96692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1623939100
transform -1 0 98808 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1623939100
transform -1 0 98808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1623939100
transform 1 0 98164 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_1047
timestamp 1623939100
transform 1 0 97428 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_1056
timestamp 1623939100
transform 1 0 98256 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_1051
timestamp 1623939100
transform 1 0 97796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _343_
timestamp 1623939100
transform 1 0 1840 0 -1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1623939100
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1623939100
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1623939100
transform 1 0 1748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1623939100
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_22
timestamp 1623939100
transform 1 0 3128 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_28
timestamp 1623939100
transform 1 0 3680 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1623939100
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1623939100
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_54
timestamp 1623939100
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1623939100
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_78
timestamp 1623939100
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1623939100
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1623939100
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_99
timestamp 1623939100
transform 1 0 10212 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_111
timestamp 1623939100
transform 1 0 11316 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1623939100
transform 1 0 12420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1623939100
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_135
timestamp 1623939100
transform 1 0 13524 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1623939100
transform 1 0 14352 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1623939100
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1623939100
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1623939100
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1623939100
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_192
timestamp 1623939100
transform 1 0 18768 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1623939100
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_213
timestamp 1623939100
transform 1 0 20700 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_225
timestamp 1623939100
transform 1 0 21804 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_237
timestamp 1623939100
transform 1 0 22908 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_249
timestamp 1623939100
transform 1 0 24012 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1623939100
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_258
timestamp 1623939100
transform 1 0 24840 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_270
timestamp 1623939100
transform 1 0 25944 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_282
timestamp 1623939100
transform 1 0 27048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _580_
timestamp 1623939100
transform 1 0 28152 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_297
timestamp 1623939100
transform 1 0 28428 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1623939100
transform 1 0 29532 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1623939100
transform 1 0 29992 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_313
timestamp 1623939100
transform 1 0 29900 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_315
timestamp 1623939100
transform 1 0 30084 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_327
timestamp 1623939100
transform 1 0 31188 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_339
timestamp 1623939100
transform 1 0 32292 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_351
timestamp 1623939100
transform 1 0 33396 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1623939100
transform 1 0 35236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_363
timestamp 1623939100
transform 1 0 34500 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_372
timestamp 1623939100
transform 1 0 35328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_384
timestamp 1623939100
transform 1 0 36432 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_396
timestamp 1623939100
transform 1 0 37536 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_408
timestamp 1623939100
transform 1 0 38640 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1623939100
transform 1 0 40480 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_420
timestamp 1623939100
transform 1 0 39744 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_429
timestamp 1623939100
transform 1 0 40572 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_441
timestamp 1623939100
transform 1 0 41676 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_453
timestamp 1623939100
transform 1 0 42780 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_465
timestamp 1623939100
transform 1 0 43884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_477
timestamp 1623939100
transform 1 0 44988 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1623939100
transform 1 0 45724 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_486
timestamp 1623939100
transform 1 0 45816 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_498
timestamp 1623939100
transform 1 0 46920 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_510
timestamp 1623939100
transform 1 0 48024 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_522
timestamp 1623939100
transform 1 0 49128 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_534
timestamp 1623939100
transform 1 0 50232 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1623939100
transform 1 0 50968 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_543
timestamp 1623939100
transform 1 0 51060 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_555
timestamp 1623939100
transform 1 0 52164 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_567
timestamp 1623939100
transform 1 0 53268 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_579
timestamp 1623939100
transform 1 0 54372 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1623939100
transform 1 0 56212 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_591
timestamp 1623939100
transform 1 0 55476 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_600
timestamp 1623939100
transform 1 0 56304 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _743_
timestamp 1623939100
transform -1 0 59524 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_77
timestamp 1623939100
transform -1 0 57776 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_612
timestamp 1623939100
transform 1 0 57408 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_635
timestamp 1623939100
transform 1 0 59524 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1623939100
transform 1 0 61456 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_647
timestamp 1623939100
transform 1 0 60628 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_655
timestamp 1623939100
transform 1 0 61364 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_657
timestamp 1623939100
transform 1 0 61548 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_669
timestamp 1623939100
transform 1 0 62652 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_681
timestamp 1623939100
transform 1 0 63756 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_693
timestamp 1623939100
transform 1 0 64860 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_705
timestamp 1623939100
transform 1 0 65964 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1623939100
transform 1 0 66700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_714
timestamp 1623939100
transform 1 0 66792 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_726
timestamp 1623939100
transform 1 0 67896 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_738
timestamp 1623939100
transform 1 0 69000 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_750
timestamp 1623939100
transform 1 0 70104 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1623939100
transform 1 0 71944 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_762
timestamp 1623939100
transform 1 0 71208 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_771
timestamp 1623939100
transform 1 0 72036 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_783
timestamp 1623939100
transform 1 0 73140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_795
timestamp 1623939100
transform 1 0 74244 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_807
timestamp 1623939100
transform 1 0 75348 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1623939100
transform 1 0 77188 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_819
timestamp 1623939100
transform 1 0 76452 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_828
timestamp 1623939100
transform 1 0 77280 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_840
timestamp 1623939100
transform 1 0 78384 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_852
timestamp 1623939100
transform 1 0 79488 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_864
timestamp 1623939100
transform 1 0 80592 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1623939100
transform 1 0 82432 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_876
timestamp 1623939100
transform 1 0 81696 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_885
timestamp 1623939100
transform 1 0 82524 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_897
timestamp 1623939100
transform 1 0 83628 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_909
timestamp 1623939100
transform 1 0 84732 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_921
timestamp 1623939100
transform 1 0 85836 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_933
timestamp 1623939100
transform 1 0 86940 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1623939100
transform 1 0 87676 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_942
timestamp 1623939100
transform 1 0 87768 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_954
timestamp 1623939100
transform 1 0 88872 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_966
timestamp 1623939100
transform 1 0 89976 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_978
timestamp 1623939100
transform 1 0 91080 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1623939100
transform 1 0 92920 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_990
timestamp 1623939100
transform 1 0 92184 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_999
timestamp 1623939100
transform 1 0 93012 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1011
timestamp 1623939100
transform 1 0 94116 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1023
timestamp 1623939100
transform 1 0 95220 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1035
timestamp 1623939100
transform 1 0 96324 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1623939100
transform -1 0 98808 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1623939100
transform 1 0 98164 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_1047
timestamp 1623939100
transform 1 0 97428 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_1056
timestamp 1623939100
transform 1 0 98256 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1623939100
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1623939100
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_15
timestamp 1623939100
transform 1 0 2484 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_4  _453_
timestamp 1623939100
transform -1 0 5060 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_79
timestamp 1623939100
transform -1 0 3588 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_81
timestamp 1623939100
transform -1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_83
timestamp 1623939100
transform -1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1623939100
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_80
timestamp 1623939100
transform -1 0 5244 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_82
timestamp 1623939100
transform -1 0 5428 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_84
timestamp 1623939100
transform -1 0 5612 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_49
timestamp 1623939100
transform 1 0 5612 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1623939100
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1623939100
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1623939100
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1623939100
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1623939100
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_106
timestamp 1623939100
transform 1 0 10856 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_115
timestamp 1623939100
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_127
timestamp 1623939100
transform 1 0 12788 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_139
timestamp 1623939100
transform 1 0 13892 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1623939100
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_163
timestamp 1623939100
transform 1 0 16100 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1623939100
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1623939100
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1623939100
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1623939100
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1623939100
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1623939100
transform 1 0 22080 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_220
timestamp 1623939100
transform 1 0 21344 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_229
timestamp 1623939100
transform 1 0 22172 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_241
timestamp 1623939100
transform 1 0 23276 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_253
timestamp 1623939100
transform 1 0 24380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_265
timestamp 1623939100
transform 1 0 25484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1623939100
transform 1 0 27324 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_277
timestamp 1623939100
transform 1 0 26588 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_286
timestamp 1623939100
transform 1 0 27416 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_298
timestamp 1623939100
transform 1 0 28520 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_310
timestamp 1623939100
transform 1 0 29624 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_322
timestamp 1623939100
transform 1 0 30728 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1623939100
transform 1 0 32568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_334
timestamp 1623939100
transform 1 0 31832 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_343
timestamp 1623939100
transform 1 0 32660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _793_
timestamp 1623939100
transform 1 0 33764 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_29_374
timestamp 1623939100
transform 1 0 35512 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_386
timestamp 1623939100
transform 1 0 36616 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _500_
timestamp 1623939100
transform 1 0 39284 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1623939100
transform 1 0 37812 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_167
timestamp 1623939100
transform 1 0 39100 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_398
timestamp 1623939100
transform 1 0 37720 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_400
timestamp 1623939100
transform 1 0 37904 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_412
timestamp 1623939100
transform 1 0 39008 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_424
timestamp 1623939100
transform 1 0 40112 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_436
timestamp 1623939100
transform 1 0 41216 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1623939100
transform 1 0 43056 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_448
timestamp 1623939100
transform 1 0 42320 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_457
timestamp 1623939100
transform 1 0 43148 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_469
timestamp 1623939100
transform 1 0 44252 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_481
timestamp 1623939100
transform 1 0 45356 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_493
timestamp 1623939100
transform 1 0 46460 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1623939100
transform 1 0 48300 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1623939100
transform 1 0 47564 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_514
timestamp 1623939100
transform 1 0 48392 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_526
timestamp 1623939100
transform 1 0 49496 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_538
timestamp 1623939100
transform 1 0 50600 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_550
timestamp 1623939100
transform 1 0 51704 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_562
timestamp 1623939100
transform 1 0 52808 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1623939100
transform 1 0 53544 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_571
timestamp 1623939100
transform 1 0 53636 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_583
timestamp 1623939100
transform 1 0 54740 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_595
timestamp 1623939100
transform 1 0 55844 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_607
timestamp 1623939100
transform 1 0 56948 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_619
timestamp 1623939100
transform 1 0 58052 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1623939100
transform 1 0 58788 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_628
timestamp 1623939100
transform 1 0 58880 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_640
timestamp 1623939100
transform 1 0 59984 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_652
timestamp 1623939100
transform 1 0 61088 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_664
timestamp 1623939100
transform 1 0 62192 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _366_
timestamp 1623939100
transform 1 0 62560 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1623939100
transform 1 0 64032 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_677
timestamp 1623939100
transform 1 0 63388 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_683
timestamp 1623939100
transform 1 0 63940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_685
timestamp 1623939100
transform 1 0 64124 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_697
timestamp 1623939100
transform 1 0 65228 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_709
timestamp 1623939100
transform 1 0 66332 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_721
timestamp 1623939100
transform 1 0 67436 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _704_
timestamp 1623939100
transform 1 0 69736 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1623939100
transform 1 0 69276 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_733
timestamp 1623939100
transform 1 0 68540 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_742
timestamp 1623939100
transform 1 0 69368 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_765
timestamp 1623939100
transform 1 0 71484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _541_
timestamp 1623939100
transform 1 0 73048 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_777
timestamp 1623939100
transform 1 0 72588 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_781
timestamp 1623939100
transform 1 0 72956 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_791
timestamp 1623939100
transform 1 0 73876 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _660_
timestamp 1623939100
transform 1 0 75716 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1623939100
transform 1 0 74520 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_797
timestamp 1623939100
transform 1 0 74428 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_799
timestamp 1623939100
transform 1 0 74612 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_814
timestamp 1623939100
transform 1 0 75992 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_826
timestamp 1623939100
transform 1 0 77096 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_838
timestamp 1623939100
transform 1 0 78200 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_850
timestamp 1623939100
transform 1 0 79304 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_854
timestamp 1623939100
transform 1 0 79672 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1623939100
transform 1 0 79764 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_856
timestamp 1623939100
transform 1 0 79856 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_868
timestamp 1623939100
transform 1 0 80960 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_880
timestamp 1623939100
transform 1 0 82064 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_892
timestamp 1623939100
transform 1 0 83168 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1623939100
transform 1 0 85008 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_904
timestamp 1623939100
transform 1 0 84272 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_913
timestamp 1623939100
transform 1 0 85100 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_925
timestamp 1623939100
transform 1 0 86204 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_937
timestamp 1623939100
transform 1 0 87308 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _422_
timestamp 1623939100
transform 1 0 89240 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_949
timestamp 1623939100
transform 1 0 88412 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_957
timestamp 1623939100
transform 1 0 89148 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1623939100
transform 1 0 90252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1623939100
transform -1 0 91264 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_964
timestamp 1623939100
transform 1 0 89792 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_968
timestamp 1623939100
transform 1 0 90160 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_970
timestamp 1623939100
transform 1 0 90344 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _709_
timestamp 1623939100
transform -1 0 93012 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_29_999
timestamp 1623939100
transform 1 0 93012 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1011
timestamp 1623939100
transform 1 0 94116 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1623939100
transform 1 0 95496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_1023
timestamp 1623939100
transform 1 0 95220 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1027
timestamp 1623939100
transform 1 0 95588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1039
timestamp 1623939100
transform 1 0 96692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1623939100
transform -1 0 98808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_1051
timestamp 1623939100
transform 1 0 97796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1623939100
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1623939100
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1623939100
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1623939100
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_113
timestamp 1623939100
transform -1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1623939100
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_30
timestamp 1623939100
transform 1 0 3864 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_38
timestamp 1623939100
transform 1 0 4600 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _763_
timestamp 1623939100
transform -1 0 6992 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_111
timestamp 1623939100
transform -1 0 5244 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_112
timestamp 1623939100
transform -1 0 7176 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_114
timestamp 1623939100
transform -1 0 7360 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1623939100
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_80
timestamp 1623939100
transform 1 0 8464 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1623939100
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1623939100
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_99
timestamp 1623939100
transform 1 0 10212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_111
timestamp 1623939100
transform 1 0 11316 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_123
timestamp 1623939100
transform 1 0 12420 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1623939100
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_135
timestamp 1623939100
transform 1 0 13524 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1623939100
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _722_
timestamp 1623939100
transform 1 0 15548 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_30_156
timestamp 1623939100
transform 1 0 15456 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_176
timestamp 1623939100
transform 1 0 17296 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1623939100
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_188
timestamp 1623939100
transform 1 0 18400 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1623939100
transform 1 0 19596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_213
timestamp 1623939100
transform 1 0 20700 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_225
timestamp 1623939100
transform 1 0 21804 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_237
timestamp 1623939100
transform 1 0 22908 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_249
timestamp 1623939100
transform 1 0 24012 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1623939100
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_258
timestamp 1623939100
transform 1 0 24840 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_270
timestamp 1623939100
transform 1 0 25944 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_282
timestamp 1623939100
transform 1 0 27048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_294
timestamp 1623939100
transform 1 0 28152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_306
timestamp 1623939100
transform 1 0 29256 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1623939100
transform 1 0 29992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_315
timestamp 1623939100
transform 1 0 30084 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_327
timestamp 1623939100
transform 1 0 31188 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_339
timestamp 1623939100
transform 1 0 32292 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_351
timestamp 1623939100
transform 1 0 33396 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1623939100
transform 1 0 35236 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_363
timestamp 1623939100
transform 1 0 34500 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_372
timestamp 1623939100
transform 1 0 35328 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_384
timestamp 1623939100
transform 1 0 36432 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_396
timestamp 1623939100
transform 1 0 37536 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_408
timestamp 1623939100
transform 1 0 38640 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1623939100
transform 1 0 40480 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_420
timestamp 1623939100
transform 1 0 39744 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_429
timestamp 1623939100
transform 1 0 40572 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_441
timestamp 1623939100
transform 1 0 41676 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_453
timestamp 1623939100
transform 1 0 42780 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_465
timestamp 1623939100
transform 1 0 43884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_477
timestamp 1623939100
transform 1 0 44988 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1623939100
transform 1 0 45724 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_486
timestamp 1623939100
transform 1 0 45816 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_498
timestamp 1623939100
transform 1 0 46920 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_510
timestamp 1623939100
transform 1 0 48024 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_522
timestamp 1623939100
transform 1 0 49128 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_534
timestamp 1623939100
transform 1 0 50232 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _513_
timestamp 1623939100
transform -1 0 53176 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1623939100
transform 1 0 50968 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_169
timestamp 1623939100
transform -1 0 52348 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_543
timestamp 1623939100
transform 1 0 51060 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_566
timestamp 1623939100
transform 1 0 53176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_578
timestamp 1623939100
transform 1 0 54280 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1623939100
transform 1 0 56212 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_590
timestamp 1623939100
transform 1 0 55384 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_598
timestamp 1623939100
transform 1 0 56120 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_600
timestamp 1623939100
transform 1 0 56304 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_612
timestamp 1623939100
transform 1 0 57408 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_624
timestamp 1623939100
transform 1 0 58512 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__inv_4  _286_
timestamp 1623939100
transform 1 0 59248 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_30_637
timestamp 1623939100
transform 1 0 59708 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1623939100
transform 1 0 61456 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_649
timestamp 1623939100
transform 1 0 60812 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_655
timestamp 1623939100
transform 1 0 61364 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_657
timestamp 1623939100
transform 1 0 61548 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_669
timestamp 1623939100
transform 1 0 62652 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_681
timestamp 1623939100
transform 1 0 63756 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_693
timestamp 1623939100
transform 1 0 64860 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_705
timestamp 1623939100
transform 1 0 65964 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1623939100
transform 1 0 66700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_714
timestamp 1623939100
transform 1 0 66792 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_726
timestamp 1623939100
transform 1 0 67896 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_738
timestamp 1623939100
transform 1 0 69000 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_750
timestamp 1623939100
transform 1 0 70104 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _387_
timestamp 1623939100
transform 1 0 70748 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1623939100
transform 1 0 71944 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_756
timestamp 1623939100
transform 1 0 70656 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_763
timestamp 1623939100
transform 1 0 71300 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_769
timestamp 1623939100
transform 1 0 71852 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_771
timestamp 1623939100
transform 1 0 72036 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_783
timestamp 1623939100
transform 1 0 73140 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _617_
timestamp 1623939100
transform 1 0 74428 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_795
timestamp 1623939100
transform 1 0 74244 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_800
timestamp 1623939100
transform 1 0 74704 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_812
timestamp 1623939100
transform 1 0 75808 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1623939100
transform 1 0 77188 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_824
timestamp 1623939100
transform 1 0 76912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_828
timestamp 1623939100
transform 1 0 77280 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_840
timestamp 1623939100
transform 1 0 78384 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_852
timestamp 1623939100
transform 1 0 79488 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_864
timestamp 1623939100
transform 1 0 80592 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1623939100
transform 1 0 82432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_876
timestamp 1623939100
transform 1 0 81696 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_885
timestamp 1623939100
transform 1 0 82524 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_897
timestamp 1623939100
transform 1 0 83628 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_909
timestamp 1623939100
transform 1 0 84732 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_921
timestamp 1623939100
transform 1 0 85836 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_933
timestamp 1623939100
transform 1 0 86940 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1623939100
transform 1 0 87676 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_942
timestamp 1623939100
transform 1 0 87768 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_954
timestamp 1623939100
transform 1 0 88872 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_966
timestamp 1623939100
transform 1 0 89976 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_978
timestamp 1623939100
transform 1 0 91080 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1623939100
transform 1 0 92920 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_990
timestamp 1623939100
transform 1 0 92184 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_999
timestamp 1623939100
transform 1 0 93012 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1011
timestamp 1623939100
transform 1 0 94116 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1023
timestamp 1623939100
transform 1 0 95220 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1035
timestamp 1623939100
transform 1 0 96324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1623939100
transform -1 0 98808 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1623939100
transform 1 0 98164 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_1047
timestamp 1623939100
transform 1 0 97428 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_1056
timestamp 1623939100
transform 1 0 98256 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1623939100
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1623939100
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1623939100
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1623939100
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1623939100
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1623939100
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_51
timestamp 1623939100
transform 1 0 5796 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_58
timestamp 1623939100
transform 1 0 6440 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_70
timestamp 1623939100
transform 1 0 7544 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_82
timestamp 1623939100
transform 1 0 8648 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1623939100
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1623939100
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_106
timestamp 1623939100
transform 1 0 10856 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1623939100
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1623939100
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1623939100
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1623939100
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_163
timestamp 1623939100
transform 1 0 16100 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1623939100
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1623939100
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1623939100
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1623939100
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1623939100
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1623939100
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_220
timestamp 1623939100
transform 1 0 21344 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1623939100
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_241
timestamp 1623939100
transform 1 0 23276 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_253
timestamp 1623939100
transform 1 0 24380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_265
timestamp 1623939100
transform 1 0 25484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1623939100
transform 1 0 27324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_277
timestamp 1623939100
transform 1 0 26588 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1623939100
transform 1 0 27416 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_298
timestamp 1623939100
transform 1 0 28520 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_310
timestamp 1623939100
transform 1 0 29624 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_322
timestamp 1623939100
transform 1 0 30728 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1623939100
transform 1 0 32568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_334
timestamp 1623939100
transform 1 0 31832 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_343
timestamp 1623939100
transform 1 0 32660 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_355
timestamp 1623939100
transform 1 0 33764 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_367
timestamp 1623939100
transform 1 0 34868 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_375
timestamp 1623939100
transform 1 0 35604 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _468_
timestamp 1623939100
transform 1 0 35880 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_31_387
timestamp 1623939100
transform 1 0 36708 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1623939100
transform 1 0 37812 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_400
timestamp 1623939100
transform 1 0 37904 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_412
timestamp 1623939100
transform 1 0 39008 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_424
timestamp 1623939100
transform 1 0 40112 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_436
timestamp 1623939100
transform 1 0 41216 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1623939100
transform 1 0 43056 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_448
timestamp 1623939100
transform 1 0 42320 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_457
timestamp 1623939100
transform 1 0 43148 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _787_
timestamp 1623939100
transform -1 0 46184 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_124
timestamp 1623939100
transform -1 0 44436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_490
timestamp 1623939100
transform 1 0 46184 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1623939100
transform 1 0 48300 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_502
timestamp 1623939100
transform 1 0 47288 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_510
timestamp 1623939100
transform 1 0 48024 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_514
timestamp 1623939100
transform 1 0 48392 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _308_
timestamp 1623939100
transform 1 0 50232 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _631_
timestamp 1623939100
transform 1 0 49128 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_135
timestamp 1623939100
transform 1 0 50048 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_525
timestamp 1623939100
transform 1 0 49404 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_531
timestamp 1623939100
transform 1 0 49956 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  _471_
timestamp 1623939100
transform 1 0 52348 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_543
timestamp 1623939100
transform 1 0 51060 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_555
timestamp 1623939100
transform 1 0 52164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1623939100
transform 1 0 53544 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_563
timestamp 1623939100
transform 1 0 52900 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_569
timestamp 1623939100
transform 1 0 53452 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_571
timestamp 1623939100
transform 1 0 53636 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_583
timestamp 1623939100
transform 1 0 54740 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_595
timestamp 1623939100
transform 1 0 55844 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_607
timestamp 1623939100
transform 1 0 56948 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_619
timestamp 1623939100
transform 1 0 58052 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _517_
timestamp 1623939100
transform 1 0 60352 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1623939100
transform 1 0 58788 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_628
timestamp 1623939100
transform 1 0 58880 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_640
timestamp 1623939100
transform 1 0 59984 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_653
timestamp 1623939100
transform 1 0 61180 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_665
timestamp 1623939100
transform 1 0 62284 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1623939100
transform 1 0 64032 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_677
timestamp 1623939100
transform 1 0 63388 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_683
timestamp 1623939100
transform 1 0 63940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_685
timestamp 1623939100
transform 1 0 64124 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_697
timestamp 1623939100
transform 1 0 65228 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_709
timestamp 1623939100
transform 1 0 66332 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_721
timestamp 1623939100
transform 1 0 67436 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1623939100
transform 1 0 69276 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_733
timestamp 1623939100
transform 1 0 68540 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_742
timestamp 1623939100
transform 1 0 69368 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_754
timestamp 1623939100
transform 1 0 70472 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_766
timestamp 1623939100
transform 1 0 71576 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_778
timestamp 1623939100
transform 1 0 72680 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_790
timestamp 1623939100
transform 1 0 73784 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1623939100
transform 1 0 74520 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_799
timestamp 1623939100
transform 1 0 74612 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_811
timestamp 1623939100
transform 1 0 75716 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_823
timestamp 1623939100
transform 1 0 76820 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_835
timestamp 1623939100
transform 1 0 77924 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_847
timestamp 1623939100
transform 1 0 79028 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1623939100
transform 1 0 79764 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_856
timestamp 1623939100
transform 1 0 79856 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_868
timestamp 1623939100
transform 1 0 80960 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_880
timestamp 1623939100
transform 1 0 82064 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_892
timestamp 1623939100
transform 1 0 83168 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1623939100
transform 1 0 85008 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_904
timestamp 1623939100
transform 1 0 84272 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_913
timestamp 1623939100
transform 1 0 85100 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_925
timestamp 1623939100
transform 1 0 86204 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_937
timestamp 1623939100
transform 1 0 87308 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_949
timestamp 1623939100
transform 1 0 88412 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1623939100
transform 1 0 90252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_961
timestamp 1623939100
transform 1 0 89516 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_970
timestamp 1623939100
transform 1 0 90344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_982
timestamp 1623939100
transform 1 0 91448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_994
timestamp 1623939100
transform 1 0 92552 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1006
timestamp 1623939100
transform 1 0 93656 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_1018
timestamp 1623939100
transform 1 0 94760 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1623939100
transform 1 0 95496 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1027
timestamp 1623939100
transform 1 0 95588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1039
timestamp 1623939100
transform 1 0 96692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _667_
timestamp 1623939100
transform 1 0 97888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1623939100
transform -1 0 98808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1051
timestamp 1623939100
transform 1 0 97796 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_1055
timestamp 1623939100
transform 1 0 98164 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1623939100
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input295
timestamp 1623939100
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_6
timestamp 1623939100
transform 1 0 1656 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_18
timestamp 1623939100
transform 1 0 2760 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1623939100
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_26
timestamp 1623939100
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_30
timestamp 1623939100
transform 1 0 3864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_42
timestamp 1623939100
transform 1 0 4968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_54
timestamp 1623939100
transform 1 0 6072 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_66
timestamp 1623939100
transform 1 0 7176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_78
timestamp 1623939100
transform 1 0 8280 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1623939100
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1623939100
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_99
timestamp 1623939100
transform 1 0 10212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_111
timestamp 1623939100
transform 1 0 11316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1623939100
transform 1 0 12420 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1623939100
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_135
timestamp 1623939100
transform 1 0 13524 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_144
timestamp 1623939100
transform 1 0 14352 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1623939100
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1623939100
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_180
timestamp 1623939100
transform 1 0 17664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1623939100
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_192
timestamp 1623939100
transform 1 0 18768 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1623939100
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_213
timestamp 1623939100
transform 1 0 20700 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_225
timestamp 1623939100
transform 1 0 21804 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_237
timestamp 1623939100
transform 1 0 22908 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_249
timestamp 1623939100
transform 1 0 24012 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1623939100
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_258
timestamp 1623939100
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_270
timestamp 1623939100
transform 1 0 25944 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_282
timestamp 1623939100
transform 1 0 27048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _510_
timestamp 1623939100
transform 1 0 28704 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_32_294
timestamp 1623939100
transform 1 0 28152 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_309
timestamp 1623939100
transform 1 0 29532 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1623939100
transform 1 0 29992 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_313
timestamp 1623939100
transform 1 0 29900 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_315
timestamp 1623939100
transform 1 0 30084 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_327
timestamp 1623939100
transform 1 0 31188 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_1_wb_clk_i
timestamp 1623939100
transform 1 0 33212 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_339
timestamp 1623939100
transform 1 0 32292 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_347
timestamp 1623939100
transform 1 0 33028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_352
timestamp 1623939100
transform 1 0 33488 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1623939100
transform 1 0 35236 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_364
timestamp 1623939100
transform 1 0 34592 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_370
timestamp 1623939100
transform 1 0 35144 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_372
timestamp 1623939100
transform 1 0 35328 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_384
timestamp 1623939100
transform 1 0 36432 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i
timestamp 1623939100
transform 1 0 38456 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_396
timestamp 1623939100
transform 1 0 37536 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_404
timestamp 1623939100
transform 1 0 38272 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_409
timestamp 1623939100
transform 1 0 38732 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1623939100
transform 1 0 40480 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_421
timestamp 1623939100
transform 1 0 39836 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_427
timestamp 1623939100
transform 1 0 40388 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_429
timestamp 1623939100
transform 1 0 40572 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_441
timestamp 1623939100
transform 1 0 41676 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_453
timestamp 1623939100
transform 1 0 42780 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_465
timestamp 1623939100
transform 1 0 43884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_477
timestamp 1623939100
transform 1 0 44988 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1623939100
transform 1 0 45724 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_486
timestamp 1623939100
transform 1 0 45816 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_498
timestamp 1623939100
transform 1 0 46920 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 48760 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_32_510
timestamp 1623939100
transform 1 0 48024 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_538
timestamp 1623939100
transform 1 0 50600 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1623939100
transform 1 0 50968 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_543
timestamp 1623939100
transform 1 0 51060 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_555
timestamp 1623939100
transform 1 0 52164 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _313_
timestamp 1623939100
transform 1 0 54648 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_32_567
timestamp 1623939100
transform 1 0 53268 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_579
timestamp 1623939100
transform 1 0 54372 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1623939100
transform 1 0 56212 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_589
timestamp 1623939100
transform 1 0 55292 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_597
timestamp 1623939100
transform 1 0 56028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_600
timestamp 1623939100
transform 1 0 56304 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_612
timestamp 1623939100
transform 1 0 57408 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_624
timestamp 1623939100
transform 1 0 58512 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1623939100
transform 1 0 59248 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_635
timestamp 1623939100
transform 1 0 59524 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1623939100
transform 1 0 61456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_647
timestamp 1623939100
transform 1 0 60628 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_655
timestamp 1623939100
transform 1 0 61364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_657
timestamp 1623939100
transform 1 0 61548 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_669
timestamp 1623939100
transform 1 0 62652 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_681
timestamp 1623939100
transform 1 0 63756 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_687
timestamp 1623939100
transform 1 0 64308 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_1_wb_clk_i
timestamp 1623939100
transform 1 0 64400 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_691
timestamp 1623939100
transform 1 0 64676 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_703
timestamp 1623939100
transform 1 0 65780 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1623939100
transform 1 0 66700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_711
timestamp 1623939100
transform 1 0 66516 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_714
timestamp 1623939100
transform 1 0 66792 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_726
timestamp 1623939100
transform 1 0 67896 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_738
timestamp 1623939100
transform 1 0 69000 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_750
timestamp 1623939100
transform 1 0 70104 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1623939100
transform 1 0 71944 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_762
timestamp 1623939100
transform 1 0 71208 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_771
timestamp 1623939100
transform 1 0 72036 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_783
timestamp 1623939100
transform 1 0 73140 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_791
timestamp 1623939100
transform 1 0 73876 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _284_
timestamp 1623939100
transform 1 0 75624 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_8  _485_
timestamp 1623939100
transform 1 0 73968 0 -1 20128
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_32_803
timestamp 1623939100
transform 1 0 74980 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_809
timestamp 1623939100
transform 1 0 75532 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1623939100
transform 1 0 77188 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_817
timestamp 1623939100
transform 1 0 76268 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_825
timestamp 1623939100
transform 1 0 77004 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_828
timestamp 1623939100
transform 1 0 77280 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_840
timestamp 1623939100
transform 1 0 78384 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_852
timestamp 1623939100
transform 1 0 79488 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_864
timestamp 1623939100
transform 1 0 80592 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1623939100
transform 1 0 82432 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_876
timestamp 1623939100
transform 1 0 81696 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_885
timestamp 1623939100
transform 1 0 82524 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_897
timestamp 1623939100
transform 1 0 83628 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_909
timestamp 1623939100
transform 1 0 84732 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_921
timestamp 1623939100
transform 1 0 85836 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_933
timestamp 1623939100
transform 1 0 86940 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1623939100
transform 1 0 87676 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_942
timestamp 1623939100
transform 1 0 87768 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_954
timestamp 1623939100
transform 1 0 88872 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_966
timestamp 1623939100
transform 1 0 89976 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_978
timestamp 1623939100
transform 1 0 91080 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1623939100
transform 1 0 92920 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_990
timestamp 1623939100
transform 1 0 92184 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_999
timestamp 1623939100
transform 1 0 93012 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1011
timestamp 1623939100
transform 1 0 94116 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1023
timestamp 1623939100
transform 1 0 95220 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_1035
timestamp 1623939100
transform 1 0 96324 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1623939100
transform -1 0 98808 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1623939100
transform 1 0 98164 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output446
timestamp 1623939100
transform 1 0 97428 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_251
timestamp 1623939100
transform 1 0 97244 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_1043
timestamp 1623939100
transform 1 0 97060 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_1051
timestamp 1623939100
transform 1 0 97796 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_1056
timestamp 1623939100
transform 1 0 98256 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _444_
timestamp 1623939100
transform -1 0 2576 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1623939100
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1623939100
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_156
timestamp 1623939100
transform -1 0 1748 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_157
timestamp 1623939100
transform -1 0 2760 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_206
timestamp 1623939100
transform -1 0 1564 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1623939100
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1623939100
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_18
timestamp 1623939100
transform 1 0 2760 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1623939100
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_172
timestamp 1623939100
transform -1 0 5060 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1623939100
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1623939100
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_26
timestamp 1623939100
transform 1 0 3496 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_30
timestamp 1623939100
transform 1 0 3864 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_38
timestamp 1623939100
transform 1 0 4600 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _522_
timestamp 1623939100
transform -1 0 6072 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1623939100
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_170
timestamp 1623939100
transform -1 0 5244 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_171
timestamp 1623939100
transform -1 0 6256 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_51
timestamp 1623939100
transform 1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_58
timestamp 1623939100
transform 1 0 6440 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1623939100
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_70
timestamp 1623939100
transform 1 0 7544 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_82
timestamp 1623939100
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1623939100
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_80
timestamp 1623939100
transform 1 0 8464 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1623939100
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1623939100
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1623939100
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1623939100
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1623939100
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_106
timestamp 1623939100
transform 1 0 10856 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1623939100
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_111
timestamp 1623939100
transform 1 0 11316 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1623939100
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1623939100
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1623939100
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1623939100
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_135
timestamp 1623939100
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_144
timestamp 1623939100
transform 1 0 14352 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _683_
timestamp 1623939100
transform 1 0 15456 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _716_
timestamp 1623939100
transform 1 0 15916 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_33_151
timestamp 1623939100
transform 1 0 14996 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1623939100
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1623939100
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_156
timestamp 1623939100
transform 1 0 15456 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_160
timestamp 1623939100
transform 1 0 15824 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1623939100
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1623939100
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1623939100
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_180
timestamp 1623939100
transform 1 0 17664 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _359_
timestamp 1623939100
transform 1 0 18584 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1623939100
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1623939100
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1623939100
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_188
timestamp 1623939100
transform 1 0 18400 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_196
timestamp 1623939100
transform 1 0 19136 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1623939100
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1623939100
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_220
timestamp 1623939100
transform 1 0 21344 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_229
timestamp 1623939100
transform 1 0 22172 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_213
timestamp 1623939100
transform 1 0 20700 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_225
timestamp 1623939100
transform 1 0 21804 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _625_
timestamp 1623939100
transform 1 0 22540 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_236
timestamp 1623939100
transform 1 0 22816 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_248
timestamp 1623939100
transform 1 0 23920 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_237
timestamp 1623939100
transform 1 0 22908 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_249
timestamp 1623939100
transform 1 0 24012 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1623939100
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_260
timestamp 1623939100
transform 1 0 25024 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1623939100
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_270
timestamp 1623939100
transform 1 0 25944 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1623939100
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_272
timestamp 1623939100
transform 1 0 26128 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_284
timestamp 1623939100
transform 1 0 27232 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_286
timestamp 1623939100
transform 1 0 27416 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_282
timestamp 1623939100
transform 1 0 27048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_298
timestamp 1623939100
transform 1 0 28520 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_310
timestamp 1623939100
transform 1 0 29624 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_294
timestamp 1623939100
transform 1 0 28152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_306
timestamp 1623939100
transform 1 0 29256 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1623939100
transform 1 0 29992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_322
timestamp 1623939100
transform 1 0 30728 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_315
timestamp 1623939100
transform 1 0 30084 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_327
timestamp 1623939100
transform 1 0 31188 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1623939100
transform 1 0 32568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_334
timestamp 1623939100
transform 1 0 31832 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1623939100
transform 1 0 32660 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_339
timestamp 1623939100
transform 1 0 32292 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_351
timestamp 1623939100
transform 1 0 33396 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _681_
timestamp 1623939100
transform 1 0 34040 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1623939100
transform 1 0 35236 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_355
timestamp 1623939100
transform 1 0 33764 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1623939100
transform 1 0 34316 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1623939100
transform 1 0 35420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_363
timestamp 1623939100
transform 1 0 34500 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_372
timestamp 1623939100
transform 1 0 35328 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_385
timestamp 1623939100
transform 1 0 36524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_384
timestamp 1623939100
transform 1 0 36432 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1623939100
transform 1 0 37812 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_397
timestamp 1623939100
transform 1 0 37628 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_400
timestamp 1623939100
transform 1 0 37904 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_412
timestamp 1623939100
transform 1 0 39008 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_396
timestamp 1623939100
transform 1 0 37536 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_408
timestamp 1623939100
transform 1 0 38640 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1623939100
transform 1 0 40480 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_424
timestamp 1623939100
transform 1 0 40112 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_436
timestamp 1623939100
transform 1 0 41216 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_420
timestamp 1623939100
transform 1 0 39744 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_429
timestamp 1623939100
transform 1 0 40572 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1623939100
transform 1 0 43056 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_448
timestamp 1623939100
transform 1 0 42320 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_457
timestamp 1623939100
transform 1 0 43148 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_441
timestamp 1623939100
transform 1 0 41676 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_453
timestamp 1623939100
transform 1 0 42780 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _493_
timestamp 1623939100
transform 1 0 44160 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_33_469
timestamp 1623939100
transform 1 0 44252 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_465
timestamp 1623939100
transform 1 0 43884 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_477
timestamp 1623939100
transform 1 0 44988 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1623939100
transform 1 0 45724 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_481
timestamp 1623939100
transform 1 0 45356 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_493
timestamp 1623939100
transform 1 0 46460 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_486
timestamp 1623939100
transform 1 0 45816 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_498
timestamp 1623939100
transform 1 0 46920 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1623939100
transform 1 0 48300 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1623939100
transform 1 0 47564 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_514
timestamp 1623939100
transform 1 0 48392 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_510
timestamp 1623939100
transform 1 0 48024 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_526
timestamp 1623939100
transform 1 0 49496 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_538
timestamp 1623939100
transform 1 0 50600 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_522
timestamp 1623939100
transform 1 0 49128 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_534
timestamp 1623939100
transform 1 0 50232 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _484_
timestamp 1623939100
transform 1 0 51980 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1623939100
transform 1 0 50968 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_550
timestamp 1623939100
transform 1 0 51704 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_559
timestamp 1623939100
transform 1 0 52532 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_543
timestamp 1623939100
transform 1 0 51060 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_555
timestamp 1623939100
transform 1 0 52164 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1623939100
transform 1 0 53544 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_567
timestamp 1623939100
transform 1 0 53268 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_571
timestamp 1623939100
transform 1 0 53636 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_583
timestamp 1623939100
transform 1 0 54740 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_567
timestamp 1623939100
transform 1 0 53268 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_579
timestamp 1623939100
transform 1 0 54372 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1623939100
transform 1 0 56212 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_595
timestamp 1623939100
transform 1 0 55844 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_591
timestamp 1623939100
transform 1 0 55476 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_600
timestamp 1623939100
transform 1 0 56304 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_607
timestamp 1623939100
transform 1 0 56948 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_619
timestamp 1623939100
transform 1 0 58052 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_612
timestamp 1623939100
transform 1 0 57408 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_624
timestamp 1623939100
transform 1 0 58512 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1623939100
transform 1 0 58788 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_628
timestamp 1623939100
transform 1 0 58880 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_640
timestamp 1623939100
transform 1 0 59984 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_636
timestamp 1623939100
transform 1 0 59616 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1623939100
transform 1 0 61456 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_652
timestamp 1623939100
transform 1 0 61088 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_664
timestamp 1623939100
transform 1 0 62192 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_648
timestamp 1623939100
transform 1 0 60720 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_657
timestamp 1623939100
transform 1 0 61548 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _353_
timestamp 1623939100
transform 1 0 63020 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _624_
timestamp 1623939100
transform 1 0 63940 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1623939100
transform 1 0 64032 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_676
timestamp 1623939100
transform 1 0 63296 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_685
timestamp 1623939100
transform 1 0 64124 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_669
timestamp 1623939100
transform 1 0 62652 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_679
timestamp 1623939100
transform 1 0 63572 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_686
timestamp 1623939100
transform 1 0 64216 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _719_
timestamp 1623939100
transform 1 0 64492 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_33_706
timestamp 1623939100
transform 1 0 66056 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_698
timestamp 1623939100
transform 1 0 65320 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _614_
timestamp 1623939100
transform 1 0 67160 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1623939100
transform 1 0 66700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_718
timestamp 1623939100
transform 1 0 67160 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_710
timestamp 1623939100
transform 1 0 66424 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_714
timestamp 1623939100
transform 1 0 66792 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_721
timestamp 1623939100
transform 1 0 67436 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _439_
timestamp 1623939100
transform 1 0 69828 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1623939100
transform 1 0 69276 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_730
timestamp 1623939100
transform 1 0 68264 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_738
timestamp 1623939100
transform 1 0 69000 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_742
timestamp 1623939100
transform 1 0 69368 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_746
timestamp 1623939100
transform 1 0 69736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_733
timestamp 1623939100
transform 1 0 68540 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_745
timestamp 1623939100
transform 1 0 69644 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _335_
timestamp 1623939100
transform -1 0 72956 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1623939100
transform 1 0 71944 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_119
timestamp 1623939100
transform -1 0 71484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_756
timestamp 1623939100
transform 1 0 70656 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_762
timestamp 1623939100
transform 1 0 71208 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_757
timestamp 1623939100
transform 1 0 70748 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_769
timestamp 1623939100
transform 1 0 71852 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_120
timestamp 1623939100
transform -1 0 73140 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_783
timestamp 1623939100
transform 1 0 73140 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_771
timestamp 1623939100
transform 1 0 72036 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_783
timestamp 1623939100
transform 1 0 73140 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1623939100
transform 1 0 74520 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_795
timestamp 1623939100
transform 1 0 74244 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_799
timestamp 1623939100
transform 1 0 74612 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_811
timestamp 1623939100
transform 1 0 75716 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_795
timestamp 1623939100
transform 1 0 74244 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_807
timestamp 1623939100
transform 1 0 75348 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1623939100
transform 1 0 77188 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_823
timestamp 1623939100
transform 1 0 76820 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_819
timestamp 1623939100
transform 1 0 76452 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_828
timestamp 1623939100
transform 1 0 77280 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_835
timestamp 1623939100
transform 1 0 77924 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_847
timestamp 1623939100
transform 1 0 79028 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_840
timestamp 1623939100
transform 1 0 78384 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_852
timestamp 1623939100
transform 1 0 79488 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _473_
timestamp 1623939100
transform -1 0 82432 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _710_
timestamp 1623939100
transform 1 0 80040 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1623939100
transform 1 0 79764 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_165
timestamp 1623939100
transform -1 0 81604 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_856
timestamp 1623939100
transform 1 0 79856 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_868
timestamp 1623939100
transform 1 0 80960 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_872
timestamp 1623939100
transform 1 0 81328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1623939100
transform 1 0 82432 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_884
timestamp 1623939100
transform 1 0 82432 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_877
timestamp 1623939100
transform 1 0 81788 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_883
timestamp 1623939100
transform 1 0 82340 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_885
timestamp 1623939100
transform 1 0 82524 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1623939100
transform 1 0 85008 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_896
timestamp 1623939100
transform 1 0 83536 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_908
timestamp 1623939100
transform 1 0 84640 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_913
timestamp 1623939100
transform 1 0 85100 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_897
timestamp 1623939100
transform 1 0 83628 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_909
timestamp 1623939100
transform 1 0 84732 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_925
timestamp 1623939100
transform 1 0 86204 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_937
timestamp 1623939100
transform 1 0 87308 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_921
timestamp 1623939100
transform 1 0 85836 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_933
timestamp 1623939100
transform 1 0 86940 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1623939100
transform 1 0 87676 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_949
timestamp 1623939100
transform 1 0 88412 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_942
timestamp 1623939100
transform 1 0 87768 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_954
timestamp 1623939100
transform 1 0 88872 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1623939100
transform 1 0 90252 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_961
timestamp 1623939100
transform 1 0 89516 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_970
timestamp 1623939100
transform 1 0 90344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_966
timestamp 1623939100
transform 1 0 89976 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_978
timestamp 1623939100
transform 1 0 91080 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1623939100
transform 1 0 92920 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_72
timestamp 1623939100
transform 1 0 93104 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_75
timestamp 1623939100
transform 1 0 92736 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_982
timestamp 1623939100
transform 1 0 91448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_994
timestamp 1623939100
transform 1 0 92552 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_990
timestamp 1623939100
transform 1 0 92184 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_999
timestamp 1623939100
transform 1 0 93012 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _435_
timestamp 1623939100
transform 1 0 93472 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _742_
timestamp 1623939100
transform 1 0 93656 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_68
timestamp 1623939100
transform 1 0 93472 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_70
timestamp 1623939100
transform 1 0 93288 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_1002
timestamp 1623939100
transform 1 0 93288 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1013
timestamp 1623939100
transform 1 0 94300 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1025
timestamp 1623939100
transform 1 0 95404 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_74
timestamp 1623939100
transform 1 0 95956 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_73
timestamp 1623939100
transform 1 0 95772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_71
timestamp 1623939100
transform 1 0 95588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_69
timestamp 1623939100
transform 1 0 95404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1623939100
transform 1 0 95496 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_1039
timestamp 1623939100
transform 1 0 96692 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_76
timestamp 1623939100
transform 1 0 96140 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1035
timestamp 1623939100
transform 1 0 96324 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1027
timestamp 1623939100
transform 1 0 95588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _450_
timestamp 1623939100
transform 1 0 97060 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1623939100
transform -1 0 98808 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1623939100
transform -1 0 98808 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1623939100
transform 1 0 98164 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_1055
timestamp 1623939100
transform 1 0 98164 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_1047
timestamp 1623939100
transform 1 0 97428 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_1056
timestamp 1623939100
transform 1 0 98256 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1623939100
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1623939100
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1623939100
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1623939100
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1623939100
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1623939100
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_51
timestamp 1623939100
transform 1 0 5796 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_58
timestamp 1623939100
transform 1 0 6440 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_70
timestamp 1623939100
transform 1 0 7544 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1623939100
transform 1 0 8648 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1623939100
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _514_
timestamp 1623939100
transform 1 0 12052 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1623939100
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_106
timestamp 1623939100
transform 1 0 10856 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_115
timestamp 1623939100
transform 1 0 11684 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_128
timestamp 1623939100
transform 1 0 12880 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_140
timestamp 1623939100
transform 1 0 13984 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_152
timestamp 1623939100
transform 1 0 15088 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_164
timestamp 1623939100
transform 1 0 16192 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1623939100
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_170
timestamp 1623939100
transform 1 0 16744 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_172
timestamp 1623939100
transform 1 0 16928 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1623939100
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1623939100
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1623939100
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1623939100
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_220
timestamp 1623939100
transform 1 0 21344 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_229
timestamp 1623939100
transform 1 0 22172 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_241
timestamp 1623939100
transform 1 0 23276 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _418_
timestamp 1623939100
transform 1 0 25852 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_35_253
timestamp 1623939100
transform 1 0 24380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_265
timestamp 1623939100
transform 1 0 25484 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1623939100
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_278
timestamp 1623939100
transform 1 0 26680 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_284
timestamp 1623939100
transform 1 0 27232 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_286
timestamp 1623939100
transform 1 0 27416 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_298
timestamp 1623939100
transform 1 0 28520 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_310
timestamp 1623939100
transform 1 0 29624 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_322
timestamp 1623939100
transform 1 0 30728 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _650_
timestamp 1623939100
transform 1 0 33028 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1623939100
transform 1 0 32568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_354
timestamp 1623939100
transform 1 0 32844 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_334
timestamp 1623939100
transform 1 0 31832 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_343
timestamp 1623939100
transform 1 0 32660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_350
timestamp 1623939100
transform 1 0 33304 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_362
timestamp 1623939100
transform 1 0 34408 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_374
timestamp 1623939100
transform 1 0 35512 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_386
timestamp 1623939100
transform 1 0 36616 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1623939100
transform 1 0 37812 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_398
timestamp 1623939100
transform 1 0 37720 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_400
timestamp 1623939100
transform 1 0 37904 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_412
timestamp 1623939100
transform 1 0 39008 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _698_
timestamp 1623939100
transform -1 0 41492 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1623939100
transform -1 0 39744 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1623939100
transform 1 0 43056 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_439
timestamp 1623939100
transform 1 0 41492 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_451
timestamp 1623939100
transform 1 0 42596 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_455
timestamp 1623939100
transform 1 0 42964 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_457
timestamp 1623939100
transform 1 0 43148 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _618_
timestamp 1623939100
transform 1 0 43792 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_463
timestamp 1623939100
transform 1 0 43700 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_467
timestamp 1623939100
transform 1 0 44068 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_479
timestamp 1623939100
transform 1 0 45172 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_491
timestamp 1623939100
transform 1 0 46276 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1623939100
transform 1 0 48300 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_503
timestamp 1623939100
transform 1 0 47380 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_511
timestamp 1623939100
transform 1 0 48116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_514
timestamp 1623939100
transform 1 0 48392 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_526
timestamp 1623939100
transform 1 0 49496 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_538
timestamp 1623939100
transform 1 0 50600 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _305_
timestamp 1623939100
transform 1 0 51888 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_550
timestamp 1623939100
transform 1 0 51704 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_561
timestamp 1623939100
transform 1 0 52716 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _762_
timestamp 1623939100
transform 1 0 54004 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1623939100
transform 1 0 53544 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_569
timestamp 1623939100
transform 1 0 53452 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_571
timestamp 1623939100
transform 1 0 53636 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_594
timestamp 1623939100
transform 1 0 55752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_606
timestamp 1623939100
transform 1 0 56856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_618
timestamp 1623939100
transform 1 0 57960 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1623939100
transform 1 0 58788 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_626
timestamp 1623939100
transform 1 0 58696 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_628
timestamp 1623939100
transform 1 0 58880 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_640
timestamp 1623939100
transform 1 0 59984 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _503_
timestamp 1623939100
transform 1 0 60628 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_35_646
timestamp 1623939100
transform 1 0 60536 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_656
timestamp 1623939100
transform 1 0 61456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1623939100
transform 1 0 64032 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_668
timestamp 1623939100
transform 1 0 62560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_680
timestamp 1623939100
transform 1 0 63664 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_685
timestamp 1623939100
transform 1 0 64124 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _553_
timestamp 1623939100
transform 1 0 65136 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_693
timestamp 1623939100
transform 1 0 64860 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_699
timestamp 1623939100
transform 1 0 65412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_711
timestamp 1623939100
transform 1 0 66516 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_723
timestamp 1623939100
transform 1 0 67620 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1623939100
transform 1 0 69276 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_735
timestamp 1623939100
transform 1 0 68724 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_742
timestamp 1623939100
transform 1 0 69368 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_754
timestamp 1623939100
transform 1 0 70472 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_766
timestamp 1623939100
transform 1 0 71576 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_778
timestamp 1623939100
transform 1 0 72680 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_790
timestamp 1623939100
transform 1 0 73784 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1623939100
transform 1 0 74520 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_799
timestamp 1623939100
transform 1 0 74612 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_811
timestamp 1623939100
transform 1 0 75716 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_823
timestamp 1623939100
transform 1 0 76820 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_835
timestamp 1623939100
transform 1 0 77924 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_847
timestamp 1623939100
transform 1 0 79028 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1623939100
transform 1 0 79764 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_856
timestamp 1623939100
transform 1 0 79856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_868
timestamp 1623939100
transform 1 0 80960 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _644_
timestamp 1623939100
transform 1 0 82340 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_880
timestamp 1623939100
transform 1 0 82064 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_886
timestamp 1623939100
transform 1 0 82616 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1623939100
transform 1 0 85008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_898
timestamp 1623939100
transform 1 0 83720 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_910
timestamp 1623939100
transform 1 0 84824 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_913
timestamp 1623939100
transform 1 0 85100 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_925
timestamp 1623939100
transform 1 0 86204 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_937
timestamp 1623939100
transform 1 0 87308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_949
timestamp 1623939100
transform 1 0 88412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1623939100
transform 1 0 90252 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_961
timestamp 1623939100
transform 1 0 89516 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_970
timestamp 1623939100
transform 1 0 90344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_982
timestamp 1623939100
transform 1 0 91448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_994
timestamp 1623939100
transform 1 0 92552 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1006
timestamp 1623939100
transform 1 0 93656 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_1018
timestamp 1623939100
transform 1 0 94760 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1623939100
transform 1 0 95496 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1027
timestamp 1623939100
transform 1 0 95588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1039
timestamp 1623939100
transform 1 0 96692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1623939100
transform -1 0 98808 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_1051
timestamp 1623939100
transform 1 0 97796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1623939100
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1623939100
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1623939100
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1623939100
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1623939100
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1623939100
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_42
timestamp 1623939100
transform 1 0 4968 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_54
timestamp 1623939100
transform 1 0 6072 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_66
timestamp 1623939100
transform 1 0 7176 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_78
timestamp 1623939100
transform 1 0 8280 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _408_
timestamp 1623939100
transform 1 0 9752 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1623939100
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_87
timestamp 1623939100
transform 1 0 9108 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_93
timestamp 1623939100
transform 1 0 9660 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_103
timestamp 1623939100
transform 1 0 10580 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_115
timestamp 1623939100
transform 1 0 11684 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1623939100
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_127
timestamp 1623939100
transform 1 0 12788 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_139
timestamp 1623939100
transform 1 0 13892 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_144
timestamp 1623939100
transform 1 0 14352 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1623939100
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1623939100
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1623939100
transform 1 0 17664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1623939100
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_192
timestamp 1623939100
transform 1 0 18768 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1623939100
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_213
timestamp 1623939100
transform 1 0 20700 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_225
timestamp 1623939100
transform 1 0 21804 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_237
timestamp 1623939100
transform 1 0 22908 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_249
timestamp 1623939100
transform 1 0 24012 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1623939100
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1623939100
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_270
timestamp 1623939100
transform 1 0 25944 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_282
timestamp 1623939100
transform 1 0 27048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_294
timestamp 1623939100
transform 1 0 28152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_306
timestamp 1623939100
transform 1 0 29256 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1623939100
transform 1 0 29992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_315
timestamp 1623939100
transform 1 0 30084 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_327
timestamp 1623939100
transform 1 0 31188 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_339
timestamp 1623939100
transform 1 0 32292 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_351
timestamp 1623939100
transform 1 0 33396 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1623939100
transform 1 0 35236 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_363
timestamp 1623939100
transform 1 0 34500 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_372
timestamp 1623939100
transform 1 0 35328 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_384
timestamp 1623939100
transform 1 0 36432 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _390_
timestamp 1623939100
transform 1 0 38088 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_147
timestamp 1623939100
transform 1 0 37904 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_396
timestamp 1623939100
transform 1 0 37536 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_409
timestamp 1623939100
transform 1 0 38732 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1623939100
transform 1 0 40480 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_421
timestamp 1623939100
transform 1 0 39836 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_427
timestamp 1623939100
transform 1 0 40388 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_429
timestamp 1623939100
transform 1 0 40572 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_441
timestamp 1623939100
transform 1 0 41676 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_453
timestamp 1623939100
transform 1 0 42780 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _303_
timestamp 1623939100
transform -1 0 44068 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_210
timestamp 1623939100
transform -1 0 43516 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_467
timestamp 1623939100
transform 1 0 44068 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_479
timestamp 1623939100
transform 1 0 45172 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1623939100
transform 1 0 45724 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_486
timestamp 1623939100
transform 1 0 45816 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_498
timestamp 1623939100
transform 1 0 46920 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_510
timestamp 1623939100
transform 1 0 48024 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_522
timestamp 1623939100
transform 1 0 49128 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_534
timestamp 1623939100
transform 1 0 50232 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _341_
timestamp 1623939100
transform 1 0 52164 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1623939100
transform 1 0 50968 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_543
timestamp 1623939100
transform 1 0 51060 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_561
timestamp 1623939100
transform 1 0 52716 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_573
timestamp 1623939100
transform 1 0 53820 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1623939100
transform 1 0 56212 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_585
timestamp 1623939100
transform 1 0 54924 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_597
timestamp 1623939100
transform 1 0 56028 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_600
timestamp 1623939100
transform 1 0 56304 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _615_
timestamp 1623939100
transform 1 0 58420 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_612
timestamp 1623939100
transform 1 0 57408 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_620
timestamp 1623939100
transform 1 0 58144 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_626
timestamp 1623939100
transform 1 0 58696 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_638
timestamp 1623939100
transform 1 0 59800 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1623939100
transform 1 0 61456 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_650
timestamp 1623939100
transform 1 0 60904 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_657
timestamp 1623939100
transform 1 0 61548 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_669
timestamp 1623939100
transform 1 0 62652 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_681
timestamp 1623939100
transform 1 0 63756 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_693
timestamp 1623939100
transform 1 0 64860 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_705
timestamp 1623939100
transform 1 0 65964 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1623939100
transform 1 0 66700 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_714
timestamp 1623939100
transform 1 0 66792 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_726
timestamp 1623939100
transform 1 0 67896 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_738
timestamp 1623939100
transform 1 0 69000 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_750
timestamp 1623939100
transform 1 0 70104 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1623939100
transform 1 0 71944 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_762
timestamp 1623939100
transform 1 0 71208 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_771
timestamp 1623939100
transform 1 0 72036 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_783
timestamp 1623939100
transform 1 0 73140 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _558_
timestamp 1623939100
transform 1 0 75164 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_795
timestamp 1623939100
transform 1 0 74244 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_803
timestamp 1623939100
transform 1 0 74980 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_808
timestamp 1623939100
transform 1 0 75440 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1623939100
transform 1 0 77188 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_820
timestamp 1623939100
transform 1 0 76544 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_826
timestamp 1623939100
transform 1 0 77096 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_828
timestamp 1623939100
transform 1 0 77280 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_840
timestamp 1623939100
transform 1 0 78384 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_852
timestamp 1623939100
transform 1 0 79488 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_864
timestamp 1623939100
transform 1 0 80592 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1623939100
transform 1 0 82432 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_876
timestamp 1623939100
transform 1 0 81696 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_885
timestamp 1623939100
transform 1 0 82524 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _370_
timestamp 1623939100
transform 1 0 85008 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_145
timestamp 1623939100
transform 1 0 84824 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_897
timestamp 1623939100
transform 1 0 83628 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_909
timestamp 1623939100
transform 1 0 84732 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_928
timestamp 1623939100
transform 1 0 86480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1623939100
transform 1 0 87676 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_940
timestamp 1623939100
transform 1 0 87584 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_942
timestamp 1623939100
transform 1 0 87768 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_954
timestamp 1623939100
transform 1 0 88872 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_966
timestamp 1623939100
transform 1 0 89976 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_978
timestamp 1623939100
transform 1 0 91080 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1623939100
transform 1 0 92920 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_990
timestamp 1623939100
transform 1 0 92184 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_999
timestamp 1623939100
transform 1 0 93012 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1011
timestamp 1623939100
transform 1 0 94116 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1023
timestamp 1623939100
transform 1 0 95220 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1035
timestamp 1623939100
transform 1 0 96324 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1623939100
transform -1 0 98808 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1623939100
transform 1 0 98164 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_1047
timestamp 1623939100
transform 1 0 97428 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_1056
timestamp 1623939100
transform 1 0 98256 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1623939100
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1623939100
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1623939100
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1623939100
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1623939100
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1623939100
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_51
timestamp 1623939100
transform 1 0 5796 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_58
timestamp 1623939100
transform 1 0 6440 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_70
timestamp 1623939100
transform 1 0 7544 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_82
timestamp 1623939100
transform 1 0 8648 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_94
timestamp 1623939100
transform 1 0 9752 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1623939100
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_106
timestamp 1623939100
transform 1 0 10856 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_115
timestamp 1623939100
transform 1 0 11684 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_127
timestamp 1623939100
transform 1 0 12788 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_139
timestamp 1623939100
transform 1 0 13892 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_145
timestamp 1623939100
transform 1 0 14444 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _639_
timestamp 1623939100
transform 1 0 14720 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_343
timestamp 1623939100
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1623939100
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_163
timestamp 1623939100
transform 1 0 16100 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1623939100
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_172
timestamp 1623939100
transform 1 0 16928 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1623939100
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1623939100
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1623939100
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1623939100
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_220
timestamp 1623939100
transform 1 0 21344 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_229
timestamp 1623939100
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_241
timestamp 1623939100
transform 1 0 23276 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_253
timestamp 1623939100
transform 1 0 24380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_265
timestamp 1623939100
transform 1 0 25484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1623939100
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_277
timestamp 1623939100
transform 1 0 26588 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_286
timestamp 1623939100
transform 1 0 27416 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_298
timestamp 1623939100
transform 1 0 28520 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_310
timestamp 1623939100
transform 1 0 29624 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_322
timestamp 1623939100
transform 1 0 30728 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _717_
timestamp 1623939100
transform 1 0 33672 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1623939100
transform 1 0 32568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1623939100
transform 1 0 33488 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_334
timestamp 1623939100
transform 1 0 31832 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_343
timestamp 1623939100
transform 1 0 32660 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_351
timestamp 1623939100
transform 1 0 33396 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1623939100
transform 1 0 35420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_385
timestamp 1623939100
transform 1 0 36524 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1623939100
transform 1 0 37812 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_397
timestamp 1623939100
transform 1 0 37628 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_400
timestamp 1623939100
transform 1 0 37904 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_412
timestamp 1623939100
transform 1 0 39008 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_424
timestamp 1623939100
transform 1 0 40112 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_436
timestamp 1623939100
transform 1 0 41216 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1623939100
transform 1 0 43056 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_448
timestamp 1623939100
transform 1 0 42320 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_457
timestamp 1623939100
transform 1 0 43148 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_469
timestamp 1623939100
transform 1 0 44252 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_481
timestamp 1623939100
transform 1 0 45356 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_493
timestamp 1623939100
transform 1 0 46460 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1623939100
transform 1 0 48300 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1623939100
transform 1 0 47564 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_514
timestamp 1623939100
transform 1 0 48392 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_526
timestamp 1623939100
transform 1 0 49496 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_538
timestamp 1623939100
transform 1 0 50600 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_550
timestamp 1623939100
transform 1 0 51704 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_562
timestamp 1623939100
transform 1 0 52808 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1623939100
transform 1 0 53544 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_571
timestamp 1623939100
transform 1 0 53636 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_583
timestamp 1623939100
transform 1 0 54740 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_595
timestamp 1623939100
transform 1 0 55844 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_607
timestamp 1623939100
transform 1 0 56948 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_619
timestamp 1623939100
transform 1 0 58052 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1623939100
transform 1 0 58788 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_628
timestamp 1623939100
transform 1 0 58880 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_640
timestamp 1623939100
transform 1 0 59984 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_652
timestamp 1623939100
transform 1 0 61088 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_664
timestamp 1623939100
transform 1 0 62192 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1623939100
transform 1 0 64032 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_676
timestamp 1623939100
transform 1 0 63296 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_685
timestamp 1623939100
transform 1 0 64124 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _394_
timestamp 1623939100
transform 1 0 65136 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_390
timestamp 1623939100
transform 1 0 64952 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_693
timestamp 1623939100
transform 1 0 64860 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_705
timestamp 1623939100
transform 1 0 65964 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_717
timestamp 1623939100
transform 1 0 67068 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_729
timestamp 1623939100
transform 1 0 68172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1623939100
transform 1 0 69276 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_742
timestamp 1623939100
transform 1 0 69368 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_754
timestamp 1623939100
transform 1 0 70472 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_766
timestamp 1623939100
transform 1 0 71576 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_778
timestamp 1623939100
transform 1 0 72680 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_790
timestamp 1623939100
transform 1 0 73784 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _502_
timestamp 1623939100
transform 1 0 74980 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1623939100
transform 1 0 74520 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_799
timestamp 1623939100
transform 1 0 74612 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_809
timestamp 1623939100
transform 1 0 75532 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _619_
timestamp 1623939100
transform 1 0 75900 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_816
timestamp 1623939100
transform 1 0 76176 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_828
timestamp 1623939100
transform 1 0 77280 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_840
timestamp 1623939100
transform 1 0 78384 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_852
timestamp 1623939100
transform 1 0 79488 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1623939100
transform 1 0 79764 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_856
timestamp 1623939100
transform 1 0 79856 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_868
timestamp 1623939100
transform 1 0 80960 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_880
timestamp 1623939100
transform 1 0 82064 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_892
timestamp 1623939100
transform 1 0 83168 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1623939100
transform 1 0 85008 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_904
timestamp 1623939100
transform 1 0 84272 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_913
timestamp 1623939100
transform 1 0 85100 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_925
timestamp 1623939100
transform 1 0 86204 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_937
timestamp 1623939100
transform 1 0 87308 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_949
timestamp 1623939100
transform 1 0 88412 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1623939100
transform 1 0 90252 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_961
timestamp 1623939100
transform 1 0 89516 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_970
timestamp 1623939100
transform 1 0 90344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_982
timestamp 1623939100
transform 1 0 91448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_994
timestamp 1623939100
transform 1 0 92552 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1006
timestamp 1623939100
transform 1 0 93656 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1018
timestamp 1623939100
transform 1 0 94760 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1623939100
transform 1 0 95496 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1027
timestamp 1623939100
transform 1 0 95588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1039
timestamp 1623939100
transform 1 0 96692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1623939100
transform -1 0 98808 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1051
timestamp 1623939100
transform 1 0 97796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1623939100
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1623939100
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1623939100
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1623939100
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1623939100
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_30
timestamp 1623939100
transform 1 0 3864 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_42
timestamp 1623939100
transform 1 0 4968 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_54
timestamp 1623939100
transform 1 0 6072 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_66
timestamp 1623939100
transform 1 0 7176 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_78
timestamp 1623939100
transform 1 0 8280 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _732_
timestamp 1623939100
transform 1 0 9476 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1623939100
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_87
timestamp 1623939100
transform 1 0 9108 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_110
timestamp 1623939100
transform 1 0 11224 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_122
timestamp 1623939100
transform 1 0 12328 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1623939100
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_134
timestamp 1623939100
transform 1 0 13432 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_142
timestamp 1623939100
transform 1 0 14168 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_144
timestamp 1623939100
transform 1 0 14352 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _372_
timestamp 1623939100
transform 1 0 14720 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_38_155
timestamp 1623939100
transform 1 0 15364 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_167
timestamp 1623939100
transform 1 0 16468 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_179
timestamp 1623939100
transform 1 0 17572 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1623939100
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_191
timestamp 1623939100
transform 1 0 18676 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_199
timestamp 1623939100
transform 1 0 19412 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_201
timestamp 1623939100
transform 1 0 19596 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_213
timestamp 1623939100
transform 1 0 20700 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_225
timestamp 1623939100
transform 1 0 21804 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_237
timestamp 1623939100
transform 1 0 22908 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_249
timestamp 1623939100
transform 1 0 24012 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _533_
timestamp 1623939100
transform 1 0 25760 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1623939100
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_258
timestamp 1623939100
transform 1 0 24840 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_266
timestamp 1623939100
transform 1 0 25576 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1623939100
transform 1 0 26588 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1623939100
transform 1 0 27692 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_301
timestamp 1623939100
transform 1 0 28796 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1623939100
transform 1 0 29992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_313
timestamp 1623939100
transform 1 0 29900 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_315
timestamp 1623939100
transform 1 0 30084 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_327
timestamp 1623939100
transform 1 0 31188 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_339
timestamp 1623939100
transform 1 0 32292 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_351
timestamp 1623939100
transform 1 0 33396 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1623939100
transform 1 0 35236 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_363
timestamp 1623939100
transform 1 0 34500 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_372
timestamp 1623939100
transform 1 0 35328 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_384
timestamp 1623939100
transform 1 0 36432 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_396
timestamp 1623939100
transform 1 0 37536 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_408
timestamp 1623939100
transform 1 0 38640 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1623939100
transform 1 0 40480 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_420
timestamp 1623939100
transform 1 0 39744 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_429
timestamp 1623939100
transform 1 0 40572 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_441
timestamp 1623939100
transform 1 0 41676 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_453
timestamp 1623939100
transform 1 0 42780 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_465
timestamp 1623939100
transform 1 0 43884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_477
timestamp 1623939100
transform 1 0 44988 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1623939100
transform 1 0 45724 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_486
timestamp 1623939100
transform 1 0 45816 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_498
timestamp 1623939100
transform 1 0 46920 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _291_
timestamp 1623939100
transform -1 0 48484 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_129
timestamp 1623939100
transform -1 0 47656 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_130
timestamp 1623939100
transform -1 0 48668 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_187
timestamp 1623939100
transform -1 0 47472 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_188
timestamp 1623939100
transform -1 0 48852 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_519
timestamp 1623939100
transform 1 0 48852 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_531
timestamp 1623939100
transform 1 0 49956 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_539
timestamp 1623939100
transform 1 0 50692 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1623939100
transform 1 0 50968 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_543
timestamp 1623939100
transform 1 0 51060 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_555
timestamp 1623939100
transform 1 0 52164 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_567
timestamp 1623939100
transform 1 0 53268 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_579
timestamp 1623939100
transform 1 0 54372 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1623939100
transform 1 0 56212 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_591
timestamp 1623939100
transform 1 0 55476 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_600
timestamp 1623939100
transform 1 0 56304 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_612
timestamp 1623939100
transform 1 0 57408 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_624
timestamp 1623939100
transform 1 0 58512 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_636
timestamp 1623939100
transform 1 0 59616 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _508_
timestamp 1623939100
transform 1 0 61916 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1623939100
transform 1 0 61456 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_168
timestamp 1623939100
transform 1 0 61732 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_648
timestamp 1623939100
transform 1 0 60720 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_657
timestamp 1623939100
transform 1 0 61548 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_670
timestamp 1623939100
transform 1 0 62744 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_682
timestamp 1623939100
transform 1 0 63848 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_694
timestamp 1623939100
transform 1 0 64952 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_706
timestamp 1623939100
transform 1 0 66056 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _737_
timestamp 1623939100
transform 1 0 67436 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1623939100
transform 1 0 66700 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_712
timestamp 1623939100
transform 1 0 66608 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_714
timestamp 1623939100
transform 1 0 66792 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_720
timestamp 1623939100
transform 1 0 67344 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  _518_
timestamp 1623939100
transform 1 0 70012 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_38_740
timestamp 1623939100
transform 1 0 69184 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_748
timestamp 1623939100
transform 1 0 69920 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1623939100
transform 1 0 71944 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_758
timestamp 1623939100
transform 1 0 70840 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _345_
timestamp 1623939100
transform 1 0 72588 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_143
timestamp 1623939100
transform 1 0 72404 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_381
timestamp 1623939100
transform 1 0 73416 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_771
timestamp 1623939100
transform 1 0 72036 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_788
timestamp 1623939100
transform 1 0 73600 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_800
timestamp 1623939100
transform 1 0 74704 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_812
timestamp 1623939100
transform 1 0 75808 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1623939100
transform 1 0 77188 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_824
timestamp 1623939100
transform 1 0 76912 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_828
timestamp 1623939100
transform 1 0 77280 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_840
timestamp 1623939100
transform 1 0 78384 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_852
timestamp 1623939100
transform 1 0 79488 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_864
timestamp 1623939100
transform 1 0 80592 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1623939100
transform 1 0 82432 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_876
timestamp 1623939100
transform 1 0 81696 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_885
timestamp 1623939100
transform 1 0 82524 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_897
timestamp 1623939100
transform 1 0 83628 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_909
timestamp 1623939100
transform 1 0 84732 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_921
timestamp 1623939100
transform 1 0 85836 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_933
timestamp 1623939100
transform 1 0 86940 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1623939100
transform 1 0 87676 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_942
timestamp 1623939100
transform 1 0 87768 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_954
timestamp 1623939100
transform 1 0 88872 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_966
timestamp 1623939100
transform 1 0 89976 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_978
timestamp 1623939100
transform 1 0 91080 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1623939100
transform 1 0 92920 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_990
timestamp 1623939100
transform 1 0 92184 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_999
timestamp 1623939100
transform 1 0 93012 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1011
timestamp 1623939100
transform 1 0 94116 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1023
timestamp 1623939100
transform 1 0 95220 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1035
timestamp 1623939100
transform 1 0 96324 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1623939100
transform -1 0 98808 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1623939100
transform 1 0 98164 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_1047
timestamp 1623939100
transform 1 0 97428 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_1056
timestamp 1623939100
transform 1 0 98256 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _282_
timestamp 1623939100
transform 1 0 2944 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1623939100
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1623939100
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1623939100
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1623939100
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1623939100
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_15
timestamp 1623939100
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_19
timestamp 1623939100
transform 1 0 2852 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _658_
timestamp 1623939100
transform 1 0 4600 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1623939100
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_361
timestamp 1623939100
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_27
timestamp 1623939100
transform 1 0 3588 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_35
timestamp 1623939100
transform 1 0 4324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_41
timestamp 1623939100
transform 1 0 4876 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_25
timestamp 1623939100
transform 1 0 3404 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_30
timestamp 1623939100
transform 1 0 3864 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1623939100
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_53
timestamp 1623939100
transform 1 0 5980 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_58
timestamp 1623939100
transform 1 0 6440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_42
timestamp 1623939100
transform 1 0 4968 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_54
timestamp 1623939100
transform 1 0 6072 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_70
timestamp 1623939100
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_82
timestamp 1623939100
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_66
timestamp 1623939100
transform 1 0 7176 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_78
timestamp 1623939100
transform 1 0 8280 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1623939100
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_94
timestamp 1623939100
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_87
timestamp 1623939100
transform 1 0 9108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_99
timestamp 1623939100
transform 1 0 10212 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1623939100
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_106
timestamp 1623939100
transform 1 0 10856 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_115
timestamp 1623939100
transform 1 0 11684 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_111
timestamp 1623939100
transform 1 0 11316 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1623939100
transform 1 0 12420 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _635_
timestamp 1623939100
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1623939100
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_127
timestamp 1623939100
transform 1 0 12788 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_139
timestamp 1623939100
transform 1 0 13892 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_135
timestamp 1623939100
transform 1 0 13524 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1623939100
transform 1 0 14352 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _479_
timestamp 1623939100
transform -1 0 17572 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_155
timestamp 1623939100
transform -1 0 16100 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_146
timestamp 1623939100
transform 1 0 14536 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_158
timestamp 1623939100
transform 1 0 15640 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_156
timestamp 1623939100
transform 1 0 15456 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_160
timestamp 1623939100
transform 1 0 15824 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1623939100
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_190
timestamp 1623939100
transform -1 0 17756 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_170
timestamp 1623939100
transform 1 0 16744 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_172
timestamp 1623939100
transform 1 0 16928 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1623939100
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_181
timestamp 1623939100
transform 1 0 17756 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1623939100
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1623939100
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1623939100
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_193
timestamp 1623939100
transform 1 0 18860 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_199
timestamp 1623939100
transform 1 0 19412 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_201
timestamp 1623939100
transform 1 0 19596 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _758_
timestamp 1623939100
transform 1 0 20424 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1623939100
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_220
timestamp 1623939100
transform 1 0 21344 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_229
timestamp 1623939100
transform 1 0 22172 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_209
timestamp 1623939100
transform 1 0 20332 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_229
timestamp 1623939100
transform 1 0 22172 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  _338_
timestamp 1623939100
transform 1 0 22540 0 -1 24480
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_39_241
timestamp 1623939100
transform 1 0 23276 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_244
timestamp 1623939100
transform 1 0 23552 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _542_
timestamp 1623939100
transform 1 0 24932 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1623939100
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_253
timestamp 1623939100
transform 1 0 24380 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_268
timestamp 1623939100
transform 1 0 25760 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_256
timestamp 1623939100
transform 1 0 24656 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_258
timestamp 1623939100
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_270
timestamp 1623939100
transform 1 0 25944 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1623939100
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_280
timestamp 1623939100
transform 1 0 26864 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_284
timestamp 1623939100
transform 1 0 27232 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_286
timestamp 1623939100
transform 1 0 27416 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_282
timestamp 1623939100
transform 1 0 27048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_298
timestamp 1623939100
transform 1 0 28520 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_310
timestamp 1623939100
transform 1 0 29624 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_294
timestamp 1623939100
transform 1 0 28152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_306
timestamp 1623939100
transform 1 0 29256 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1623939100
transform 1 0 29992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_322
timestamp 1623939100
transform 1 0 30728 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_315
timestamp 1623939100
transform 1 0 30084 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_327
timestamp 1623939100
transform 1 0 31188 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1623939100
transform 1 0 32568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_334
timestamp 1623939100
transform 1 0 31832 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_343
timestamp 1623939100
transform 1 0 32660 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_339
timestamp 1623939100
transform 1 0 32292 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_351
timestamp 1623939100
transform 1 0 33396 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1623939100
transform 1 0 35236 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_355
timestamp 1623939100
transform 1 0 33764 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_367
timestamp 1623939100
transform 1 0 34868 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_363
timestamp 1623939100
transform 1 0 34500 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_372
timestamp 1623939100
transform 1 0 35328 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _638_
timestamp 1623939100
transform 1 0 36156 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_379
timestamp 1623939100
transform 1 0 35972 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_391
timestamp 1623939100
transform 1 0 37076 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_380
timestamp 1623939100
transform 1 0 36064 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_384
timestamp 1623939100
transform 1 0 36432 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1623939100
transform 1 0 37812 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_400
timestamp 1623939100
transform 1 0 37904 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_412
timestamp 1623939100
transform 1 0 39008 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_396
timestamp 1623939100
transform 1 0 37536 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_408
timestamp 1623939100
transform 1 0 38640 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1623939100
transform 1 0 40480 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  repeater608
timestamp 1623939100
transform 1 0 40940 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_424
timestamp 1623939100
transform 1 0 40112 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_436
timestamp 1623939100
transform 1 0 41216 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_420
timestamp 1623939100
transform 1 0 39744 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_429
timestamp 1623939100
transform 1 0 40572 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_437
timestamp 1623939100
transform 1 0 41308 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1623939100
transform 1 0 43056 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_448
timestamp 1623939100
transform 1 0 42320 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_457
timestamp 1623939100
transform 1 0 43148 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_449
timestamp 1623939100
transform 1 0 42412 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_469
timestamp 1623939100
transform 1 0 44252 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_461
timestamp 1623939100
transform 1 0 43516 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_473
timestamp 1623939100
transform 1 0 44620 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _329_
timestamp 1623939100
transform 1 0 46184 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1623939100
transform 1 0 45724 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_481
timestamp 1623939100
transform 1 0 45356 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_493
timestamp 1623939100
transform 1 0 46460 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_486
timestamp 1623939100
transform 1 0 45816 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_497
timestamp 1623939100
transform 1 0 46828 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _768_
timestamp 1623939100
transform 1 0 48760 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1623939100
transform 1 0 48300 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1623939100
transform 1 0 47564 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_514
timestamp 1623939100
transform 1 0 48392 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_509
timestamp 1623939100
transform 1 0 47932 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_537
timestamp 1623939100
transform 1 0 50508 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_521
timestamp 1623939100
transform 1 0 49036 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_533
timestamp 1623939100
transform 1 0 50140 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_541
timestamp 1623939100
transform 1 0 50876 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1623939100
transform 1 0 50968 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_549
timestamp 1623939100
transform 1 0 51612 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_561
timestamp 1623939100
transform 1 0 52716 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_543
timestamp 1623939100
transform 1 0 51060 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_555
timestamp 1623939100
transform 1 0 52164 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1623939100
transform 1 0 53544 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_569
timestamp 1623939100
transform 1 0 53452 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_571
timestamp 1623939100
transform 1 0 53636 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_583
timestamp 1623939100
transform 1 0 54740 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_567
timestamp 1623939100
transform 1 0 53268 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_579
timestamp 1623939100
transform 1 0 54372 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1623939100
transform 1 0 56212 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_595
timestamp 1623939100
transform 1 0 55844 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_591
timestamp 1623939100
transform 1 0 55476 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_600
timestamp 1623939100
transform 1 0 56304 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_607
timestamp 1623939100
transform 1 0 56948 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_619
timestamp 1623939100
transform 1 0 58052 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_612
timestamp 1623939100
transform 1 0 57408 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_624
timestamp 1623939100
transform 1 0 58512 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1623939100
transform 1 0 58788 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_628
timestamp 1623939100
transform 1 0 58880 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_640
timestamp 1623939100
transform 1 0 59984 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_636
timestamp 1623939100
transform 1 0 59616 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1623939100
transform 1 0 61456 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_652
timestamp 1623939100
transform 1 0 61088 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_664
timestamp 1623939100
transform 1 0 62192 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_648
timestamp 1623939100
transform 1 0 60720 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_657
timestamp 1623939100
transform 1 0 61548 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1623939100
transform 1 0 64032 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_676
timestamp 1623939100
transform 1 0 63296 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_685
timestamp 1623939100
transform 1 0 64124 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_669
timestamp 1623939100
transform 1 0 62652 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_681
timestamp 1623939100
transform 1 0 63756 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _596_
timestamp 1623939100
transform 1 0 65320 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform -1 0 66516 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1623939100
transform -1 0 65688 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_697
timestamp 1623939100
transform 1 0 65228 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_693
timestamp 1623939100
transform 1 0 64860 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_697
timestamp 1623939100
transform 1 0 65228 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_701
timestamp 1623939100
transform 1 0 65596 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1623939100
transform 1 0 66700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_711
timestamp 1623939100
transform 1 0 66516 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_723
timestamp 1623939100
transform 1 0 67620 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_714
timestamp 1623939100
transform 1 0 66792 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_726
timestamp 1623939100
transform 1 0 67896 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _597_
timestamp 1623939100
transform 1 0 69736 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1623939100
transform 1 0 69276 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_735
timestamp 1623939100
transform 1 0 68724 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_742
timestamp 1623939100
transform 1 0 69368 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_749
timestamp 1623939100
transform 1 0 70012 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_738
timestamp 1623939100
transform 1 0 69000 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_750
timestamp 1623939100
transform 1 0 70104 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1623939100
transform 1 0 71944 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_761
timestamp 1623939100
transform 1 0 71116 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_769
timestamp 1623939100
transform 1 0 71852 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_762
timestamp 1623939100
transform 1 0 71208 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _428_
timestamp 1623939100
transform 1 0 72220 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_154
timestamp 1623939100
transform 1 0 72036 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_779
timestamp 1623939100
transform 1 0 72772 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_791
timestamp 1623939100
transform 1 0 73876 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_771
timestamp 1623939100
transform 1 0 72036 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_783
timestamp 1623939100
transform 1 0 73140 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _403_
timestamp 1623939100
transform 1 0 75532 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _759_
timestamp 1623939100
transform 1 0 74980 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1623939100
transform 1 0 74520 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_149
timestamp 1623939100
transform 1 0 75348 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_797
timestamp 1623939100
transform 1 0 74428 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_799
timestamp 1623939100
transform 1 0 74612 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_795
timestamp 1623939100
transform 1 0 74244 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _349_
timestamp 1623939100
transform 1 0 76912 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1623939100
transform 1 0 77188 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_140
timestamp 1623939100
transform 1 0 76728 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_185
timestamp 1623939100
transform 1 0 76176 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_820
timestamp 1623939100
transform 1 0 76544 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_830
timestamp 1623939100
transform 1 0 77464 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_818
timestamp 1623939100
transform 1 0 76360 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_826
timestamp 1623939100
transform 1 0 77096 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_828
timestamp 1623939100
transform 1 0 77280 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _569_
timestamp 1623939100
transform 1 0 78936 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_842
timestamp 1623939100
transform 1 0 78568 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_849
timestamp 1623939100
transform 1 0 79212 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_840
timestamp 1623939100
transform 1 0 78384 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_852
timestamp 1623939100
transform 1 0 79488 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _573_
timestamp 1623939100
transform -1 0 80500 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1623939100
transform 1 0 79764 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_331
timestamp 1623939100
transform -1 0 80224 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_856
timestamp 1623939100
transform 1 0 79856 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_863
timestamp 1623939100
transform 1 0 80500 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_875
timestamp 1623939100
transform 1 0 81604 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_864
timestamp 1623939100
transform 1 0 80592 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _404_
timestamp 1623939100
transform 1 0 82984 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1623939100
transform 1 0 82432 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_887
timestamp 1623939100
transform 1 0 82708 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_876
timestamp 1623939100
transform 1 0 81696 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_885
timestamp 1623939100
transform 1 0 82524 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_889
timestamp 1623939100
transform 1 0 82892 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1623939100
transform 1 0 85008 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_899
timestamp 1623939100
transform 1 0 83812 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_911
timestamp 1623939100
transform 1 0 84916 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_913
timestamp 1623939100
transform 1 0 85100 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_899
timestamp 1623939100
transform 1 0 83812 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_911
timestamp 1623939100
transform 1 0 84916 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_925
timestamp 1623939100
transform 1 0 86204 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_937
timestamp 1623939100
transform 1 0 87308 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_923
timestamp 1623939100
transform 1 0 86020 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_935
timestamp 1623939100
transform 1 0 87124 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1623939100
transform 1 0 87676 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_949
timestamp 1623939100
transform 1 0 88412 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_942
timestamp 1623939100
transform 1 0 87768 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_954
timestamp 1623939100
transform 1 0 88872 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1623939100
transform 1 0 90252 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_961
timestamp 1623939100
transform 1 0 89516 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_970
timestamp 1623939100
transform 1 0 90344 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_966
timestamp 1623939100
transform 1 0 89976 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_978
timestamp 1623939100
transform 1 0 91080 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1623939100
transform 1 0 92920 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_982
timestamp 1623939100
transform 1 0 91448 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_994
timestamp 1623939100
transform 1 0 92552 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_990
timestamp 1623939100
transform 1 0 92184 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_999
timestamp 1623939100
transform 1 0 93012 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1006
timestamp 1623939100
transform 1 0 93656 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1018
timestamp 1623939100
transform 1 0 94760 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1011
timestamp 1623939100
transform 1 0 94116 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _729_
timestamp 1623939100
transform 1 0 95956 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1623939100
transform 1 0 95496 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1623939100
transform 1 0 95772 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1623939100
transform 1 0 95588 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_57
timestamp 1623939100
transform 1 0 95312 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1023
timestamp 1623939100
transform 1 0 95220 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1035
timestamp 1623939100
transform 1 0 96324 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1623939100
transform -1 0 98808 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1623939100
transform -1 0 98808 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1623939100
transform 1 0 98164 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1623939100
transform 1 0 97704 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1623939100
transform 1 0 97888 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1623939100
transform 1 0 98072 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_1056
timestamp 1623939100
transform 1 0 98256 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_1047
timestamp 1623939100
transform 1 0 97428 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_1056
timestamp 1623939100
transform 1 0 98256 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_4  _369_
timestamp 1623939100
transform 1 0 2668 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__o221a_2  _489_
timestamp 1623939100
transform 1 0 1472 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1623939100
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_166
timestamp 1623939100
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_198
timestamp 1623939100
transform 1 0 2484 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_3
timestamp 1623939100
transform 1 0 1380 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_31
timestamp 1623939100
transform 1 0 3956 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1623939100
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_43
timestamp 1623939100
transform 1 0 5060 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_55
timestamp 1623939100
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_58
timestamp 1623939100
transform 1 0 6440 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_70
timestamp 1623939100
transform 1 0 7544 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_82
timestamp 1623939100
transform 1 0 8648 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1623939100
transform 1 0 9752 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _663_
timestamp 1623939100
transform 1 0 12236 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1623939100
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_368
timestamp 1623939100
transform 1 0 12052 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_106
timestamp 1623939100
transform 1 0 10856 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_115
timestamp 1623939100
transform 1 0 11684 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_124
timestamp 1623939100
transform 1 0 12512 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_136
timestamp 1623939100
transform 1 0 13616 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_148
timestamp 1623939100
transform 1 0 14720 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp 1623939100
transform 1 0 15824 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1623939100
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_168
timestamp 1623939100
transform 1 0 16560 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_172
timestamp 1623939100
transform 1 0 16928 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1623939100
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1623939100
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1623939100
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1623939100
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_220
timestamp 1623939100
transform 1 0 21344 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_229
timestamp 1623939100
transform 1 0 22172 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_241
timestamp 1623939100
transform 1 0 23276 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_253
timestamp 1623939100
transform 1 0 24380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_265
timestamp 1623939100
transform 1 0 25484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1623939100
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_277
timestamp 1623939100
transform 1 0 26588 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_286
timestamp 1623939100
transform 1 0 27416 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  _525_
timestamp 1623939100
transform 1 0 29808 0 1 24480
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_41_298
timestamp 1623939100
transform 1 0 28520 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_310
timestamp 1623939100
transform 1 0 29624 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_323
timestamp 1623939100
transform 1 0 30820 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1623939100
transform 1 0 32568 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_335
timestamp 1623939100
transform 1 0 31924 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_341
timestamp 1623939100
transform 1 0 32476 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_343
timestamp 1623939100
transform 1 0 32660 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_355
timestamp 1623939100
transform 1 0 33764 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_367
timestamp 1623939100
transform 1 0 34868 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_379
timestamp 1623939100
transform 1 0 35972 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_391
timestamp 1623939100
transform 1 0 37076 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_912
timestamp 1623939100
transform 1 0 37812 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_400
timestamp 1623939100
transform 1 0 37904 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_412
timestamp 1623939100
transform 1 0 39008 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_424
timestamp 1623939100
transform 1 0 40112 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_436
timestamp 1623939100
transform 1 0 41216 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_913
timestamp 1623939100
transform 1 0 43056 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_448
timestamp 1623939100
transform 1 0 42320 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_457
timestamp 1623939100
transform 1 0 43148 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _741_
timestamp 1623939100
transform 1 0 43516 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_41_480
timestamp 1623939100
transform 1 0 45264 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_492
timestamp 1623939100
transform 1 0 46368 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_914
timestamp 1623939100
transform 1 0 48300 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_504
timestamp 1623939100
transform 1 0 47472 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_512
timestamp 1623939100
transform 1 0 48208 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_514
timestamp 1623939100
transform 1 0 48392 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _735_
timestamp 1623939100
transform 1 0 50876 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_41_526
timestamp 1623939100
transform 1 0 49496 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_538
timestamp 1623939100
transform 1 0 50600 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_560
timestamp 1623939100
transform 1 0 52624 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_915
timestamp 1623939100
transform 1 0 53544 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_568
timestamp 1623939100
transform 1 0 53360 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_571
timestamp 1623939100
transform 1 0 53636 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_583
timestamp 1623939100
transform 1 0 54740 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_595
timestamp 1623939100
transform 1 0 55844 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_607
timestamp 1623939100
transform 1 0 56948 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_619
timestamp 1623939100
transform 1 0 58052 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_916
timestamp 1623939100
transform 1 0 58788 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_628
timestamp 1623939100
transform 1 0 58880 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_640
timestamp 1623939100
transform 1 0 59984 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_652
timestamp 1623939100
transform 1 0 61088 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_664
timestamp 1623939100
transform 1 0 62192 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_917
timestamp 1623939100
transform 1 0 64032 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_676
timestamp 1623939100
transform 1 0 63296 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_685
timestamp 1623939100
transform 1 0 64124 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_697
timestamp 1623939100
transform 1 0 65228 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_709
timestamp 1623939100
transform 1 0 66332 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_721
timestamp 1623939100
transform 1 0 67436 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_918
timestamp 1623939100
transform 1 0 69276 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_733
timestamp 1623939100
transform 1 0 68540 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_742
timestamp 1623939100
transform 1 0 69368 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _689_
timestamp 1623939100
transform 1 0 71208 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_754
timestamp 1623939100
transform 1 0 70472 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_765
timestamp 1623939100
transform 1 0 71484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_777
timestamp 1623939100
transform 1 0 72588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_789
timestamp 1623939100
transform 1 0 73692 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_919
timestamp 1623939100
transform 1 0 74520 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_797
timestamp 1623939100
transform 1 0 74428 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_799
timestamp 1623939100
transform 1 0 74612 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_811
timestamp 1623939100
transform 1 0 75716 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _747_
timestamp 1623939100
transform -1 0 78384 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_85
timestamp 1623939100
transform -1 0 76636 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_87
timestamp 1623939100
transform -1 0 76452 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_89
timestamp 1623939100
transform -1 0 76268 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_86
timestamp 1623939100
transform -1 0 78568 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_88
timestamp 1623939100
transform -1 0 78752 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_90
timestamp 1623939100
transform -1 0 78936 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_846
timestamp 1623939100
transform 1 0 78936 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_854
timestamp 1623939100
transform 1 0 79672 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_920
timestamp 1623939100
transform 1 0 79764 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_856
timestamp 1623939100
transform 1 0 79856 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_868
timestamp 1623939100
transform 1 0 80960 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_880
timestamp 1623939100
transform 1 0 82064 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_892
timestamp 1623939100
transform 1 0 83168 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_921
timestamp 1623939100
transform 1 0 85008 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_904
timestamp 1623939100
transform 1 0 84272 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_913
timestamp 1623939100
transform 1 0 85100 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_925
timestamp 1623939100
transform 1 0 86204 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_937
timestamp 1623939100
transform 1 0 87308 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_949
timestamp 1623939100
transform 1 0 88412 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_922
timestamp 1623939100
transform 1 0 90252 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_961
timestamp 1623939100
transform 1 0 89516 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_970
timestamp 1623939100
transform 1 0 90344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_982
timestamp 1623939100
transform 1 0 91448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_994
timestamp 1623939100
transform 1 0 92552 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1006
timestamp 1623939100
transform 1 0 93656 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_1018
timestamp 1623939100
transform 1 0 94760 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_923
timestamp 1623939100
transform 1 0 95496 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1027
timestamp 1623939100
transform 1 0 95588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1039
timestamp 1623939100
transform 1 0 96692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1623939100
transform -1 0 98808 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_1051
timestamp 1623939100
transform 1 0 97796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1623939100
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1623939100
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1623939100
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_924
timestamp 1623939100
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_27
timestamp 1623939100
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_30
timestamp 1623939100
transform 1 0 3864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_42
timestamp 1623939100
transform 1 0 4968 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_54
timestamp 1623939100
transform 1 0 6072 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_66
timestamp 1623939100
transform 1 0 7176 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_78
timestamp 1623939100
transform 1 0 8280 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_925
timestamp 1623939100
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_87
timestamp 1623939100
transform 1 0 9108 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_99
timestamp 1623939100
transform 1 0 10212 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_111
timestamp 1623939100
transform 1 0 11316 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_123
timestamp 1623939100
transform 1 0 12420 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_926
timestamp 1623939100
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_135
timestamp 1623939100
transform 1 0 13524 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_144
timestamp 1623939100
transform 1 0 14352 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1623939100
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1623939100
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1623939100
transform 1 0 17664 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_927
timestamp 1623939100
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_192
timestamp 1623939100
transform 1 0 18768 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1623939100
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _306_
timestamp 1623939100
transform -1 0 22080 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_209
timestamp 1623939100
transform -1 0 21528 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_213
timestamp 1623939100
transform 1 0 20700 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_219
timestamp 1623939100
transform 1 0 21252 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_228
timestamp 1623939100
transform 1 0 22080 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_240
timestamp 1623939100
transform 1 0 23184 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_928
timestamp 1623939100
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_252
timestamp 1623939100
transform 1 0 24288 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_256
timestamp 1623939100
transform 1 0 24656 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_258
timestamp 1623939100
transform 1 0 24840 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_270
timestamp 1623939100
transform 1 0 25944 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _616_
timestamp 1623939100
transform 1 0 27508 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_282
timestamp 1623939100
transform 1 0 27048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_286
timestamp 1623939100
transform 1 0 27416 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_290
timestamp 1623939100
transform 1 0 27784 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_302
timestamp 1623939100
transform 1 0 28888 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_929
timestamp 1623939100
transform 1 0 29992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_315
timestamp 1623939100
transform 1 0 30084 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_327
timestamp 1623939100
transform 1 0 31188 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_339
timestamp 1623939100
transform 1 0 32292 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_351
timestamp 1623939100
transform 1 0 33396 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_930
timestamp 1623939100
transform 1 0 35236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_363
timestamp 1623939100
transform 1 0 34500 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_372
timestamp 1623939100
transform 1 0 35328 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_384
timestamp 1623939100
transform 1 0 36432 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_396
timestamp 1623939100
transform 1 0 37536 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_408
timestamp 1623939100
transform 1 0 38640 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _785_
timestamp 1623939100
transform 1 0 40940 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_931
timestamp 1623939100
transform 1 0 40480 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_420
timestamp 1623939100
transform 1 0 39744 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_429
timestamp 1623939100
transform 1 0 40572 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_380
timestamp 1623939100
transform -1 0 43424 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_452
timestamp 1623939100
transform 1 0 42688 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _351_
timestamp 1623939100
transform -1 0 44252 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_42_469
timestamp 1623939100
transform 1 0 44252 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_932
timestamp 1623939100
transform 1 0 45724 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_481
timestamp 1623939100
transform 1 0 45356 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_486
timestamp 1623939100
transform 1 0 45816 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_498
timestamp 1623939100
transform 1 0 46920 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_510
timestamp 1623939100
transform 1 0 48024 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_522
timestamp 1623939100
transform 1 0 49128 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_534
timestamp 1623939100
transform 1 0 50232 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _342_
timestamp 1623939100
transform 1 0 52808 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _399_
timestamp 1623939100
transform 1 0 51612 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_933
timestamp 1623939100
transform 1 0 50968 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_543
timestamp 1623939100
transform 1 0 51060 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_558
timestamp 1623939100
transform 1 0 52440 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_568
timestamp 1623939100
transform 1 0 53360 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_580
timestamp 1623939100
transform 1 0 54464 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_934
timestamp 1623939100
transform 1 0 56212 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_592
timestamp 1623939100
transform 1 0 55568 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_598
timestamp 1623939100
transform 1 0 56120 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_600
timestamp 1623939100
transform 1 0 56304 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_612
timestamp 1623939100
transform 1 0 57408 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_624
timestamp 1623939100
transform 1 0 58512 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_636
timestamp 1623939100
transform 1 0 59616 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_935
timestamp 1623939100
transform 1 0 61456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_648
timestamp 1623939100
transform 1 0 60720 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_657
timestamp 1623939100
transform 1 0 61548 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_669
timestamp 1623939100
transform 1 0 62652 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_681
timestamp 1623939100
transform 1 0 63756 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_693
timestamp 1623939100
transform 1 0 64860 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_705
timestamp 1623939100
transform 1 0 65964 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_936
timestamp 1623939100
transform 1 0 66700 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_714
timestamp 1623939100
transform 1 0 66792 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_726
timestamp 1623939100
transform 1 0 67896 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_738
timestamp 1623939100
transform 1 0 69000 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_750
timestamp 1623939100
transform 1 0 70104 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_937
timestamp 1623939100
transform 1 0 71944 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_762
timestamp 1623939100
transform 1 0 71208 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  _528_
timestamp 1623939100
transform 1 0 73600 0 -1 25568
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_42_771
timestamp 1623939100
transform 1 0 72036 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_783
timestamp 1623939100
transform 1 0 73140 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_787
timestamp 1623939100
transform 1 0 73508 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_799
timestamp 1623939100
transform 1 0 74612 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_811
timestamp 1623939100
transform 1 0 75716 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_938
timestamp 1623939100
transform 1 0 77188 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_823
timestamp 1623939100
transform 1 0 76820 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_828
timestamp 1623939100
transform 1 0 77280 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_840
timestamp 1623939100
transform 1 0 78384 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_852
timestamp 1623939100
transform 1 0 79488 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_864
timestamp 1623939100
transform 1 0 80592 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_939
timestamp 1623939100
transform 1 0 82432 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_876
timestamp 1623939100
transform 1 0 81696 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_885
timestamp 1623939100
transform 1 0 82524 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_897
timestamp 1623939100
transform 1 0 83628 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_909
timestamp 1623939100
transform 1 0 84732 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_921
timestamp 1623939100
transform 1 0 85836 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_933
timestamp 1623939100
transform 1 0 86940 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_940
timestamp 1623939100
transform 1 0 87676 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_942
timestamp 1623939100
transform 1 0 87768 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_954
timestamp 1623939100
transform 1 0 88872 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _440_
timestamp 1623939100
transform 1 0 90620 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_94
timestamp 1623939100
transform 1 0 90436 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_96
timestamp 1623939100
transform 1 0 90252 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_98
timestamp 1623939100
transform 1 0 90068 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_966
timestamp 1623939100
transform 1 0 89976 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_941
timestamp 1623939100
transform 1 0 92920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_95
timestamp 1623939100
transform 1 0 92092 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_97
timestamp 1623939100
transform 1 0 92276 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_99
timestamp 1623939100
transform 1 0 92460 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_995
timestamp 1623939100
transform 1 0 92644 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_999
timestamp 1623939100
transform 1 0 93012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1011
timestamp 1623939100
transform 1 0 94116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1023
timestamp 1623939100
transform 1 0 95220 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1035
timestamp 1623939100
transform 1 0 96324 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1623939100
transform -1 0 98808 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_942
timestamp 1623939100
transform 1 0 98164 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_1047
timestamp 1623939100
transform 1 0 97428 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_1056
timestamp 1623939100
transform 1 0 98256 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1623939100
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1623939100
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1623939100
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1623939100
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1623939100
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_943
timestamp 1623939100
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_51
timestamp 1623939100
transform 1 0 5796 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_58
timestamp 1623939100
transform 1 0 6440 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_70
timestamp 1623939100
transform 1 0 7544 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_82
timestamp 1623939100
transform 1 0 8648 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_94
timestamp 1623939100
transform 1 0 9752 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_944
timestamp 1623939100
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_106
timestamp 1623939100
transform 1 0 10856 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_115
timestamp 1623939100
transform 1 0 11684 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_127
timestamp 1623939100
transform 1 0 12788 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_139
timestamp 1623939100
transform 1 0 13892 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_151
timestamp 1623939100
transform 1 0 14996 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_163
timestamp 1623939100
transform 1 0 16100 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_945
timestamp 1623939100
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_172
timestamp 1623939100
transform 1 0 16928 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_184
timestamp 1623939100
transform 1 0 18032 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _773_
timestamp 1623939100
transform 1 0 19044 0 1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_43_192
timestamp 1623939100
transform 1 0 18768 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_946
timestamp 1623939100
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_212
timestamp 1623939100
transform 1 0 20608 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_224
timestamp 1623939100
transform 1 0 21712 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_229
timestamp 1623939100
transform 1 0 22172 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _585_
timestamp 1623939100
transform 1 0 22724 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_238
timestamp 1623939100
transform 1 0 23000 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_250
timestamp 1623939100
transform 1 0 24104 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_262
timestamp 1623939100
transform 1 0 25208 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_947
timestamp 1623939100
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_274
timestamp 1623939100
transform 1 0 26312 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_282
timestamp 1623939100
transform 1 0 27048 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_286
timestamp 1623939100
transform 1 0 27416 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_298
timestamp 1623939100
transform 1 0 28520 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_310
timestamp 1623939100
transform 1 0 29624 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_322
timestamp 1623939100
transform 1 0 30728 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_948
timestamp 1623939100
transform 1 0 32568 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_334
timestamp 1623939100
transform 1 0 31832 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_343
timestamp 1623939100
transform 1 0 32660 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_355
timestamp 1623939100
transform 1 0 33764 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_367
timestamp 1623939100
transform 1 0 34868 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_379
timestamp 1623939100
transform 1 0 35972 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_391
timestamp 1623939100
transform 1 0 37076 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_4  _505_
timestamp 1623939100
transform 1 0 39192 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_949
timestamp 1623939100
transform 1 0 37812 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_400
timestamp 1623939100
transform 1 0 37904 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_412
timestamp 1623939100
transform 1 0 39008 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_430
timestamp 1623939100
transform 1 0 40664 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_950
timestamp 1623939100
transform 1 0 43056 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_442
timestamp 1623939100
transform 1 0 41768 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_454
timestamp 1623939100
transform 1 0 42872 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_457
timestamp 1623939100
transform 1 0 43148 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_469
timestamp 1623939100
transform 1 0 44252 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_481
timestamp 1623939100
transform 1 0 45356 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_493
timestamp 1623939100
transform 1 0 46460 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_951
timestamp 1623939100
transform 1 0 48300 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1623939100
transform 1 0 47564 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_514
timestamp 1623939100
transform 1 0 48392 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_526
timestamp 1623939100
transform 1 0 49496 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_538
timestamp 1623939100
transform 1 0 50600 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_550
timestamp 1623939100
transform 1 0 51704 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_562
timestamp 1623939100
transform 1 0 52808 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_952
timestamp 1623939100
transform 1 0 53544 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_571
timestamp 1623939100
transform 1 0 53636 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_583
timestamp 1623939100
transform 1 0 54740 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_595
timestamp 1623939100
transform 1 0 55844 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_607
timestamp 1623939100
transform 1 0 56948 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_619
timestamp 1623939100
transform 1 0 58052 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_953
timestamp 1623939100
transform 1 0 58788 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_628
timestamp 1623939100
transform 1 0 58880 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_640
timestamp 1623939100
transform 1 0 59984 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _605_
timestamp 1623939100
transform 1 0 61456 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_652
timestamp 1623939100
transform 1 0 61088 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_659
timestamp 1623939100
transform 1 0 61732 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_954
timestamp 1623939100
transform 1 0 64032 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_671
timestamp 1623939100
transform 1 0 62836 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_683
timestamp 1623939100
transform 1 0 63940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_685
timestamp 1623939100
transform 1 0 64124 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _653_
timestamp 1623939100
transform 1 0 66148 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_697
timestamp 1623939100
transform 1 0 65228 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_705
timestamp 1623939100
transform 1 0 65964 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _781_
timestamp 1623939100
transform 1 0 67160 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_43_710
timestamp 1623939100
transform 1 0 66424 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_955
timestamp 1623939100
transform 1 0 69276 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_737
timestamp 1623939100
transform 1 0 68908 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_742
timestamp 1623939100
transform 1 0 69368 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_754
timestamp 1623939100
transform 1 0 70472 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_766
timestamp 1623939100
transform 1 0 71576 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_778
timestamp 1623939100
transform 1 0 72680 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_790
timestamp 1623939100
transform 1 0 73784 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_956
timestamp 1623939100
transform 1 0 74520 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_799
timestamp 1623939100
transform 1 0 74612 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_811
timestamp 1623939100
transform 1 0 75716 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_823
timestamp 1623939100
transform 1 0 76820 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_835
timestamp 1623939100
transform 1 0 77924 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_847
timestamp 1623939100
transform 1 0 79028 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _652_
timestamp 1623939100
transform 1 0 80224 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_957
timestamp 1623939100
transform 1 0 79764 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_856
timestamp 1623939100
transform 1 0 79856 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_863
timestamp 1623939100
transform 1 0 80500 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_875
timestamp 1623939100
transform 1 0 81604 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_887
timestamp 1623939100
transform 1 0 82708 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_958
timestamp 1623939100
transform 1 0 85008 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_899
timestamp 1623939100
transform 1 0 83812 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_911
timestamp 1623939100
transform 1 0 84916 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_913
timestamp 1623939100
transform 1 0 85100 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_925
timestamp 1623939100
transform 1 0 86204 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_937
timestamp 1623939100
transform 1 0 87308 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_949
timestamp 1623939100
transform 1 0 88412 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_959
timestamp 1623939100
transform 1 0 90252 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_961
timestamp 1623939100
transform 1 0 89516 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_970
timestamp 1623939100
transform 1 0 90344 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_982
timestamp 1623939100
transform 1 0 91448 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_994
timestamp 1623939100
transform 1 0 92552 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1006
timestamp 1623939100
transform 1 0 93656 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_1018
timestamp 1623939100
transform 1 0 94760 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_960
timestamp 1623939100
transform 1 0 95496 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1027
timestamp 1623939100
transform 1 0 95588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1039
timestamp 1623939100
transform 1 0 96692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1623939100
transform -1 0 98808 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_1051
timestamp 1623939100
transform 1 0 97796 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1623939100
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1623939100
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1623939100
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _531_
timestamp 1623939100
transform 1 0 4692 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_961
timestamp 1623939100
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_199
timestamp 1623939100
transform 1 0 4508 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_27
timestamp 1623939100
transform 1 0 3588 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_30
timestamp 1623939100
transform 1 0 3864 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_36
timestamp 1623939100
transform 1 0 4416 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _593_
timestamp 1623939100
transform 1 0 6716 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_302
timestamp 1623939100
transform 1 0 6532 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_48
timestamp 1623939100
transform 1 0 5520 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_56
timestamp 1623939100
transform 1 0 6256 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_64
timestamp 1623939100
transform 1 0 6992 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_76
timestamp 1623939100
transform 1 0 8096 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_962
timestamp 1623939100
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_84
timestamp 1623939100
transform 1 0 8832 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_87
timestamp 1623939100
transform 1 0 9108 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_99
timestamp 1623939100
transform 1 0 10212 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_111
timestamp 1623939100
transform 1 0 11316 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_123
timestamp 1623939100
transform 1 0 12420 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_963
timestamp 1623939100
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_135
timestamp 1623939100
transform 1 0 13524 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_144
timestamp 1623939100
transform 1 0 14352 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _778_
timestamp 1623939100
transform 1 0 15088 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_44_171
timestamp 1623939100
transform 1 0 16836 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_183
timestamp 1623939100
transform 1 0 17940 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _309_
timestamp 1623939100
transform 1 0 19964 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_964
timestamp 1623939100
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_195
timestamp 1623939100
transform 1 0 19044 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_199
timestamp 1623939100
transform 1 0 19412 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_201
timestamp 1623939100
transform 1 0 19596 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_214
timestamp 1623939100
transform 1 0 20792 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_226
timestamp 1623939100
transform 1 0 21896 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_238
timestamp 1623939100
transform 1 0 23000 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_250
timestamp 1623939100
transform 1 0 24104 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_965
timestamp 1623939100
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_256
timestamp 1623939100
transform 1 0 24656 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_258
timestamp 1623939100
transform 1 0 24840 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_270
timestamp 1623939100
transform 1 0 25944 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_282
timestamp 1623939100
transform 1 0 27048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_294
timestamp 1623939100
transform 1 0 28152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_306
timestamp 1623939100
transform 1 0 29256 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _389_
timestamp 1623939100
transform -1 0 31004 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_966
timestamp 1623939100
transform 1 0 29992 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_146
timestamp 1623939100
transform -1 0 30452 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_315
timestamp 1623939100
transform 1 0 30084 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_325
timestamp 1623939100
transform 1 0 31004 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_337
timestamp 1623939100
transform 1 0 32108 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_349
timestamp 1623939100
transform 1 0 33212 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_967
timestamp 1623939100
transform 1 0 35236 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_150
timestamp 1623939100
transform 1 0 35512 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_361
timestamp 1623939100
transform 1 0 34316 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_369
timestamp 1623939100
transform 1 0 35052 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_372
timestamp 1623939100
transform 1 0 35328 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _412_
timestamp 1623939100
transform 1 0 35696 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_44_385
timestamp 1623939100
transform 1 0 36524 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_397
timestamp 1623939100
transform 1 0 37628 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_409
timestamp 1623939100
transform 1 0 38732 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_968
timestamp 1623939100
transform 1 0 40480 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_421
timestamp 1623939100
transform 1 0 39836 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_427
timestamp 1623939100
transform 1 0 40388 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_429
timestamp 1623939100
transform 1 0 40572 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_441
timestamp 1623939100
transform 1 0 41676 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_453
timestamp 1623939100
transform 1 0 42780 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_465
timestamp 1623939100
transform 1 0 43884 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_477
timestamp 1623939100
transform 1 0 44988 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_969
timestamp 1623939100
transform 1 0 45724 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_486
timestamp 1623939100
transform 1 0 45816 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_498
timestamp 1623939100
transform 1 0 46920 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_4  _391_
timestamp 1623939100
transform 1 0 47840 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_44_506
timestamp 1623939100
transform 1 0 47656 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _307_
timestamp 1623939100
transform 1 0 49956 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_44_524
timestamp 1623939100
transform 1 0 49312 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_530
timestamp 1623939100
transform 1 0 49864 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_538
timestamp 1623939100
transform 1 0 50600 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_970
timestamp 1623939100
transform 1 0 50968 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_543
timestamp 1623939100
transform 1 0 51060 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_555
timestamp 1623939100
transform 1 0 52164 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_567
timestamp 1623939100
transform 1 0 53268 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_579
timestamp 1623939100
transform 1 0 54372 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_971
timestamp 1623939100
transform 1 0 56212 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_591
timestamp 1623939100
transform 1 0 55476 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_600
timestamp 1623939100
transform 1 0 56304 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_612
timestamp 1623939100
transform 1 0 57408 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_624
timestamp 1623939100
transform 1 0 58512 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_636
timestamp 1623939100
transform 1 0 59616 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_972
timestamp 1623939100
transform 1 0 61456 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_648
timestamp 1623939100
transform 1 0 60720 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_657
timestamp 1623939100
transform 1 0 61548 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_669
timestamp 1623939100
transform 1 0 62652 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_681
timestamp 1623939100
transform 1 0 63756 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_693
timestamp 1623939100
transform 1 0 64860 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_705
timestamp 1623939100
transform 1 0 65964 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_973
timestamp 1623939100
transform 1 0 66700 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_714
timestamp 1623939100
transform 1 0 66792 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_726
timestamp 1623939100
transform 1 0 67896 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_738
timestamp 1623939100
transform 1 0 69000 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_750
timestamp 1623939100
transform 1 0 70104 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_974
timestamp 1623939100
transform 1 0 71944 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_762
timestamp 1623939100
transform 1 0 71208 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _324_
timestamp 1623939100
transform 1 0 73324 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_44_771
timestamp 1623939100
transform 1 0 72036 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_783
timestamp 1623939100
transform 1 0 73140 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_794
timestamp 1623939100
transform 1 0 74152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_806
timestamp 1623939100
transform 1 0 75256 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_975
timestamp 1623939100
transform 1 0 77188 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_818
timestamp 1623939100
transform 1 0 76360 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_826
timestamp 1623939100
transform 1 0 77096 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_828
timestamp 1623939100
transform 1 0 77280 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_840
timestamp 1623939100
transform 1 0 78384 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_852
timestamp 1623939100
transform 1 0 79488 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_864
timestamp 1623939100
transform 1 0 80592 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_976
timestamp 1623939100
transform 1 0 82432 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_876
timestamp 1623939100
transform 1 0 81696 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_885
timestamp 1623939100
transform 1 0 82524 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_897
timestamp 1623939100
transform 1 0 83628 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_909
timestamp 1623939100
transform 1 0 84732 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _534_
timestamp 1623939100
transform -1 0 87032 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_226
timestamp 1623939100
transform -1 0 86204 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_921
timestamp 1623939100
transform 1 0 85836 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_934
timestamp 1623939100
transform 1 0 87032 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _578_
timestamp 1623939100
transform -1 0 88412 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_977
timestamp 1623939100
transform 1 0 87676 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_272
timestamp 1623939100
transform -1 0 88136 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_940
timestamp 1623939100
transform 1 0 87584 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_942
timestamp 1623939100
transform 1 0 87768 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_949
timestamp 1623939100
transform 1 0 88412 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_4  _407_
timestamp 1623939100
transform 1 0 90620 0 -1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA_184
timestamp 1623939100
transform 1 0 90436 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_961
timestamp 1623939100
transform 1 0 89516 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_969
timestamp 1623939100
transform 1 0 90252 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_978
timestamp 1623939100
transform 1 0 92920 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_987
timestamp 1623939100
transform 1 0 91908 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_995
timestamp 1623939100
transform 1 0 92644 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_999
timestamp 1623939100
transform 1 0 93012 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1011
timestamp 1623939100
transform 1 0 94116 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1023
timestamp 1623939100
transform 1 0 95220 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1035
timestamp 1623939100
transform 1 0 96324 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1623939100
transform -1 0 98808 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_979
timestamp 1623939100
transform 1 0 98164 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_1047
timestamp 1623939100
transform 1 0 97428 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_1056
timestamp 1623939100
transform 1 0 98256 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1623939100
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1623939100
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1623939100
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1623939100
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1623939100
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_980
timestamp 1623939100
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_51
timestamp 1623939100
transform 1 0 5796 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_58
timestamp 1623939100
transform 1 0 6440 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_70
timestamp 1623939100
transform 1 0 7544 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_82
timestamp 1623939100
transform 1 0 8648 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_94
timestamp 1623939100
transform 1 0 9752 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_981
timestamp 1623939100
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_106
timestamp 1623939100
transform 1 0 10856 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_115
timestamp 1623939100
transform 1 0 11684 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_127
timestamp 1623939100
transform 1 0 12788 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_139
timestamp 1623939100
transform 1 0 13892 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_151
timestamp 1623939100
transform 1 0 14996 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_163
timestamp 1623939100
transform 1 0 16100 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_982
timestamp 1623939100
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_172
timestamp 1623939100
transform 1 0 16928 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1623939100
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1623939100
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1623939100
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_983
timestamp 1623939100
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_220
timestamp 1623939100
transform 1 0 21344 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_229
timestamp 1623939100
transform 1 0 22172 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_241
timestamp 1623939100
transform 1 0 23276 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1623939100
transform 1 0 24380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_265
timestamp 1623939100
transform 1 0 25484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_984
timestamp 1623939100
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_277
timestamp 1623939100
transform 1 0 26588 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_286
timestamp 1623939100
transform 1 0 27416 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_298
timestamp 1623939100
transform 1 0 28520 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_310
timestamp 1623939100
transform 1 0 29624 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_322
timestamp 1623939100
transform 1 0 30728 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_985
timestamp 1623939100
transform 1 0 32568 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_334
timestamp 1623939100
transform 1 0 31832 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_343
timestamp 1623939100
transform 1 0 32660 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_355
timestamp 1623939100
transform 1 0 33764 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_367
timestamp 1623939100
transform 1 0 34868 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_379
timestamp 1623939100
transform 1 0 35972 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_391
timestamp 1623939100
transform 1 0 37076 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _395_
timestamp 1623939100
transform 1 0 39192 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_986
timestamp 1623939100
transform 1 0 37812 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_400
timestamp 1623939100
transform 1 0 37904 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_412
timestamp 1623939100
transform 1 0 39008 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_423
timestamp 1623939100
transform 1 0 40020 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_435
timestamp 1623939100
transform 1 0 41124 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_987
timestamp 1623939100
transform 1 0 43056 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_447
timestamp 1623939100
transform 1 0 42228 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_455
timestamp 1623939100
transform 1 0 42964 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_457
timestamp 1623939100
transform 1 0 43148 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_469
timestamp 1623939100
transform 1 0 44252 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_481
timestamp 1623939100
transform 1 0 45356 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_493
timestamp 1623939100
transform 1 0 46460 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_988
timestamp 1623939100
transform 1 0 48300 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1623939100
transform 1 0 47564 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_514
timestamp 1623939100
transform 1 0 48392 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_526
timestamp 1623939100
transform 1 0 49496 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_538
timestamp 1623939100
transform 1 0 50600 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_550
timestamp 1623939100
transform 1 0 51704 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_562
timestamp 1623939100
transform 1 0 52808 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_989
timestamp 1623939100
transform 1 0 53544 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_571
timestamp 1623939100
transform 1 0 53636 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_583
timestamp 1623939100
transform 1 0 54740 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_595
timestamp 1623939100
transform 1 0 55844 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_607
timestamp 1623939100
transform 1 0 56948 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_619
timestamp 1623939100
transform 1 0 58052 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _726_
timestamp 1623939100
transform 1 0 59616 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_990
timestamp 1623939100
transform 1 0 58788 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_628
timestamp 1623939100
transform 1 0 58880 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_655
timestamp 1623939100
transform 1 0 61364 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_991
timestamp 1623939100
transform 1 0 64032 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_667
timestamp 1623939100
transform 1 0 62468 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_679
timestamp 1623939100
transform 1 0 63572 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_683
timestamp 1623939100
transform 1 0 63940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_685
timestamp 1623939100
transform 1 0 64124 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_697
timestamp 1623939100
transform 1 0 65228 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_709
timestamp 1623939100
transform 1 0 66332 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_721
timestamp 1623939100
transform 1 0 67436 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_992
timestamp 1623939100
transform 1 0 69276 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_733
timestamp 1623939100
transform 1 0 68540 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_742
timestamp 1623939100
transform 1 0 69368 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_754
timestamp 1623939100
transform 1 0 70472 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_766
timestamp 1623939100
transform 1 0 71576 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_778
timestamp 1623939100
transform 1 0 72680 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_790
timestamp 1623939100
transform 1 0 73784 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_993
timestamp 1623939100
transform 1 0 74520 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_799
timestamp 1623939100
transform 1 0 74612 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_811
timestamp 1623939100
transform 1 0 75716 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_823
timestamp 1623939100
transform 1 0 76820 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_831
timestamp 1623939100
transform 1 0 77556 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _546_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 78016 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA_175
timestamp 1623939100
transform 1 0 77832 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_177
timestamp 1623939100
transform 1 0 78476 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_843
timestamp 1623939100
transform 1 0 78660 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_994
timestamp 1623939100
transform 1 0 79764 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_856
timestamp 1623939100
transform 1 0 79856 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_868
timestamp 1623939100
transform 1 0 80960 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_880
timestamp 1623939100
transform 1 0 82064 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_892
timestamp 1623939100
transform 1 0 83168 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_995
timestamp 1623939100
transform 1 0 85008 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_904
timestamp 1623939100
transform 1 0 84272 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_913
timestamp 1623939100
transform 1 0 85100 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _705_
timestamp 1623939100
transform 1 0 86296 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_45_925
timestamp 1623939100
transform 1 0 86204 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_945
timestamp 1623939100
transform 1 0 88044 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_957
timestamp 1623939100
transform 1 0 89148 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_996
timestamp 1623939100
transform 1 0 90252 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_970
timestamp 1623939100
transform 1 0 90344 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_982
timestamp 1623939100
transform 1 0 91448 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_994
timestamp 1623939100
transform 1 0 92552 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _298_
timestamp 1623939100
transform 1 0 94208 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1006
timestamp 1623939100
transform 1 0 93656 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1019
timestamp 1623939100
transform 1 0 94852 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_4  _478_
timestamp 1623939100
transform 1 0 96692 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_997
timestamp 1623939100
transform 1 0 95496 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1025
timestamp 1623939100
transform 1 0 95404 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1027
timestamp 1623939100
transform 1 0 95588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1623939100
transform -1 0 98808 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1055
timestamp 1623939100
transform 1 0 98164 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1623939100
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1623939100
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1623939100
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1623939100
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1623939100
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_15
timestamp 1623939100
transform 1 0 2484 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _311_
timestamp 1623939100
transform 1 0 3588 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_998
timestamp 1623939100
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_208
timestamp 1623939100
transform 1 0 3404 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_27
timestamp 1623939100
transform 1 0 3588 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_30
timestamp 1623939100
transform 1 0 3864 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_23
timestamp 1623939100
transform 1 0 3220 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_33
timestamp 1623939100
transform 1 0 4140 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1017
timestamp 1623939100
transform 1 0 6348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_42
timestamp 1623939100
transform 1 0 4968 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_54
timestamp 1623939100
transform 1 0 6072 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_45
timestamp 1623939100
transform 1 0 5244 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_58
timestamp 1623939100
transform 1 0 6440 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_66
timestamp 1623939100
transform 1 0 7176 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_78
timestamp 1623939100
transform 1 0 8280 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_70
timestamp 1623939100
transform 1 0 7544 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_82
timestamp 1623939100
transform 1 0 8648 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_999
timestamp 1623939100
transform 1 0 9016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_87
timestamp 1623939100
transform 1 0 9108 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_99
timestamp 1623939100
transform 1 0 10212 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_94
timestamp 1623939100
transform 1 0 9752 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4_2  _295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 10948 0 -1 27744
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _506_
timestamp 1623939100
transform 1 0 12236 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1018
timestamp 1623939100
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_117
timestamp 1623939100
transform 1 0 11868 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_106
timestamp 1623939100
transform 1 0 10856 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_115
timestamp 1623939100
transform 1 0 11684 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_2  _419_
timestamp 1623939100
transform -1 0 14628 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1000
timestamp 1623939100
transform 1 0 14260 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_205
timestamp 1623939100
transform -1 0 13984 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_130
timestamp 1623939100
transform 1 0 13064 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_142
timestamp 1623939100
transform 1 0 14168 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_144
timestamp 1623939100
transform 1 0 14352 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_127
timestamp 1623939100
transform 1 0 12788 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_135
timestamp 1623939100
transform 1 0 13524 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _592_
timestamp 1623939100
transform 1 0 15088 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _699_
timestamp 1623939100
transform 1 0 15824 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_300
timestamp 1623939100
transform 1 0 14904 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_155
timestamp 1623939100
transform 1 0 15364 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_159
timestamp 1623939100
transform 1 0 15732 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_147
timestamp 1623939100
transform 1 0 14628 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_159
timestamp 1623939100
transform 1 0 15732 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _702_
timestamp 1623939100
transform -1 0 19044 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1019
timestamp 1623939100
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1623939100
transform -1 0 17296 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1623939100
transform -1 0 17112 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_179
timestamp 1623939100
transform 1 0 17572 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _536_
timestamp 1623939100
transform 1 0 19780 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1001
timestamp 1623939100
transform 1 0 19504 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1623939100
transform -1 0 19228 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_191
timestamp 1623939100
transform 1 0 18676 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_199
timestamp 1623939100
transform 1 0 19412 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_201
timestamp 1623939100
transform 1 0 19596 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_197
timestamp 1623939100
transform 1 0 19228 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1020
timestamp 1623939100
transform 1 0 22080 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_213
timestamp 1623939100
transform 1 0 20700 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1623939100
transform 1 0 21804 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_212
timestamp 1623939100
transform 1 0 20608 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_224
timestamp 1623939100
transform 1 0 21712 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_229
timestamp 1623939100
transform 1 0 22172 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _642_
timestamp 1623939100
transform 1 0 23460 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_237
timestamp 1623939100
transform 1 0 22908 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_246
timestamp 1623939100
transform 1 0 23736 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_241
timestamp 1623939100
transform 1 0 23276 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1002
timestamp 1623939100
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_254
timestamp 1623939100
transform 1 0 24472 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_258
timestamp 1623939100
transform 1 0 24840 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_270
timestamp 1623939100
transform 1 0 25944 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_253
timestamp 1623939100
transform 1 0 24380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_265
timestamp 1623939100
transform 1 0 25484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _782_
timestamp 1623939100
transform 1 0 27508 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1021
timestamp 1623939100
transform 1 0 27324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_282
timestamp 1623939100
transform 1 0 27048 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_286
timestamp 1623939100
transform 1 0 27416 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_277
timestamp 1623939100
transform 1 0 26588 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_286
timestamp 1623939100
transform 1 0 27416 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_306
timestamp 1623939100
transform 1 0 29256 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_298
timestamp 1623939100
transform 1 0 28520 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_310
timestamp 1623939100
transform 1 0 29624 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1003
timestamp 1623939100
transform 1 0 29992 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_315
timestamp 1623939100
transform 1 0 30084 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_327
timestamp 1623939100
transform 1 0 31188 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_322
timestamp 1623939100
transform 1 0 30728 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _483_
timestamp 1623939100
transform 1 0 33028 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1022
timestamp 1623939100
transform 1 0 32568 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_339
timestamp 1623939100
transform 1 0 32292 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_351
timestamp 1623939100
transform 1 0 33396 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_334
timestamp 1623939100
transform 1 0 31832 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_343
timestamp 1623939100
transform 1 0 32660 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1004
timestamp 1623939100
transform 1 0 35236 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_363
timestamp 1623939100
transform 1 0 34500 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_372
timestamp 1623939100
transform 1 0 35328 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_356
timestamp 1623939100
transform 1 0 33856 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_368
timestamp 1623939100
transform 1 0 34960 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_384
timestamp 1623939100
transform 1 0 36432 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_380
timestamp 1623939100
transform 1 0 36064 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_392
timestamp 1623939100
transform 1 0 37168 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_400
timestamp 1623939100
transform 1 0 37904 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_398
timestamp 1623939100
transform 1 0 37720 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1023
timestamp 1623939100
transform 1 0 37812 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_408
timestamp 1623939100
transform 1 0 38640 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_408
timestamp 1623939100
transform 1 0 38640 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_329
timestamp 1623939100
transform 1 0 38824 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _627_
timestamp 1623939100
transform 1 0 39008 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _529_
timestamp 1623939100
transform 1 0 38916 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_47_415
timestamp 1623939100
transform 1 0 39284 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_396
timestamp 1623939100
transform 1 0 37536 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _330_
timestamp 1623939100
transform -1 0 42136 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1005
timestamp 1623939100
transform 1 0 40480 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_383
timestamp 1623939100
transform -1 0 41308 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_420
timestamp 1623939100
transform 1 0 39744 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_429
timestamp 1623939100
transform 1 0 40572 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_427
timestamp 1623939100
transform 1 0 40388 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1024
timestamp 1623939100
transform 1 0 43056 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_446
timestamp 1623939100
transform 1 0 42136 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_458
timestamp 1623939100
transform 1 0 43240 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_439
timestamp 1623939100
transform 1 0 41492 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_451
timestamp 1623939100
transform 1 0 42596 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_455
timestamp 1623939100
transform 1 0 42964 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_457
timestamp 1623939100
transform 1 0 43148 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_470
timestamp 1623939100
transform 1 0 44344 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_469
timestamp 1623939100
transform 1 0 44252 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1006
timestamp 1623939100
transform 1 0 45724 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_482
timestamp 1623939100
transform 1 0 45448 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_486
timestamp 1623939100
transform 1 0 45816 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_498
timestamp 1623939100
transform 1 0 46920 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_481
timestamp 1623939100
transform 1 0 45356 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_493
timestamp 1623939100
transform 1 0 46460 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1025
timestamp 1623939100
transform 1 0 48300 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_510
timestamp 1623939100
transform 1 0 48024 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1623939100
transform 1 0 47564 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_514
timestamp 1623939100
transform 1 0 48392 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_522
timestamp 1623939100
transform 1 0 49128 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_534
timestamp 1623939100
transform 1 0 50232 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_526
timestamp 1623939100
transform 1 0 49496 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_538
timestamp 1623939100
transform 1 0 50600 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1007
timestamp 1623939100
transform 1 0 50968 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_543
timestamp 1623939100
transform 1 0 51060 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_555
timestamp 1623939100
transform 1 0 52164 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_550
timestamp 1623939100
transform 1 0 51704 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_562
timestamp 1623939100
transform 1 0 52808 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _361_
timestamp 1623939100
transform 1 0 53176 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1026
timestamp 1623939100
transform 1 0 53544 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_563
timestamp 1623939100
transform 1 0 52900 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_575
timestamp 1623939100
transform 1 0 54004 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_571
timestamp 1623939100
transform 1 0 53636 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_583
timestamp 1623939100
transform 1 0 54740 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1008
timestamp 1623939100
transform 1 0 56212 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_587
timestamp 1623939100
transform 1 0 55108 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_600
timestamp 1623939100
transform 1 0 56304 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_595
timestamp 1623939100
transform 1 0 55844 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_612
timestamp 1623939100
transform 1 0 57408 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_624
timestamp 1623939100
transform 1 0 58512 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_607
timestamp 1623939100
transform 1 0 56948 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_619
timestamp 1623939100
transform 1 0 58052 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1027
timestamp 1623939100
transform 1 0 58788 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_636
timestamp 1623939100
transform 1 0 59616 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_628
timestamp 1623939100
transform 1 0 58880 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_640
timestamp 1623939100
transform 1 0 59984 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1009
timestamp 1623939100
transform 1 0 61456 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_648
timestamp 1623939100
transform 1 0 60720 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_657
timestamp 1623939100
transform 1 0 61548 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_652
timestamp 1623939100
transform 1 0 61088 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_664
timestamp 1623939100
transform 1 0 62192 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1028
timestamp 1623939100
transform 1 0 64032 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_669
timestamp 1623939100
transform 1 0 62652 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_681
timestamp 1623939100
transform 1 0 63756 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_676
timestamp 1623939100
transform 1 0 63296 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_685
timestamp 1623939100
transform 1 0 64124 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_693
timestamp 1623939100
transform 1 0 64860 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_705
timestamp 1623939100
transform 1 0 65964 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_697
timestamp 1623939100
transform 1 0 65228 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1010
timestamp 1623939100
transform 1 0 66700 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_714
timestamp 1623939100
transform 1 0 66792 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_726
timestamp 1623939100
transform 1 0 67896 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_709
timestamp 1623939100
transform 1 0 66332 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_721
timestamp 1623939100
transform 1 0 67436 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1029
timestamp 1623939100
transform 1 0 69276 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_738
timestamp 1623939100
transform 1 0 69000 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_750
timestamp 1623939100
transform 1 0 70104 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_733
timestamp 1623939100
transform 1 0 68540 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_742
timestamp 1623939100
transform 1 0 69368 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1011
timestamp 1623939100
transform 1 0 71944 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_762
timestamp 1623939100
transform 1 0 71208 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_754
timestamp 1623939100
transform 1 0 70472 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_766
timestamp 1623939100
transform 1 0 71576 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_771
timestamp 1623939100
transform 1 0 72036 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_783
timestamp 1623939100
transform 1 0 73140 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_778
timestamp 1623939100
transform 1 0 72680 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_790
timestamp 1623939100
transform 1 0 73784 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1030
timestamp 1623939100
transform 1 0 74520 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_795
timestamp 1623939100
transform 1 0 74244 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_807
timestamp 1623939100
transform 1 0 75348 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_799
timestamp 1623939100
transform 1 0 74612 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_811
timestamp 1623939100
transform 1 0 75716 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1012
timestamp 1623939100
transform 1 0 77188 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_819
timestamp 1623939100
transform 1 0 76452 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_828
timestamp 1623939100
transform 1 0 77280 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_823
timestamp 1623939100
transform 1 0 76820 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _738_
timestamp 1623939100
transform 1 0 79304 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_46_840
timestamp 1623939100
transform 1 0 78384 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_848
timestamp 1623939100
transform 1 0 79120 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_835
timestamp 1623939100
transform 1 0 77924 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_847
timestamp 1623939100
transform 1 0 79028 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1031
timestamp 1623939100
transform 1 0 79764 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_869
timestamp 1623939100
transform 1 0 81052 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_856
timestamp 1623939100
transform 1 0 79856 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_868
timestamp 1623939100
transform 1 0 80960 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1013
timestamp 1623939100
transform 1 0 82432 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_881
timestamp 1623939100
transform 1 0 82156 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_885
timestamp 1623939100
transform 1 0 82524 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_880
timestamp 1623939100
transform 1 0 82064 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_892
timestamp 1623939100
transform 1 0 83168 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1032
timestamp 1623939100
transform 1 0 85008 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_897
timestamp 1623939100
transform 1 0 83628 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_909
timestamp 1623939100
transform 1 0 84732 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_904
timestamp 1623939100
transform 1 0 84272 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_913
timestamp 1623939100
transform 1 0 85100 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _516_
timestamp 1623939100
transform -1 0 87860 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_229
timestamp 1623939100
transform -1 0 87032 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_921
timestamp 1623939100
transform 1 0 85836 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_933
timestamp 1623939100
transform 1 0 86940 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_925
timestamp 1623939100
transform 1 0 86204 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_931
timestamp 1623939100
transform 1 0 86756 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1014
timestamp 1623939100
transform 1 0 87676 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_942
timestamp 1623939100
transform 1 0 87768 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_954
timestamp 1623939100
transform 1 0 88872 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_943
timestamp 1623939100
transform 1 0 87860 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_955
timestamp 1623939100
transform 1 0 88964 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1033
timestamp 1623939100
transform 1 0 90252 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_966
timestamp 1623939100
transform 1 0 89976 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_978
timestamp 1623939100
transform 1 0 91080 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_967
timestamp 1623939100
transform 1 0 90068 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_970
timestamp 1623939100
transform 1 0 90344 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1015
timestamp 1623939100
transform 1 0 92920 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_990
timestamp 1623939100
transform 1 0 92184 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_999
timestamp 1623939100
transform 1 0 93012 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_982
timestamp 1623939100
transform 1 0 91448 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_994
timestamp 1623939100
transform 1 0 92552 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1011
timestamp 1623939100
transform 1 0 94116 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1006
timestamp 1623939100
transform 1 0 93656 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_1018
timestamp 1623939100
transform 1 0 94760 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1034
timestamp 1623939100
transform 1 0 95496 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1023
timestamp 1623939100
transform 1 0 95220 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1035
timestamp 1623939100
transform 1 0 96324 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1027
timestamp 1623939100
transform 1 0 95588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1039
timestamp 1623939100
transform 1 0 96692 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1623939100
transform -1 0 98808 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1623939100
transform -1 0 98808 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1016
timestamp 1623939100
transform 1 0 98164 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1047
timestamp 1623939100
transform 1 0 97428 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_1056
timestamp 1623939100
transform 1 0 98256 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_1051
timestamp 1623939100
transform 1 0 97796 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _780_
timestamp 1623939100
transform 1 0 1656 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1623939100
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_3
timestamp 1623939100
transform 1 0 1380 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1035
timestamp 1623939100
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_25
timestamp 1623939100
transform 1 0 3404 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_30
timestamp 1623939100
transform 1 0 3864 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _572_
timestamp 1623939100
transform 1 0 5520 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_321
timestamp 1623939100
transform 1 0 5336 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_42
timestamp 1623939100
transform 1 0 4968 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_51
timestamp 1623939100
transform 1 0 5796 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_63
timestamp 1623939100
transform 1 0 6900 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_75
timestamp 1623939100
transform 1 0 8004 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_83
timestamp 1623939100
transform 1 0 8740 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1036
timestamp 1623939100
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_87
timestamp 1623939100
transform 1 0 9108 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_99
timestamp 1623939100
transform 1 0 10212 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_111
timestamp 1623939100
transform 1 0 11316 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_123
timestamp 1623939100
transform 1 0 12420 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1037
timestamp 1623939100
transform 1 0 14260 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_135
timestamp 1623939100
transform 1 0 13524 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_144
timestamp 1623939100
transform 1 0 14352 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _755_
timestamp 1623939100
transform 1 0 15640 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_100
timestamp 1623939100
transform 1 0 15456 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_102
timestamp 1623939100
transform 1 0 15272 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_104
timestamp 1623939100
transform 1 0 15088 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_101
timestamp 1623939100
transform 1 0 17388 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_103
timestamp 1623939100
transform 1 0 17572 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_105
timestamp 1623939100
transform 1 0 17756 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_183
timestamp 1623939100
transform 1 0 17940 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1038
timestamp 1623939100
transform 1 0 19504 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_195
timestamp 1623939100
transform 1 0 19044 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_199
timestamp 1623939100
transform 1 0 19412 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_201
timestamp 1623939100
transform 1 0 19596 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _462_
timestamp 1623939100
transform 1 0 20700 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_48_222
timestamp 1623939100
transform 1 0 21528 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_234
timestamp 1623939100
transform 1 0 22632 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_246
timestamp 1623939100
transform 1 0 23736 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1039
timestamp 1623939100
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_254
timestamp 1623939100
transform 1 0 24472 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_258
timestamp 1623939100
transform 1 0 24840 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_270
timestamp 1623939100
transform 1 0 25944 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_282
timestamp 1623939100
transform 1 0 27048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_294
timestamp 1623939100
transform 1 0 28152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_306
timestamp 1623939100
transform 1 0 29256 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1040
timestamp 1623939100
transform 1 0 29992 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_315
timestamp 1623939100
transform 1 0 30084 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_327
timestamp 1623939100
transform 1 0 31188 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _360_
timestamp 1623939100
transform 1 0 33304 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_231
timestamp 1623939100
transform 1 0 33120 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_339
timestamp 1623939100
transform 1 0 32292 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_347
timestamp 1623939100
transform 1 0 33028 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1041
timestamp 1623939100
transform 1 0 35236 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_357
timestamp 1623939100
transform 1 0 33948 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_369
timestamp 1623939100
transform 1 0 35052 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_372
timestamp 1623939100
transform 1 0 35328 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _290_
timestamp 1623939100
transform -1 0 37812 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_211
timestamp 1623939100
transform -1 0 37260 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_384
timestamp 1623939100
transform 1 0 36432 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_390
timestamp 1623939100
transform 1 0 36984 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_399
timestamp 1623939100
transform 1 0 37812 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_411
timestamp 1623939100
transform 1 0 38916 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1042
timestamp 1623939100
transform 1 0 40480 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_423
timestamp 1623939100
transform 1 0 40020 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_427
timestamp 1623939100
transform 1 0 40388 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_429
timestamp 1623939100
transform 1 0 40572 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_441
timestamp 1623939100
transform 1 0 41676 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_453
timestamp 1623939100
transform 1 0 42780 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_465
timestamp 1623939100
transform 1 0 43884 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_477
timestamp 1623939100
transform 1 0 44988 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1043
timestamp 1623939100
transform 1 0 45724 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_486
timestamp 1623939100
transform 1 0 45816 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_498
timestamp 1623939100
transform 1 0 46920 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _701_
timestamp 1623939100
transform -1 0 49496 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1623939100
transform -1 0 47748 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_504
timestamp 1623939100
transform 1 0 47472 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_526
timestamp 1623939100
transform 1 0 49496 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_538
timestamp 1623939100
transform 1 0 50600 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1044
timestamp 1623939100
transform 1 0 50968 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_543
timestamp 1623939100
transform 1 0 51060 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_555
timestamp 1623939100
transform 1 0 52164 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_567
timestamp 1623939100
transform 1 0 53268 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_579
timestamp 1623939100
transform 1 0 54372 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1045
timestamp 1623939100
transform 1 0 56212 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_591
timestamp 1623939100
transform 1 0 55476 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_600
timestamp 1623939100
transform 1 0 56304 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_612
timestamp 1623939100
transform 1 0 57408 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_624
timestamp 1623939100
transform 1 0 58512 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_636
timestamp 1623939100
transform 1 0 59616 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1046
timestamp 1623939100
transform 1 0 61456 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_wb_clk_i
timestamp 1623939100
transform 1 0 61916 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_648
timestamp 1623939100
transform 1 0 60720 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_657
timestamp 1623939100
transform 1 0 61548 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_664
timestamp 1623939100
transform 1 0 62192 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_676
timestamp 1623939100
transform 1 0 63296 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_688
timestamp 1623939100
transform 1 0 64400 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_700
timestamp 1623939100
transform 1 0 65504 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1047
timestamp 1623939100
transform 1 0 66700 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_712
timestamp 1623939100
transform 1 0 66608 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_714
timestamp 1623939100
transform 1 0 66792 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_726
timestamp 1623939100
transform 1 0 67896 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_738
timestamp 1623939100
transform 1 0 69000 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_750
timestamp 1623939100
transform 1 0 70104 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1048
timestamp 1623939100
transform 1 0 71944 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_762
timestamp 1623939100
transform 1 0 71208 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_771
timestamp 1623939100
transform 1 0 72036 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_783
timestamp 1623939100
transform 1 0 73140 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_795
timestamp 1623939100
transform 1 0 74244 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_807
timestamp 1623939100
transform 1 0 75348 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1049
timestamp 1623939100
transform 1 0 77188 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_819
timestamp 1623939100
transform 1 0 76452 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_828
timestamp 1623939100
transform 1 0 77280 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _499_
timestamp 1623939100
transform -1 0 79028 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_196
timestamp 1623939100
transform -1 0 78200 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_847
timestamp 1623939100
transform 1 0 79028 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_wb_clk_i
timestamp 1623939100
transform 1 0 80868 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_859
timestamp 1623939100
transform 1 0 80132 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_870
timestamp 1623939100
transform 1 0 81144 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1050
timestamp 1623939100
transform 1 0 82432 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_882
timestamp 1623939100
transform 1 0 82248 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_885
timestamp 1623939100
transform 1 0 82524 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_897
timestamp 1623939100
transform 1 0 83628 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_909
timestamp 1623939100
transform 1 0 84732 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_921
timestamp 1623939100
transform 1 0 85836 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_933
timestamp 1623939100
transform 1 0 86940 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1051
timestamp 1623939100
transform 1 0 87676 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_942
timestamp 1623939100
transform 1 0 87768 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_954
timestamp 1623939100
transform 1 0 88872 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_966
timestamp 1623939100
transform 1 0 89976 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_978
timestamp 1623939100
transform 1 0 91080 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1052
timestamp 1623939100
transform 1 0 92920 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_990
timestamp 1623939100
transform 1 0 92184 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_999
timestamp 1623939100
transform 1 0 93012 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1011
timestamp 1623939100
transform 1 0 94116 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1023
timestamp 1623939100
transform 1 0 95220 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1035
timestamp 1623939100
transform 1 0 96324 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1623939100
transform -1 0 98808 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1053
timestamp 1623939100
transform 1 0 98164 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_1047
timestamp 1623939100
transform 1 0 97428 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_1056
timestamp 1623939100
transform 1 0 98256 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1623939100
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1623939100
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1623939100
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1623939100
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1623939100
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1054
timestamp 1623939100
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_51
timestamp 1623939100
transform 1 0 5796 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_58
timestamp 1623939100
transform 1 0 6440 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _725_
timestamp 1623939100
transform 1 0 8096 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_49_70
timestamp 1623939100
transform 1 0 7544 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_95
timestamp 1623939100
transform 1 0 9844 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1055
timestamp 1623939100
transform 1 0 11592 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_107
timestamp 1623939100
transform 1 0 10948 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_113
timestamp 1623939100
transform 1 0 11500 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_115
timestamp 1623939100
transform 1 0 11684 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _520_
timestamp 1623939100
transform 1 0 13892 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_49_127
timestamp 1623939100
transform 1 0 12788 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _571_
timestamp 1623939100
transform 1 0 15640 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_315
timestamp 1623939100
transform 1 0 15456 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_148
timestamp 1623939100
transform 1 0 14720 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_161
timestamp 1623939100
transform 1 0 15916 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1056
timestamp 1623939100
transform 1 0 16836 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_wb_clk_i
timestamp 1623939100
transform 1 0 17296 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1623939100
transform 1 0 16652 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_172
timestamp 1623939100
transform 1 0 16928 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_179
timestamp 1623939100
transform 1 0 17572 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_191
timestamp 1623939100
transform 1 0 18676 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_203
timestamp 1623939100
transform 1 0 19780 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1057
timestamp 1623939100
transform 1 0 22080 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_215
timestamp 1623939100
transform 1 0 20884 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_227
timestamp 1623939100
transform 1 0 21988 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_229
timestamp 1623939100
transform 1 0 22172 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _668_
timestamp 1623939100
transform 1 0 24012 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_254
timestamp 1623939100
transform 1 0 23828 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_241
timestamp 1623939100
transform 1 0 23276 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_252
timestamp 1623939100
transform 1 0 24288 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_264
timestamp 1623939100
transform 1 0 25392 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1058
timestamp 1623939100
transform 1 0 27324 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1623939100
transform 1 0 26128 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_275
timestamp 1623939100
transform 1 0 26404 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_283
timestamp 1623939100
transform 1 0 27140 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_286
timestamp 1623939100
transform 1 0 27416 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_298
timestamp 1623939100
transform 1 0 28520 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_310
timestamp 1623939100
transform 1 0 29624 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_322
timestamp 1623939100
transform 1 0 30728 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1059
timestamp 1623939100
transform 1 0 32568 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_334
timestamp 1623939100
transform 1 0 31832 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_343
timestamp 1623939100
transform 1 0 32660 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _756_
timestamp 1623939100
transform 1 0 35604 0 1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_49_355
timestamp 1623939100
transform 1 0 33764 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_367
timestamp 1623939100
transform 1 0 34868 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_392
timestamp 1623939100
transform 1 0 37168 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1060
timestamp 1623939100
transform 1 0 37812 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_398
timestamp 1623939100
transform 1 0 37720 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_400
timestamp 1623939100
transform 1 0 37904 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_412
timestamp 1623939100
transform 1 0 39008 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_424
timestamp 1623939100
transform 1 0 40112 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_436
timestamp 1623939100
transform 1 0 41216 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _637_
timestamp 1623939100
transform 1 0 42228 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1061
timestamp 1623939100
transform 1 0 43056 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_339
timestamp 1623939100
transform 1 0 42044 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_444
timestamp 1623939100
transform 1 0 41952 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_450
timestamp 1623939100
transform 1 0 42504 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_457
timestamp 1623939100
transform 1 0 43148 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_469
timestamp 1623939100
transform 1 0 44252 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_481
timestamp 1623939100
transform 1 0 45356 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_493
timestamp 1623939100
transform 1 0 46460 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1062
timestamp 1623939100
transform 1 0 48300 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1623939100
transform 1 0 47564 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_514
timestamp 1623939100
transform 1 0 48392 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_526
timestamp 1623939100
transform 1 0 49496 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_538
timestamp 1623939100
transform 1 0 50600 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_550
timestamp 1623939100
transform 1 0 51704 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_562
timestamp 1623939100
transform 1 0 52808 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1063
timestamp 1623939100
transform 1 0 53544 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_571
timestamp 1623939100
transform 1 0 53636 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_583
timestamp 1623939100
transform 1 0 54740 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_595
timestamp 1623939100
transform 1 0 55844 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_607
timestamp 1623939100
transform 1 0 56948 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_619
timestamp 1623939100
transform 1 0 58052 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1064
timestamp 1623939100
transform 1 0 58788 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_628
timestamp 1623939100
transform 1 0 58880 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_640
timestamp 1623939100
transform 1 0 59984 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_652
timestamp 1623939100
transform 1 0 61088 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_664
timestamp 1623939100
transform 1 0 62192 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1065
timestamp 1623939100
transform 1 0 64032 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_676
timestamp 1623939100
transform 1 0 63296 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_685
timestamp 1623939100
transform 1 0 64124 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_697
timestamp 1623939100
transform 1 0 65228 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _302_
timestamp 1623939100
transform -1 0 68908 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_132
timestamp 1623939100
transform -1 0 68080 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_709
timestamp 1623939100
transform 1 0 66332 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_721
timestamp 1623939100
transform 1 0 67436 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_725
timestamp 1623939100
transform 1 0 67804 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1066
timestamp 1623939100
transform 1 0 69276 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_737
timestamp 1623939100
transform 1 0 68908 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_742
timestamp 1623939100
transform 1 0 69368 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1623939100
transform 1 0 71024 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_754
timestamp 1623939100
transform 1 0 70472 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_763
timestamp 1623939100
transform 1 0 71300 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_775
timestamp 1623939100
transform 1 0 72404 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_787
timestamp 1623939100
transform 1 0 73508 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1067
timestamp 1623939100
transform 1 0 74520 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_795
timestamp 1623939100
transform 1 0 74244 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_799
timestamp 1623939100
transform 1 0 74612 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_811
timestamp 1623939100
transform 1 0 75716 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _630_
timestamp 1623939100
transform -1 0 76360 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_334
timestamp 1623939100
transform -1 0 76084 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_818
timestamp 1623939100
transform 1 0 76360 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_830
timestamp 1623939100
transform 1 0 77464 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_842
timestamp 1623939100
transform 1 0 78568 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_854
timestamp 1623939100
transform 1 0 79672 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1068
timestamp 1623939100
transform 1 0 79764 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_856
timestamp 1623939100
transform 1 0 79856 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_868
timestamp 1623939100
transform 1 0 80960 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_880
timestamp 1623939100
transform 1 0 82064 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_892
timestamp 1623939100
transform 1 0 83168 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1069
timestamp 1623939100
transform 1 0 85008 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_904
timestamp 1623939100
transform 1 0 84272 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_913
timestamp 1623939100
transform 1 0 85100 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _786_
timestamp 1623939100
transform -1 0 88596 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_123
timestamp 1623939100
transform -1 0 86848 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_925
timestamp 1623939100
transform 1 0 86204 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_929
timestamp 1623939100
transform 1 0 86572 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_951
timestamp 1623939100
transform 1 0 88596 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1070
timestamp 1623939100
transform 1 0 90252 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_963
timestamp 1623939100
transform 1 0 89700 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_970
timestamp 1623939100
transform 1 0 90344 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_982
timestamp 1623939100
transform 1 0 91448 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_994
timestamp 1623939100
transform 1 0 92552 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1006
timestamp 1623939100
transform 1 0 93656 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_1018
timestamp 1623939100
transform 1 0 94760 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1071
timestamp 1623939100
transform 1 0 95496 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_144
timestamp 1623939100
transform -1 0 97060 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1027
timestamp 1623939100
transform 1 0 95588 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_1039
timestamp 1623939100
transform 1 0 96692 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _375_
timestamp 1623939100
transform -1 0 98164 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1623939100
transform -1 0 98808 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_1055
timestamp 1623939100
transform 1 0 98164 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _693_
timestamp 1623939100
transform 1 0 2300 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1623939100
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_287
timestamp 1623939100
transform 1 0 2116 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1623939100
transform 1 0 1380 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_16
timestamp 1623939100
transform 1 0 2576 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1072
timestamp 1623939100
transform 1 0 3772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_28
timestamp 1623939100
transform 1 0 3680 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_30
timestamp 1623939100
transform 1 0 3864 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_42
timestamp 1623939100
transform 1 0 4968 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_54
timestamp 1623939100
transform 1 0 6072 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_66
timestamp 1623939100
transform 1 0 7176 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_78
timestamp 1623939100
transform 1 0 8280 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1073
timestamp 1623939100
transform 1 0 9016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_87
timestamp 1623939100
transform 1 0 9108 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_99
timestamp 1623939100
transform 1 0 10212 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_111
timestamp 1623939100
transform 1 0 11316 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_123
timestamp 1623939100
transform 1 0 12420 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1074
timestamp 1623939100
transform 1 0 14260 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_135
timestamp 1623939100
transform 1 0 13524 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_144
timestamp 1623939100
transform 1 0 14352 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_156
timestamp 1623939100
transform 1 0 15456 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_168
timestamp 1623939100
transform 1 0 16560 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_180
timestamp 1623939100
transform 1 0 17664 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1075
timestamp 1623939100
transform 1 0 19504 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_192
timestamp 1623939100
transform 1 0 18768 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_201
timestamp 1623939100
transform 1 0 19596 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _606_
timestamp 1623939100
transform 1 0 20884 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_310
timestamp 1623939100
transform 1 0 20700 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_218
timestamp 1623939100
transform 1 0 21160 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_230
timestamp 1623939100
transform 1 0 22264 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_242
timestamp 1623939100
transform 1 0 23368 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1076
timestamp 1623939100
transform 1 0 24748 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_254
timestamp 1623939100
transform 1 0 24472 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_258
timestamp 1623939100
transform 1 0 24840 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_270
timestamp 1623939100
transform 1 0 25944 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_282
timestamp 1623939100
transform 1 0 27048 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_294
timestamp 1623939100
transform 1 0 28152 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_306
timestamp 1623939100
transform 1 0 29256 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1077
timestamp 1623939100
transform 1 0 29992 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_315
timestamp 1623939100
transform 1 0 30084 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_327
timestamp 1623939100
transform 1 0 31188 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_339
timestamp 1623939100
transform 1 0 32292 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_351
timestamp 1623939100
transform 1 0 33396 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1078
timestamp 1623939100
transform 1 0 35236 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_363
timestamp 1623939100
transform 1 0 34500 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_372
timestamp 1623939100
transform 1 0 35328 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _657_
timestamp 1623939100
transform 1 0 36984 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_wb_clk_i
timestamp 1623939100
transform 1 0 36156 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_359
timestamp 1623939100
transform 1 0 36800 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_380
timestamp 1623939100
transform 1 0 36064 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_384
timestamp 1623939100
transform 1 0 36432 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_393
timestamp 1623939100
transform 1 0 37260 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _476_
timestamp 1623939100
transform 1 0 37996 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _636_
timestamp 1623939100
transform 1 0 39192 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_336
timestamp 1623939100
transform 1 0 39008 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_410
timestamp 1623939100
transform 1 0 38824 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1079
timestamp 1623939100
transform 1 0 40480 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_417
timestamp 1623939100
transform 1 0 39468 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_425
timestamp 1623939100
transform 1 0 40204 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_429
timestamp 1623939100
transform 1 0 40572 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_441
timestamp 1623939100
transform 1 0 41676 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_453
timestamp 1623939100
transform 1 0 42780 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_465
timestamp 1623939100
transform 1 0 43884 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_477
timestamp 1623939100
transform 1 0 44988 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _413_
timestamp 1623939100
transform 1 0 46184 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1080
timestamp 1623939100
transform 1 0 45724 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_486
timestamp 1623939100
transform 1 0 45816 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_497
timestamp 1623939100
transform 1 0 46828 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_509
timestamp 1623939100
transform 1 0 47932 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_521
timestamp 1623939100
transform 1 0 49036 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_533
timestamp 1623939100
transform 1 0 50140 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_541
timestamp 1623939100
transform 1 0 50876 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1081
timestamp 1623939100
transform 1 0 50968 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_543
timestamp 1623939100
transform 1 0 51060 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_555
timestamp 1623939100
transform 1 0 52164 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_567
timestamp 1623939100
transform 1 0 53268 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_579
timestamp 1623939100
transform 1 0 54372 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1082
timestamp 1623939100
transform 1 0 56212 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_591
timestamp 1623939100
transform 1 0 55476 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_600
timestamp 1623939100
transform 1 0 56304 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_612
timestamp 1623939100
transform 1 0 57408 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_624
timestamp 1623939100
transform 1 0 58512 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_636
timestamp 1623939100
transform 1 0 59616 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1083
timestamp 1623939100
transform 1 0 61456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_648
timestamp 1623939100
transform 1 0 60720 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_657
timestamp 1623939100
transform 1 0 61548 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_669
timestamp 1623939100
transform 1 0 62652 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_681
timestamp 1623939100
transform 1 0 63756 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_693
timestamp 1623939100
transform 1 0 64860 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_705
timestamp 1623939100
transform 1 0 65964 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _761_
timestamp 1623939100
transform 1 0 67160 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1084
timestamp 1623939100
transform 1 0 66700 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_106
timestamp 1623939100
transform 1 0 66976 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_714
timestamp 1623939100
transform 1 0 66792 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_737
timestamp 1623939100
transform 1 0 68908 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_749
timestamp 1623939100
transform 1 0 70012 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1085
timestamp 1623939100
transform 1 0 71944 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_761
timestamp 1623939100
transform 1 0 71116 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_769
timestamp 1623939100
transform 1 0 71852 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_771
timestamp 1623939100
transform 1 0 72036 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_783
timestamp 1623939100
transform 1 0 73140 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_795
timestamp 1623939100
transform 1 0 74244 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_807
timestamp 1623939100
transform 1 0 75348 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1086
timestamp 1623939100
transform 1 0 77188 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_819
timestamp 1623939100
transform 1 0 76452 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_828
timestamp 1623939100
transform 1 0 77280 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_840
timestamp 1623939100
transform 1 0 78384 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_852
timestamp 1623939100
transform 1 0 79488 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_864
timestamp 1623939100
transform 1 0 80592 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1087
timestamp 1623939100
transform 1 0 82432 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_876
timestamp 1623939100
transform 1 0 81696 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_885
timestamp 1623939100
transform 1 0 82524 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_897
timestamp 1623939100
transform 1 0 83628 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_909
timestamp 1623939100
transform 1 0 84732 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_921
timestamp 1623939100
transform 1 0 85836 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_933
timestamp 1623939100
transform 1 0 86940 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _749_
timestamp 1623939100
transform -1 0 90068 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1088
timestamp 1623939100
transform 1 0 87676 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_91
timestamp 1623939100
transform -1 0 88320 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_942
timestamp 1623939100
transform 1 0 87768 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_967
timestamp 1623939100
transform 1 0 90068 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_979
timestamp 1623939100
transform 1 0 91172 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1089
timestamp 1623939100
transform 1 0 92920 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_991
timestamp 1623939100
transform 1 0 92276 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_997
timestamp 1623939100
transform 1 0 92828 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_999
timestamp 1623939100
transform 1 0 93012 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1011
timestamp 1623939100
transform 1 0 94116 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1023
timestamp 1623939100
transform 1 0 95220 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1035
timestamp 1623939100
transform 1 0 96324 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1623939100
transform -1 0 98808 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1090
timestamp 1623939100
transform 1 0 98164 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_1047
timestamp 1623939100
transform 1 0 97428 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_1056
timestamp 1623939100
transform 1 0 98256 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1623939100
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1623939100
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1623939100
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1623939100
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1623939100
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1091
timestamp 1623939100
transform 1 0 6348 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_51
timestamp 1623939100
transform 1 0 5796 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_58
timestamp 1623939100
transform 1 0 6440 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_70
timestamp 1623939100
transform 1 0 7544 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_82
timestamp 1623939100
transform 1 0 8648 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _445_
timestamp 1623939100
transform 1 0 9752 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _775_
timestamp 1623939100
transform 1 0 12052 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1092
timestamp 1623939100
transform 1 0 11592 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_106
timestamp 1623939100
transform 1 0 10856 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_115
timestamp 1623939100
transform 1 0 11684 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_138
timestamp 1623939100
transform 1 0 13800 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_150
timestamp 1623939100
transform 1 0 14904 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_162
timestamp 1623939100
transform 1 0 16008 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1093
timestamp 1623939100
transform 1 0 16836 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_170
timestamp 1623939100
transform 1 0 16744 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_172
timestamp 1623939100
transform 1 0 16928 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1623939100
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1623939100
transform 1 0 19136 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1623939100
transform 1 0 20240 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1094
timestamp 1623939100
transform 1 0 22080 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_220
timestamp 1623939100
transform 1 0 21344 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_229
timestamp 1623939100
transform 1 0 22172 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _333_
timestamp 1623939100
transform 1 0 24012 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_51_241
timestamp 1623939100
transform 1 0 23276 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_258
timestamp 1623939100
transform 1 0 24840 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_270
timestamp 1623939100
transform 1 0 25944 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1095
timestamp 1623939100
transform 1 0 27324 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_282
timestamp 1623939100
transform 1 0 27048 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_286
timestamp 1623939100
transform 1 0 27416 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_298
timestamp 1623939100
transform 1 0 28520 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_310
timestamp 1623939100
transform 1 0 29624 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_322
timestamp 1623939100
transform 1 0 30728 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1096
timestamp 1623939100
transform 1 0 32568 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_334
timestamp 1623939100
transform 1 0 31832 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_343
timestamp 1623939100
transform 1 0 32660 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_355
timestamp 1623939100
transform 1 0 33764 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1623939100
transform 1 0 34868 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1623939100
transform 1 0 35972 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_391
timestamp 1623939100
transform 1 0 37076 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1097
timestamp 1623939100
transform 1 0 37812 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_400
timestamp 1623939100
transform 1 0 37904 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_412
timestamp 1623939100
transform 1 0 39008 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_424
timestamp 1623939100
transform 1 0 40112 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_436
timestamp 1623939100
transform 1 0 41216 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1098
timestamp 1623939100
transform 1 0 43056 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_448
timestamp 1623939100
transform 1 0 42320 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_457
timestamp 1623939100
transform 1 0 43148 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _397_
timestamp 1623939100
transform 1 0 43516 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_51_470
timestamp 1623939100
transform 1 0 44344 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_482
timestamp 1623939100
transform 1 0 45448 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_494
timestamp 1623939100
transform 1 0 46552 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1099
timestamp 1623939100
transform 1 0 48300 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_506
timestamp 1623939100
transform 1 0 47656 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_512
timestamp 1623939100
transform 1 0 48208 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_514
timestamp 1623939100
transform 1 0 48392 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_526
timestamp 1623939100
transform 1 0 49496 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_538
timestamp 1623939100
transform 1 0 50600 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_550
timestamp 1623939100
transform 1 0 51704 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_562
timestamp 1623939100
transform 1 0 52808 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1100
timestamp 1623939100
transform 1 0 53544 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_571
timestamp 1623939100
transform 1 0 53636 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_583
timestamp 1623939100
transform 1 0 54740 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_595
timestamp 1623939100
transform 1 0 55844 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_607
timestamp 1623939100
transform 1 0 56948 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_619
timestamp 1623939100
transform 1 0 58052 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1101
timestamp 1623939100
transform 1 0 58788 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_628
timestamp 1623939100
transform 1 0 58880 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_640
timestamp 1623939100
transform 1 0 59984 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_652
timestamp 1623939100
transform 1 0 61088 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_664
timestamp 1623939100
transform 1 0 62192 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _623_
timestamp 1623939100
transform -1 0 62928 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1102
timestamp 1623939100
transform 1 0 64032 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_326
timestamp 1623939100
transform -1 0 62652 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_672
timestamp 1623939100
transform 1 0 62928 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_685
timestamp 1623939100
transform 1 0 64124 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_697
timestamp 1623939100
transform 1 0 65228 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_709
timestamp 1623939100
transform 1 0 66332 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_721
timestamp 1623939100
transform 1 0 67436 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1103
timestamp 1623939100
transform 1 0 69276 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_733
timestamp 1623939100
transform 1 0 68540 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_742
timestamp 1623939100
transform 1 0 69368 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _664_
timestamp 1623939100
transform 1 0 71024 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_370
timestamp 1623939100
transform 1 0 70840 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_754
timestamp 1623939100
transform 1 0 70472 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_763
timestamp 1623939100
transform 1 0 71300 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_775
timestamp 1623939100
transform 1 0 72404 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_787
timestamp 1623939100
transform 1 0 73508 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1104
timestamp 1623939100
transform 1 0 74520 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_795
timestamp 1623939100
transform 1 0 74244 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_799
timestamp 1623939100
transform 1 0 74612 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_811
timestamp 1623939100
transform 1 0 75716 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_823
timestamp 1623939100
transform 1 0 76820 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_835
timestamp 1623939100
transform 1 0 77924 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_847
timestamp 1623939100
transform 1 0 79028 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _724_
timestamp 1623939100
transform 1 0 80224 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1105
timestamp 1623939100
transform 1 0 79764 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_856
timestamp 1623939100
transform 1 0 79856 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_879
timestamp 1623939100
transform 1 0 81972 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_891
timestamp 1623939100
transform 1 0 83076 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1106
timestamp 1623939100
transform 1 0 85008 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_903
timestamp 1623939100
transform 1 0 84180 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_911
timestamp 1623939100
transform 1 0 84916 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_913
timestamp 1623939100
transform 1 0 85100 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_925
timestamp 1623939100
transform 1 0 86204 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_937
timestamp 1623939100
transform 1 0 87308 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _753_
timestamp 1623939100
transform 1 0 87584 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _757_
timestamp 1623939100
transform 1 0 90988 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1107
timestamp 1623939100
transform 1 0 90252 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_959
timestamp 1623939100
transform 1 0 89332 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_967
timestamp 1623939100
transform 1 0 90068 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_970
timestamp 1623939100
transform 1 0 90344 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_976
timestamp 1623939100
transform 1 0 90896 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_996
timestamp 1623939100
transform 1 0 92736 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1008
timestamp 1623939100
transform 1 0 93840 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1020
timestamp 1623939100
transform 1 0 94944 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1108
timestamp 1623939100
transform 1 0 95496 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1027
timestamp 1623939100
transform 1 0 95588 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1039
timestamp 1623939100
transform 1 0 96692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1623939100
transform -1 0 98808 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_1051
timestamp 1623939100
transform 1 0 97796 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1623939100
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1623939100
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1623939100
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1623939100
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1623939100
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1623939100
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1109
timestamp 1623939100
transform 1 0 3772 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_27
timestamp 1623939100
transform 1 0 3588 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_30
timestamp 1623939100
transform 1 0 3864 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1623939100
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1623939100
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1128
timestamp 1623939100
transform 1 0 6348 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_42
timestamp 1623939100
transform 1 0 4968 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_54
timestamp 1623939100
transform 1 0 6072 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_51
timestamp 1623939100
transform 1 0 5796 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_58
timestamp 1623939100
transform 1 0 6440 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_66
timestamp 1623939100
transform 1 0 7176 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_78
timestamp 1623939100
transform 1 0 8280 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_70
timestamp 1623939100
transform 1 0 7544 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_82
timestamp 1623939100
transform 1 0 8648 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1110
timestamp 1623939100
transform 1 0 9016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_87
timestamp 1623939100
transform 1 0 9108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_99
timestamp 1623939100
transform 1 0 10212 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_94
timestamp 1623939100
transform 1 0 9752 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1129
timestamp 1623939100
transform 1 0 11592 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_111
timestamp 1623939100
transform 1 0 11316 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_123
timestamp 1623939100
transform 1 0 12420 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_106
timestamp 1623939100
transform 1 0 10856 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_115
timestamp 1623939100
transform 1 0 11684 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1111
timestamp 1623939100
transform 1 0 14260 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_135
timestamp 1623939100
transform 1 0 13524 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_144
timestamp 1623939100
transform 1 0 14352 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_127
timestamp 1623939100
transform 1 0 12788 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_139
timestamp 1623939100
transform 1 0 13892 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_156
timestamp 1623939100
transform 1 0 15456 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_151
timestamp 1623939100
transform 1 0 14996 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_163
timestamp 1623939100
transform 1 0 16100 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _784_
timestamp 1623939100
transform -1 0 19412 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1130
timestamp 1623939100
transform 1 0 16836 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_121
timestamp 1623939100
transform -1 0 17664 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_168
timestamp 1623939100
transform 1 0 16560 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_180
timestamp 1623939100
transform 1 0 17664 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_172
timestamp 1623939100
transform 1 0 16928 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1112
timestamp 1623939100
transform 1 0 19504 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_122
timestamp 1623939100
transform -1 0 19596 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_192
timestamp 1623939100
transform 1 0 18768 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_201
timestamp 1623939100
transform 1 0 19596 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_201
timestamp 1623939100
transform 1 0 19596 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1131
timestamp 1623939100
transform 1 0 22080 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_213
timestamp 1623939100
transform 1 0 20700 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_225
timestamp 1623939100
transform 1 0 21804 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_213
timestamp 1623939100
transform 1 0 20700 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_225
timestamp 1623939100
transform 1 0 21804 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_229
timestamp 1623939100
transform 1 0 22172 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _609_
timestamp 1623939100
transform 1 0 23828 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_317
timestamp 1623939100
transform 1 0 23644 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_237
timestamp 1623939100
transform 1 0 22908 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_250
timestamp 1623939100
transform 1 0 24104 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_241
timestamp 1623939100
transform 1 0 23276 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1113
timestamp 1623939100
transform 1 0 24748 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_256
timestamp 1623939100
transform 1 0 24656 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_258
timestamp 1623939100
transform 1 0 24840 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_270
timestamp 1623939100
transform 1 0 25944 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_253
timestamp 1623939100
transform 1 0 24380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_265
timestamp 1623939100
transform 1 0 25484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _567_
timestamp 1623939100
transform 1 0 27784 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1132
timestamp 1623939100
transform 1 0 27324 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_250
timestamp 1623939100
transform 1 0 27600 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_282
timestamp 1623939100
transform 1 0 27048 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_277
timestamp 1623939100
transform 1 0 26588 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_286
timestamp 1623939100
transform 1 0 27416 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_294
timestamp 1623939100
transform 1 0 28152 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_306
timestamp 1623939100
transform 1 0 29256 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1623939100
transform 1 0 28060 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1623939100
transform 1 0 29164 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1114
timestamp 1623939100
transform 1 0 29992 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_315
timestamp 1623939100
transform 1 0 30084 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_327
timestamp 1623939100
transform 1 0 31188 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1623939100
transform 1 0 30268 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_329
timestamp 1623939100
transform 1 0 31372 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1133
timestamp 1623939100
transform 1 0 32568 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_339
timestamp 1623939100
transform 1 0 32292 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_351
timestamp 1623939100
transform 1 0 33396 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_341
timestamp 1623939100
transform 1 0 32476 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_343
timestamp 1623939100
transform 1 0 32660 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1115
timestamp 1623939100
transform 1 0 35236 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_363
timestamp 1623939100
transform 1 0 34500 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_372
timestamp 1623939100
transform 1 0 35328 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_355
timestamp 1623939100
transform 1 0 33764 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1623939100
transform 1 0 34868 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_384
timestamp 1623939100
transform 1 0 36432 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1623939100
transform 1 0 35972 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_391
timestamp 1623939100
transform 1 0 37076 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1134
timestamp 1623939100
transform 1 0 37812 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_396
timestamp 1623939100
transform 1 0 37536 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_408
timestamp 1623939100
transform 1 0 38640 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_400
timestamp 1623939100
transform 1 0 37904 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_412
timestamp 1623939100
transform 1 0 39008 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1116
timestamp 1623939100
transform 1 0 40480 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_420
timestamp 1623939100
transform 1 0 39744 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_429
timestamp 1623939100
transform 1 0 40572 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_424
timestamp 1623939100
transform 1 0 40112 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_436
timestamp 1623939100
transform 1 0 41216 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1135
timestamp 1623939100
transform 1 0 43056 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_441
timestamp 1623939100
transform 1 0 41676 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_453
timestamp 1623939100
transform 1 0 42780 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_448
timestamp 1623939100
transform 1 0 42320 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_457
timestamp 1623939100
transform 1 0 43148 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _680_
timestamp 1623939100
transform 1 0 43700 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _682_
timestamp 1623939100
transform 1 0 43976 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_274
timestamp 1623939100
transform 1 0 43516 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_276
timestamp 1623939100
transform 1 0 43792 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_466
timestamp 1623939100
transform 1 0 43976 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_478
timestamp 1623939100
transform 1 0 45080 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_463
timestamp 1623939100
transform 1 0 43700 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_469
timestamp 1623939100
transform 1 0 44252 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _423_
timestamp 1623939100
transform -1 0 47196 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1117
timestamp 1623939100
transform 1 0 45724 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_152
timestamp 1623939100
transform -1 0 46368 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_484
timestamp 1623939100
transform 1 0 45632 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_486
timestamp 1623939100
transform 1 0 45816 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_481
timestamp 1623939100
transform 1 0 45356 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_493
timestamp 1623939100
transform 1 0 46460 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1136
timestamp 1623939100
transform 1 0 48300 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1623939100
transform 1 0 47196 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1623939100
transform 1 0 48300 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1623939100
transform 1 0 47564 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_514
timestamp 1623939100
transform 1 0 48392 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_525
timestamp 1623939100
transform 1 0 49404 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_537
timestamp 1623939100
transform 1 0 50508 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_541
timestamp 1623939100
transform 1 0 50876 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_526
timestamp 1623939100
transform 1 0 49496 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_538
timestamp 1623939100
transform 1 0 50600 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1118
timestamp 1623939100
transform 1 0 50968 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_543
timestamp 1623939100
transform 1 0 51060 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_555
timestamp 1623939100
transform 1 0 52164 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_550
timestamp 1623939100
transform 1 0 51704 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_562
timestamp 1623939100
transform 1 0 52808 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _700_
timestamp 1623939100
transform 1 0 54740 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1137
timestamp 1623939100
transform 1 0 53544 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_567
timestamp 1623939100
transform 1 0 53268 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_579
timestamp 1623939100
transform 1 0 54372 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_571
timestamp 1623939100
transform 1 0 53636 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1119
timestamp 1623939100
transform 1 0 56212 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_591
timestamp 1623939100
transform 1 0 55476 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_600
timestamp 1623939100
transform 1 0 56304 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_602
timestamp 1623939100
transform 1 0 56488 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_612
timestamp 1623939100
transform 1 0 57408 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_624
timestamp 1623939100
transform 1 0 58512 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_614
timestamp 1623939100
transform 1 0 57592 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _448_
timestamp 1623939100
transform 1 0 60168 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1138
timestamp 1623939100
transform 1 0 58788 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_158
timestamp 1623939100
transform 1 0 59984 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_160
timestamp 1623939100
transform 1 0 59800 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_636
timestamp 1623939100
transform 1 0 59616 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_626
timestamp 1623939100
transform 1 0 58696 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_628
timestamp 1623939100
transform 1 0 58880 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_636
timestamp 1623939100
transform 1 0 59616 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1120
timestamp 1623939100
transform 1 0 61456 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_159
timestamp 1623939100
transform 1 0 60996 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_648
timestamp 1623939100
transform 1 0 60720 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_657
timestamp 1623939100
transform 1 0 61548 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_653
timestamp 1623939100
transform 1 0 61180 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_665
timestamp 1623939100
transform 1 0 62284 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1139
timestamp 1623939100
transform 1 0 64032 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_669
timestamp 1623939100
transform 1 0 62652 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_681
timestamp 1623939100
transform 1 0 63756 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_677
timestamp 1623939100
transform 1 0 63388 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_683
timestamp 1623939100
transform 1 0 63940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_685
timestamp 1623939100
transform 1 0 64124 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_693
timestamp 1623939100
transform 1 0 64860 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_705
timestamp 1623939100
transform 1 0 65964 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_697
timestamp 1623939100
transform 1 0 65228 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _568_
timestamp 1623939100
transform -1 0 67436 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1121
timestamp 1623939100
transform 1 0 66700 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_252
timestamp 1623939100
transform -1 0 67160 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_714
timestamp 1623939100
transform 1 0 66792 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_721
timestamp 1623939100
transform 1 0 67436 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_709
timestamp 1623939100
transform 1 0 66332 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_721
timestamp 1623939100
transform 1 0 67436 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1140
timestamp 1623939100
transform 1 0 69276 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_733
timestamp 1623939100
transform 1 0 68540 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_745
timestamp 1623939100
transform 1 0 69644 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_733
timestamp 1623939100
transform 1 0 68540 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_742
timestamp 1623939100
transform 1 0 69368 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1122
timestamp 1623939100
transform 1 0 71944 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_757
timestamp 1623939100
transform 1 0 70748 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_769
timestamp 1623939100
transform 1 0 71852 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_754
timestamp 1623939100
transform 1 0 70472 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_766
timestamp 1623939100
transform 1 0 71576 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _433_
timestamp 1623939100
transform 1 0 72404 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_771
timestamp 1623939100
transform 1 0 72036 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_783
timestamp 1623939100
transform 1 0 73140 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_778
timestamp 1623939100
transform 1 0 72680 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_790
timestamp 1623939100
transform 1 0 73784 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1141
timestamp 1623939100
transform 1 0 74520 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_795
timestamp 1623939100
transform 1 0 74244 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_807
timestamp 1623939100
transform 1 0 75348 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_799
timestamp 1623939100
transform 1 0 74612 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_811
timestamp 1623939100
transform 1 0 75716 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1123
timestamp 1623939100
transform 1 0 77188 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_819
timestamp 1623939100
transform 1 0 76452 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_828
timestamp 1623939100
transform 1 0 77280 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_823
timestamp 1623939100
transform 1 0 76820 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_840
timestamp 1623939100
transform 1 0 78384 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_852
timestamp 1623939100
transform 1 0 79488 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_835
timestamp 1623939100
transform 1 0 77924 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_847
timestamp 1623939100
transform 1 0 79028 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1142
timestamp 1623939100
transform 1 0 79764 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_864
timestamp 1623939100
transform 1 0 80592 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_856
timestamp 1623939100
transform 1 0 79856 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_868
timestamp 1623939100
transform 1 0 80960 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1124
timestamp 1623939100
transform 1 0 82432 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_876
timestamp 1623939100
transform 1 0 81696 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_885
timestamp 1623939100
transform 1 0 82524 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_880
timestamp 1623939100
transform 1 0 82064 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_892
timestamp 1623939100
transform 1 0 83168 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1143
timestamp 1623939100
transform 1 0 85008 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_897
timestamp 1623939100
transform 1 0 83628 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_909
timestamp 1623939100
transform 1 0 84732 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_904
timestamp 1623939100
transform 1 0 84272 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_913
timestamp 1623939100
transform 1 0 85100 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _355_
timestamp 1623939100
transform 1 0 86204 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _669_
timestamp 1623939100
transform -1 0 87492 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_182
timestamp 1623939100
transform 1 0 86020 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_256
timestamp 1623939100
transform -1 0 87216 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_921
timestamp 1623939100
transform 1 0 85836 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_933
timestamp 1623939100
transform 1 0 86940 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_925
timestamp 1623939100
transform 1 0 86204 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_933
timestamp 1623939100
transform 1 0 86940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _613_
timestamp 1623939100
transform -1 0 89056 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1125
timestamp 1623939100
transform 1 0 87676 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_319
timestamp 1623939100
transform -1 0 88780 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_942
timestamp 1623939100
transform 1 0 87768 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_950
timestamp 1623939100
transform 1 0 88504 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_956
timestamp 1623939100
transform 1 0 89056 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_939
timestamp 1623939100
transform 1 0 87492 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_951
timestamp 1623939100
transform 1 0 88596 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1144
timestamp 1623939100
transform 1 0 90252 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_968
timestamp 1623939100
transform 1 0 90160 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_963
timestamp 1623939100
transform 1 0 89700 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_970
timestamp 1623939100
transform 1 0 90344 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1126
timestamp 1623939100
transform 1 0 92920 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_980
timestamp 1623939100
transform 1 0 91264 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_992
timestamp 1623939100
transform 1 0 92368 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_999
timestamp 1623939100
transform 1 0 93012 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_982
timestamp 1623939100
transform 1 0 91448 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_994
timestamp 1623939100
transform 1 0 92552 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _398_
timestamp 1623939100
transform 1 0 94024 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_186
timestamp 1623939100
transform 1 0 93840 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_245
timestamp 1623939100
transform 1 0 94760 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1011
timestamp 1623939100
transform 1 0 94116 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_1006
timestamp 1623939100
transform 1 0 93656 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1020
timestamp 1623939100
transform 1 0 94944 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1145
timestamp 1623939100
transform 1 0 95496 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1023
timestamp 1623939100
transform 1 0 95220 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1035
timestamp 1623939100
transform 1 0 96324 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1027
timestamp 1623939100
transform 1 0 95588 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1039
timestamp 1623939100
transform 1 0 96692 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1623939100
transform -1 0 98808 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1623939100
transform -1 0 98808 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1127
timestamp 1623939100
transform 1 0 98164 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_1047
timestamp 1623939100
transform 1 0 97428 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_1056
timestamp 1623939100
transform 1 0 98256 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_1051
timestamp 1623939100
transform 1 0 97796 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1623939100
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1623939100
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1623939100
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1146
timestamp 1623939100
transform 1 0 3772 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_27
timestamp 1623939100
transform 1 0 3588 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_30
timestamp 1623939100
transform 1 0 3864 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_42
timestamp 1623939100
transform 1 0 4968 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_54
timestamp 1623939100
transform 1 0 6072 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_66
timestamp 1623939100
transform 1 0 7176 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_78
timestamp 1623939100
transform 1 0 8280 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1147
timestamp 1623939100
transform 1 0 9016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_87
timestamp 1623939100
transform 1 0 9108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_99
timestamp 1623939100
transform 1 0 10212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_111
timestamp 1623939100
transform 1 0 11316 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_123
timestamp 1623939100
transform 1 0 12420 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _367_
timestamp 1623939100
transform 1 0 13064 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1148
timestamp 1623939100
transform 1 0 14260 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_129
timestamp 1623939100
transform 1 0 12972 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_139
timestamp 1623939100
transform 1 0 13892 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_144
timestamp 1623939100
transform 1 0 14352 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_156
timestamp 1623939100
transform 1 0 15456 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _540_
timestamp 1623939100
transform 1 0 16744 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_54_168
timestamp 1623939100
transform 1 0 16560 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_179
timestamp 1623939100
transform 1 0 17572 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1149
timestamp 1623939100
transform 1 0 19504 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_191
timestamp 1623939100
transform 1 0 18676 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_199
timestamp 1623939100
transform 1 0 19412 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_201
timestamp 1623939100
transform 1 0 19596 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_213
timestamp 1623939100
transform 1 0 20700 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_225
timestamp 1623939100
transform 1 0 21804 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_237
timestamp 1623939100
transform 1 0 22908 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_249
timestamp 1623939100
transform 1 0 24012 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1150
timestamp 1623939100
transform 1 0 24748 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_258
timestamp 1623939100
transform 1 0 24840 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_270
timestamp 1623939100
transform 1 0 25944 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_282
timestamp 1623939100
transform 1 0 27048 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_294
timestamp 1623939100
transform 1 0 28152 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_306
timestamp 1623939100
transform 1 0 29256 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1151
timestamp 1623939100
transform 1 0 29992 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_315
timestamp 1623939100
transform 1 0 30084 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_327
timestamp 1623939100
transform 1 0 31188 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _316_
timestamp 1623939100
transform 1 0 33488 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_339
timestamp 1623939100
transform 1 0 32292 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_351
timestamp 1623939100
transform 1 0 33396 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1152
timestamp 1623939100
transform 1 0 35236 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_358
timestamp 1623939100
transform 1 0 34040 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_370
timestamp 1623939100
transform 1 0 35144 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_372
timestamp 1623939100
transform 1 0 35328 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_384
timestamp 1623939100
transform 1 0 36432 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_396
timestamp 1623939100
transform 1 0 37536 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_408
timestamp 1623939100
transform 1 0 38640 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1153
timestamp 1623939100
transform 1 0 40480 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_420
timestamp 1623939100
transform 1 0 39744 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_429
timestamp 1623939100
transform 1 0 40572 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_441
timestamp 1623939100
transform 1 0 41676 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_453
timestamp 1623939100
transform 1 0 42780 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _688_
timestamp 1623939100
transform 1 0 45080 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_282
timestamp 1623939100
transform 1 0 44896 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_465
timestamp 1623939100
transform 1 0 43884 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_473
timestamp 1623939100
transform 1 0 44620 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1154
timestamp 1623939100
transform 1 0 45724 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_481
timestamp 1623939100
transform 1 0 45356 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_486
timestamp 1623939100
transform 1 0 45816 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_498
timestamp 1623939100
transform 1 0 46920 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_510
timestamp 1623939100
transform 1 0 48024 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_522
timestamp 1623939100
transform 1 0 49128 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_534
timestamp 1623939100
transform 1 0 50232 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _769_
timestamp 1623939100
transform 1 0 52808 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1155
timestamp 1623939100
transform 1 0 50968 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_543
timestamp 1623939100
transform 1 0 51060 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_555
timestamp 1623939100
transform 1 0 52164 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_561
timestamp 1623939100
transform 1 0 52716 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_581
timestamp 1623939100
transform 1 0 54556 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1156
timestamp 1623939100
transform 1 0 56212 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_593
timestamp 1623939100
transform 1 0 55660 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_600
timestamp 1623939100
transform 1 0 56304 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _537_
timestamp 1623939100
transform 1 0 57960 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_54_612
timestamp 1623939100
transform 1 0 57408 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_627
timestamp 1623939100
transform 1 0 58788 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_639
timestamp 1623939100
transform 1 0 59892 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1157
timestamp 1623939100
transform 1 0 61456 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_651
timestamp 1623939100
transform 1 0 60996 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_655
timestamp 1623939100
transform 1 0 61364 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_657
timestamp 1623939100
transform 1 0 61548 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_669
timestamp 1623939100
transform 1 0 62652 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_681
timestamp 1623939100
transform 1 0 63756 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_693
timestamp 1623939100
transform 1 0 64860 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_705
timestamp 1623939100
transform 1 0 65964 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1158
timestamp 1623939100
transform 1 0 66700 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_714
timestamp 1623939100
transform 1 0 66792 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_726
timestamp 1623939100
transform 1 0 67896 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_738
timestamp 1623939100
transform 1 0 69000 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_750
timestamp 1623939100
transform 1 0 70104 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1159
timestamp 1623939100
transform 1 0 71944 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_762
timestamp 1623939100
transform 1 0 71208 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_771
timestamp 1623939100
transform 1 0 72036 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_783
timestamp 1623939100
transform 1 0 73140 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_795
timestamp 1623939100
transform 1 0 74244 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_807
timestamp 1623939100
transform 1 0 75348 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1160
timestamp 1623939100
transform 1 0 77188 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_819
timestamp 1623939100
transform 1 0 76452 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_828
timestamp 1623939100
transform 1 0 77280 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_840
timestamp 1623939100
transform 1 0 78384 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_852
timestamp 1623939100
transform 1 0 79488 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_864
timestamp 1623939100
transform 1 0 80592 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1161
timestamp 1623939100
transform 1 0 82432 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_876
timestamp 1623939100
transform 1 0 81696 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_885
timestamp 1623939100
transform 1 0 82524 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_897
timestamp 1623939100
transform 1 0 83628 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_909
timestamp 1623939100
transform 1 0 84732 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_921
timestamp 1623939100
transform 1 0 85836 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_933
timestamp 1623939100
transform 1 0 86940 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_4  _415_
timestamp 1623939100
transform 1 0 89148 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1162
timestamp 1623939100
transform 1 0 87676 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_151
timestamp 1623939100
transform 1 0 88964 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_942
timestamp 1623939100
transform 1 0 87768 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_954
timestamp 1623939100
transform 1 0 88872 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _590_
timestamp 1623939100
transform -1 0 91264 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_298
timestamp 1623939100
transform -1 0 90988 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_973
timestamp 1623939100
transform 1 0 90620 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1163
timestamp 1623939100
transform 1 0 92920 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_980
timestamp 1623939100
transform 1 0 91264 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_992
timestamp 1623939100
transform 1 0 92368 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_999
timestamp 1623939100
transform 1 0 93012 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1623939100
transform 1 0 94944 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_230
timestamp 1623939100
transform 1 0 94760 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1011
timestamp 1623939100
transform 1 0 94116 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1017
timestamp 1623939100
transform 1 0 94668 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_4  _515_
timestamp 1623939100
transform 1 0 95864 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1623939100
transform 1 0 95680 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1623939100
transform 1 0 95496 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1623939100
transform 1 0 95312 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1623939100
transform 1 0 95128 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1623939100
transform -1 0 98808 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1164
timestamp 1623939100
transform 1 0 98164 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1623939100
transform 1 0 97336 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1623939100
transform 1 0 97520 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1623939100
transform 1 0 97704 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1623939100
transform 1 0 97888 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1054
timestamp 1623939100
transform 1 0 98072 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_1056
timestamp 1623939100
transform 1 0 98256 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1623939100
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1623939100
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1623939100
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1623939100
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1623939100
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1165
timestamp 1623939100
transform 1 0 6348 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_51
timestamp 1623939100
transform 1 0 5796 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_58
timestamp 1623939100
transform 1 0 6440 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_70
timestamp 1623939100
transform 1 0 7544 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_82
timestamp 1623939100
transform 1 0 8648 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_94
timestamp 1623939100
transform 1 0 9752 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1166
timestamp 1623939100
transform 1 0 11592 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_106
timestamp 1623939100
transform 1 0 10856 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_115
timestamp 1623939100
transform 1 0 11684 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _577_
timestamp 1623939100
transform 1 0 13524 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_375
timestamp 1623939100
transform 1 0 13340 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_127
timestamp 1623939100
transform 1 0 12788 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_138
timestamp 1623939100
transform 1 0 13800 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_150
timestamp 1623939100
transform 1 0 14904 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_162
timestamp 1623939100
transform 1 0 16008 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1167
timestamp 1623939100
transform 1 0 16836 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_170
timestamp 1623939100
transform 1 0 16744 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_172
timestamp 1623939100
transform 1 0 16928 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1623939100
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1623939100
transform 1 0 19136 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1623939100
transform 1 0 20240 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1168
timestamp 1623939100
transform 1 0 22080 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_220
timestamp 1623939100
transform 1 0 21344 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_229
timestamp 1623939100
transform 1 0 22172 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_1  _328_
timestamp 1623939100
transform -1 0 23092 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_207
timestamp 1623939100
transform -1 0 22540 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_239
timestamp 1623939100
transform 1 0 23092 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_251
timestamp 1623939100
transform 1 0 24196 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_263
timestamp 1623939100
transform 1 0 25300 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _379_
timestamp 1623939100
transform 1 0 27784 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1169
timestamp 1623939100
transform 1 0 27324 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_275
timestamp 1623939100
transform 1 0 26404 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_283
timestamp 1623939100
transform 1 0 27140 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_286
timestamp 1623939100
transform 1 0 27416 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_299
timestamp 1623939100
transform 1 0 28612 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_311
timestamp 1623939100
transform 1 0 29716 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _673_
timestamp 1623939100
transform 1 0 31648 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_262
timestamp 1623939100
transform 1 0 31464 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_323
timestamp 1623939100
transform 1 0 30820 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_329
timestamp 1623939100
transform 1 0 31372 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1170
timestamp 1623939100
transform 1 0 32568 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_335
timestamp 1623939100
transform 1 0 31924 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_341
timestamp 1623939100
transform 1 0 32476 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_343
timestamp 1623939100
transform 1 0 32660 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_355
timestamp 1623939100
transform 1 0 33764 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1623939100
transform 1 0 34868 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1623939100
transform 1 0 35972 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_391
timestamp 1623939100
transform 1 0 37076 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1171
timestamp 1623939100
transform 1 0 37812 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_400
timestamp 1623939100
transform 1 0 37904 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_412
timestamp 1623939100
transform 1 0 39008 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _746_
timestamp 1623939100
transform 1 0 40112 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1172
timestamp 1623939100
transform 1 0 43056 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_443
timestamp 1623939100
transform 1 0 41860 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_455
timestamp 1623939100
transform 1 0 42964 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_457
timestamp 1623939100
transform 1 0 43148 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_469
timestamp 1623939100
transform 1 0 44252 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_481
timestamp 1623939100
transform 1 0 45356 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_493
timestamp 1623939100
transform 1 0 46460 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1173
timestamp 1623939100
transform 1 0 48300 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1623939100
transform 1 0 47564 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_514
timestamp 1623939100
transform 1 0 48392 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_526
timestamp 1623939100
transform 1 0 49496 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_538
timestamp 1623939100
transform 1 0 50600 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_550
timestamp 1623939100
transform 1 0 51704 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_562
timestamp 1623939100
transform 1 0 52808 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1174
timestamp 1623939100
transform 1 0 53544 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_571
timestamp 1623939100
transform 1 0 53636 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_583
timestamp 1623939100
transform 1 0 54740 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_4  _523_
timestamp 1623939100
transform 1 0 55752 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_55_591
timestamp 1623939100
transform 1 0 55476 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_610
timestamp 1623939100
transform 1 0 57224 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_622
timestamp 1623939100
transform 1 0 58328 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1175
timestamp 1623939100
transform 1 0 58788 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_626
timestamp 1623939100
transform 1 0 58696 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_628
timestamp 1623939100
transform 1 0 58880 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_640
timestamp 1623939100
transform 1 0 59984 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_652
timestamp 1623939100
transform 1 0 61088 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_664
timestamp 1623939100
transform 1 0 62192 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1176
timestamp 1623939100
transform 1 0 64032 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_676
timestamp 1623939100
transform 1 0 63296 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_685
timestamp 1623939100
transform 1 0 64124 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_697
timestamp 1623939100
transform 1 0 65228 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_709
timestamp 1623939100
transform 1 0 66332 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_721
timestamp 1623939100
transform 1 0 67436 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1177
timestamp 1623939100
transform 1 0 69276 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_733
timestamp 1623939100
transform 1 0 68540 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_742
timestamp 1623939100
transform 1 0 69368 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_754
timestamp 1623939100
transform 1 0 70472 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_766
timestamp 1623939100
transform 1 0 71576 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_778
timestamp 1623939100
transform 1 0 72680 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_790
timestamp 1623939100
transform 1 0 73784 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1178
timestamp 1623939100
transform 1 0 74520 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_799
timestamp 1623939100
transform 1 0 74612 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_811
timestamp 1623939100
transform 1 0 75716 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_823
timestamp 1623939100
transform 1 0 76820 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_835
timestamp 1623939100
transform 1 0 77924 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_847
timestamp 1623939100
transform 1 0 79028 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1179
timestamp 1623939100
transform 1 0 79764 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_856
timestamp 1623939100
transform 1 0 79856 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_868
timestamp 1623939100
transform 1 0 80960 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_880
timestamp 1623939100
transform 1 0 82064 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_892
timestamp 1623939100
transform 1 0 83168 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1180
timestamp 1623939100
transform 1 0 85008 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_904
timestamp 1623939100
transform 1 0 84272 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_913
timestamp 1623939100
transform 1 0 85100 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_925
timestamp 1623939100
transform 1 0 86204 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_937
timestamp 1623939100
transform 1 0 87308 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_949
timestamp 1623939100
transform 1 0 88412 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1181
timestamp 1623939100
transform 1 0 90252 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_961
timestamp 1623939100
transform 1 0 89516 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_970
timestamp 1623939100
transform 1 0 90344 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_982
timestamp 1623939100
transform 1 0 91448 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_994
timestamp 1623939100
transform 1 0 92552 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1006
timestamp 1623939100
transform 1 0 93656 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_1018
timestamp 1623939100
transform 1 0 94760 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1182
timestamp 1623939100
transform 1 0 95496 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1027
timestamp 1623939100
transform 1 0 95588 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1039
timestamp 1623939100
transform 1 0 96692 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1623939100
transform -1 0 98808 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_1051
timestamp 1623939100
transform 1 0 97796 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1623939100
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1623939100
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1623939100
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1183
timestamp 1623939100
transform 1 0 3772 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_27
timestamp 1623939100
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_30
timestamp 1623939100
transform 1 0 3864 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _587_
timestamp 1623939100
transform 1 0 6532 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_293
timestamp 1623939100
transform 1 0 6348 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_42
timestamp 1623939100
transform 1 0 4968 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_54
timestamp 1623939100
transform 1 0 6072 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_62
timestamp 1623939100
transform 1 0 6808 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_74
timestamp 1623939100
transform 1 0 7912 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1184
timestamp 1623939100
transform 1 0 9016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_87
timestamp 1623939100
transform 1 0 9108 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_99
timestamp 1623939100
transform 1 0 10212 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_111
timestamp 1623939100
transform 1 0 11316 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_123
timestamp 1623939100
transform 1 0 12420 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _588_
timestamp 1623939100
transform 1 0 13432 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1185
timestamp 1623939100
transform 1 0 14260 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_296
timestamp 1623939100
transform 1 0 13248 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_131
timestamp 1623939100
transform 1 0 13156 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_137
timestamp 1623939100
transform 1 0 13708 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_144
timestamp 1623939100
transform 1 0 14352 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_156
timestamp 1623939100
transform 1 0 15456 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_168
timestamp 1623939100
transform 1 0 16560 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_180
timestamp 1623939100
transform 1 0 17664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1186
timestamp 1623939100
transform 1 0 19504 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_192
timestamp 1623939100
transform 1 0 18768 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_201
timestamp 1623939100
transform 1 0 19596 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _492_
timestamp 1623939100
transform 1 0 21988 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_56_213
timestamp 1623939100
transform 1 0 20700 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_225
timestamp 1623939100
transform 1 0 21804 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_236
timestamp 1623939100
transform 1 0 22816 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_248
timestamp 1623939100
transform 1 0 23920 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1187
timestamp 1623939100
transform 1 0 24748 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_256
timestamp 1623939100
transform 1 0 24656 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_258
timestamp 1623939100
transform 1 0 24840 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_270
timestamp 1623939100
transform 1 0 25944 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_282
timestamp 1623939100
transform 1 0 27048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_294
timestamp 1623939100
transform 1 0 28152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_306
timestamp 1623939100
transform 1 0 29256 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1188
timestamp 1623939100
transform 1 0 29992 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_315
timestamp 1623939100
transform 1 0 30084 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_327
timestamp 1623939100
transform 1 0 31188 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_339
timestamp 1623939100
transform 1 0 32292 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_351
timestamp 1623939100
transform 1 0 33396 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1189
timestamp 1623939100
transform 1 0 35236 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_363
timestamp 1623939100
transform 1 0 34500 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_372
timestamp 1623939100
transform 1 0 35328 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_384
timestamp 1623939100
transform 1 0 36432 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _314_
timestamp 1623939100
transform 1 0 39008 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_136
timestamp 1623939100
transform 1 0 38824 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_396
timestamp 1623939100
transform 1 0 37536 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_408
timestamp 1623939100
transform 1 0 38640 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1190
timestamp 1623939100
transform 1 0 40480 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_421
timestamp 1623939100
transform 1 0 39836 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_427
timestamp 1623939100
transform 1 0 40388 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_429
timestamp 1623939100
transform 1 0 40572 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _416_
timestamp 1623939100
transform 1 0 41860 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_441
timestamp 1623939100
transform 1 0 41676 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_449
timestamp 1623939100
transform 1 0 42412 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_461
timestamp 1623939100
transform 1 0 43516 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_473
timestamp 1623939100
transform 1 0 44620 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _402_
timestamp 1623939100
transform 1 0 46828 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1191
timestamp 1623939100
transform 1 0 45724 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_486
timestamp 1623939100
transform 1 0 45816 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_494
timestamp 1623939100
transform 1 0 46552 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_506
timestamp 1623939100
transform 1 0 47656 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_518
timestamp 1623939100
transform 1 0 48760 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_530
timestamp 1623939100
transform 1 0 49864 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1192
timestamp 1623939100
transform 1 0 50968 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_543
timestamp 1623939100
transform 1 0 51060 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_555
timestamp 1623939100
transform 1 0 52164 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_567
timestamp 1623939100
transform 1 0 53268 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_579
timestamp 1623939100
transform 1 0 54372 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1193
timestamp 1623939100
transform 1 0 56212 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_591
timestamp 1623939100
transform 1 0 55476 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_600
timestamp 1623939100
transform 1 0 56304 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_612
timestamp 1623939100
transform 1 0 57408 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_624
timestamp 1623939100
transform 1 0 58512 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_636
timestamp 1623939100
transform 1 0 59616 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1194
timestamp 1623939100
transform 1 0 61456 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_648
timestamp 1623939100
transform 1 0 60720 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_657
timestamp 1623939100
transform 1 0 61548 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_669
timestamp 1623939100
transform 1 0 62652 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_681
timestamp 1623939100
transform 1 0 63756 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_693
timestamp 1623939100
transform 1 0 64860 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_705
timestamp 1623939100
transform 1 0 65964 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1195
timestamp 1623939100
transform 1 0 66700 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_714
timestamp 1623939100
transform 1 0 66792 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_726
timestamp 1623939100
transform 1 0 67896 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_738
timestamp 1623939100
transform 1 0 69000 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_750
timestamp 1623939100
transform 1 0 70104 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1196
timestamp 1623939100
transform 1 0 71944 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_762
timestamp 1623939100
transform 1 0 71208 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_771
timestamp 1623939100
transform 1 0 72036 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_783
timestamp 1623939100
transform 1 0 73140 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_795
timestamp 1623939100
transform 1 0 74244 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_807
timestamp 1623939100
transform 1 0 75348 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1197
timestamp 1623939100
transform 1 0 77188 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_819
timestamp 1623939100
transform 1 0 76452 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_828
timestamp 1623939100
transform 1 0 77280 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_840
timestamp 1623939100
transform 1 0 78384 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_852
timestamp 1623939100
transform 1 0 79488 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_864
timestamp 1623939100
transform 1 0 80592 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1198
timestamp 1623939100
transform 1 0 82432 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_876
timestamp 1623939100
transform 1 0 81696 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_885
timestamp 1623939100
transform 1 0 82524 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_897
timestamp 1623939100
transform 1 0 83628 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_909
timestamp 1623939100
transform 1 0 84732 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_921
timestamp 1623939100
transform 1 0 85836 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_933
timestamp 1623939100
transform 1 0 86940 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1199
timestamp 1623939100
transform 1 0 87676 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_942
timestamp 1623939100
transform 1 0 87768 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_954
timestamp 1623939100
transform 1 0 88872 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _332_
timestamp 1623939100
transform 1 0 90252 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_56_966
timestamp 1623939100
transform 1 0 89976 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_975
timestamp 1623939100
transform 1 0 90804 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1200
timestamp 1623939100
transform 1 0 92920 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_987
timestamp 1623939100
transform 1 0 91908 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_995
timestamp 1623939100
transform 1 0 92644 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_999
timestamp 1623939100
transform 1 0 93012 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1011
timestamp 1623939100
transform 1 0 94116 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1023
timestamp 1623939100
transform 1 0 95220 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1035
timestamp 1623939100
transform 1 0 96324 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1623939100
transform -1 0 98808 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1201
timestamp 1623939100
transform 1 0 98164 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_1047
timestamp 1623939100
transform 1 0 97428 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_1056
timestamp 1623939100
transform 1 0 98256 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1623939100
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1623939100
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1623939100
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1623939100
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1623939100
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1202
timestamp 1623939100
transform 1 0 6348 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_51
timestamp 1623939100
transform 1 0 5796 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_58
timestamp 1623939100
transform 1 0 6440 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_70
timestamp 1623939100
transform 1 0 7544 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_82
timestamp 1623939100
transform 1 0 8648 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_94
timestamp 1623939100
transform 1 0 9752 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1203
timestamp 1623939100
transform 1 0 11592 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_106
timestamp 1623939100
transform 1 0 10856 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_115
timestamp 1623939100
transform 1 0 11684 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_127
timestamp 1623939100
transform 1 0 12788 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_139
timestamp 1623939100
transform 1 0 13892 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_151
timestamp 1623939100
transform 1 0 14996 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_163
timestamp 1623939100
transform 1 0 16100 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _765_
timestamp 1623939100
transform 1 0 17296 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1204
timestamp 1623939100
transform 1 0 16836 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_172
timestamp 1623939100
transform 1 0 16928 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_4  _486_
timestamp 1623939100
transform 1 0 20240 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1623939100
transform 1 0 20056 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1623939100
transform 1 0 19872 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1623939100
transform 1 0 19688 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_233
timestamp 1623939100
transform 1 0 19504 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_195
timestamp 1623939100
transform 1 0 19044 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_199
timestamp 1623939100
transform 1 0 19412 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1205
timestamp 1623939100
transform 1 0 22080 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1623939100
transform 1 0 21712 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1623939100
transform 1 0 21896 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1623939100
transform 1 0 22172 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_231
timestamp 1623939100
transform 1 0 22356 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_243
timestamp 1623939100
transform 1 0 23460 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _455_
timestamp 1623939100
transform 1 0 24380 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_57_251
timestamp 1623939100
transform 1 0 24196 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_262
timestamp 1623939100
transform 1 0 25208 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1206
timestamp 1623939100
transform 1 0 27324 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_274
timestamp 1623939100
transform 1 0 26312 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_282
timestamp 1623939100
transform 1 0 27048 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_286
timestamp 1623939100
transform 1 0 27416 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_298
timestamp 1623939100
transform 1 0 28520 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_310
timestamp 1623939100
transform 1 0 29624 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _382_
timestamp 1623939100
transform 1 0 30176 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_57_323
timestamp 1623939100
transform 1 0 30820 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1207
timestamp 1623939100
transform 1 0 32568 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_335
timestamp 1623939100
transform 1 0 31924 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_341
timestamp 1623939100
transform 1 0 32476 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_343
timestamp 1623939100
transform 1 0 32660 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_355
timestamp 1623939100
transform 1 0 33764 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1623939100
transform 1 0 34868 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_379
timestamp 1623939100
transform 1 0 35972 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_391
timestamp 1623939100
transform 1 0 37076 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1208
timestamp 1623939100
transform 1 0 37812 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_400
timestamp 1623939100
transform 1 0 37904 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_412
timestamp 1623939100
transform 1 0 39008 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _777_
timestamp 1623939100
transform 1 0 40112 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_117
timestamp 1623939100
transform 1 0 39928 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_420
timestamp 1623939100
transform 1 0 39744 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1209
timestamp 1623939100
transform 1 0 43056 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_443
timestamp 1623939100
transform 1 0 41860 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_455
timestamp 1623939100
transform 1 0 42964 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_457
timestamp 1623939100
transform 1 0 43148 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_469
timestamp 1623939100
transform 1 0 44252 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_481
timestamp 1623939100
transform 1 0 45356 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_493
timestamp 1623939100
transform 1 0 46460 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1210
timestamp 1623939100
transform 1 0 48300 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1623939100
transform 1 0 47564 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_514
timestamp 1623939100
transform 1 0 48392 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _344_
timestamp 1623939100
transform 1 0 49220 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_522
timestamp 1623939100
transform 1 0 49128 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1623939100
transform 1 0 49772 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1623939100
transform 1 0 50876 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_553
timestamp 1623939100
transform 1 0 51980 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1211
timestamp 1623939100
transform 1 0 53544 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_565
timestamp 1623939100
transform 1 0 53084 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_569
timestamp 1623939100
transform 1 0 53452 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_571
timestamp 1623939100
transform 1 0 53636 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_583
timestamp 1623939100
transform 1 0 54740 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_595
timestamp 1623939100
transform 1 0 55844 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_607
timestamp 1623939100
transform 1 0 56948 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_619
timestamp 1623939100
transform 1 0 58052 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _315_
timestamp 1623939100
transform 1 0 59248 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _443_
timestamp 1623939100
transform 1 0 60444 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1212
timestamp 1623939100
transform 1 0 58788 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_628
timestamp 1623939100
transform 1 0 58880 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_641
timestamp 1623939100
transform 1 0 60076 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_654
timestamp 1623939100
transform 1 0 61272 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_666
timestamp 1623939100
transform 1 0 62376 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1213
timestamp 1623939100
transform 1 0 64032 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_678
timestamp 1623939100
transform 1 0 63480 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_685
timestamp 1623939100
transform 1 0 64124 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_697
timestamp 1623939100
transform 1 0 65228 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_709
timestamp 1623939100
transform 1 0 66332 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_721
timestamp 1623939100
transform 1 0 67436 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1214
timestamp 1623939100
transform 1 0 69276 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_733
timestamp 1623939100
transform 1 0 68540 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_742
timestamp 1623939100
transform 1 0 69368 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_754
timestamp 1623939100
transform 1 0 70472 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_766
timestamp 1623939100
transform 1 0 71576 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_778
timestamp 1623939100
transform 1 0 72680 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_790
timestamp 1623939100
transform 1 0 73784 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1215
timestamp 1623939100
transform 1 0 74520 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_799
timestamp 1623939100
transform 1 0 74612 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_811
timestamp 1623939100
transform 1 0 75716 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_823
timestamp 1623939100
transform 1 0 76820 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_835
timestamp 1623939100
transform 1 0 77924 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_847
timestamp 1623939100
transform 1 0 79028 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1216
timestamp 1623939100
transform 1 0 79764 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_856
timestamp 1623939100
transform 1 0 79856 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_868
timestamp 1623939100
transform 1 0 80960 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_880
timestamp 1623939100
transform 1 0 82064 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_892
timestamp 1623939100
transform 1 0 83168 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1217
timestamp 1623939100
transform 1 0 85008 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_904
timestamp 1623939100
transform 1 0 84272 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_913
timestamp 1623939100
transform 1 0 85100 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_925
timestamp 1623939100
transform 1 0 86204 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_937
timestamp 1623939100
transform 1 0 87308 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_949
timestamp 1623939100
transform 1 0 88412 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1218
timestamp 1623939100
transform 1 0 90252 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_961
timestamp 1623939100
transform 1 0 89516 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_970
timestamp 1623939100
transform 1 0 90344 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_982
timestamp 1623939100
transform 1 0 91448 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_994
timestamp 1623939100
transform 1 0 92552 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1006
timestamp 1623939100
transform 1 0 93656 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_1018
timestamp 1623939100
transform 1 0 94760 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1219
timestamp 1623939100
transform 1 0 95496 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1027
timestamp 1623939100
transform 1 0 95588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1039
timestamp 1623939100
transform 1 0 96692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1623939100
transform -1 0 98808 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_1051
timestamp 1623939100
transform 1 0 97796 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1623939100
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1623939100
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1623939100
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1220
timestamp 1623939100
transform 1 0 3772 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_27
timestamp 1623939100
transform 1 0 3588 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_30
timestamp 1623939100
transform 1 0 3864 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_42
timestamp 1623939100
transform 1 0 4968 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_54
timestamp 1623939100
transform 1 0 6072 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_66
timestamp 1623939100
transform 1 0 7176 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_78
timestamp 1623939100
transform 1 0 8280 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _368_
timestamp 1623939100
transform 1 0 9476 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1221
timestamp 1623939100
transform 1 0 9016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_87
timestamp 1623939100
transform 1 0 9108 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_103
timestamp 1623939100
transform 1 0 10580 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_115
timestamp 1623939100
transform 1 0 11684 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1222
timestamp 1623939100
transform 1 0 14260 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_127
timestamp 1623939100
transform 1 0 12788 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_139
timestamp 1623939100
transform 1 0 13892 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_144
timestamp 1623939100
transform 1 0 14352 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_156
timestamp 1623939100
transform 1 0 15456 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _547_
timestamp 1623939100
transform -1 0 18768 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_133
timestamp 1623939100
transform -1 0 17940 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_168
timestamp 1623939100
transform 1 0 16560 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_180
timestamp 1623939100
transform 1 0 17664 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1223
timestamp 1623939100
transform 1 0 19504 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_192
timestamp 1623939100
transform 1 0 18768 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_201
timestamp 1623939100
transform 1 0 19596 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _792_
timestamp 1623939100
transform 1 0 21528 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_58_213
timestamp 1623939100
transform 1 0 20700 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_221
timestamp 1623939100
transform 1 0 21436 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_241
timestamp 1623939100
transform 1 0 23276 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1224
timestamp 1623939100
transform 1 0 24748 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1623939100
transform 1 0 24380 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_258
timestamp 1623939100
transform 1 0 24840 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_270
timestamp 1623939100
transform 1 0 25944 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _648_
timestamp 1623939100
transform 1 0 27692 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_351
timestamp 1623939100
transform 1 0 27508 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_282
timestamp 1623939100
transform 1 0 27048 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_286
timestamp 1623939100
transform 1 0 27416 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_292
timestamp 1623939100
transform 1 0 27968 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_304
timestamp 1623939100
transform 1 0 29072 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_312
timestamp 1623939100
transform 1 0 29808 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1225
timestamp 1623939100
transform 1 0 29992 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_315
timestamp 1623939100
transform 1 0 30084 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_327
timestamp 1623939100
transform 1 0 31188 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_339
timestamp 1623939100
transform 1 0 32292 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_351
timestamp 1623939100
transform 1 0 33396 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1226
timestamp 1623939100
transform 1 0 35236 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_363
timestamp 1623939100
transform 1 0 34500 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_372
timestamp 1623939100
transform 1 0 35328 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_384
timestamp 1623939100
transform 1 0 36432 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_396
timestamp 1623939100
transform 1 0 37536 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_408
timestamp 1623939100
transform 1 0 38640 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1227
timestamp 1623939100
transform 1 0 40480 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_420
timestamp 1623939100
transform 1 0 39744 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_429
timestamp 1623939100
transform 1 0 40572 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_2  _406_
timestamp 1623939100
transform 1 0 41952 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_58_441
timestamp 1623939100
transform 1 0 41676 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_451
timestamp 1623939100
transform 1 0 42596 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_463
timestamp 1623939100
transform 1 0 43700 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_475
timestamp 1623939100
transform 1 0 44804 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1228
timestamp 1623939100
transform 1 0 45724 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_483
timestamp 1623939100
transform 1 0 45540 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_486
timestamp 1623939100
transform 1 0 45816 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_498
timestamp 1623939100
transform 1 0 46920 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_510
timestamp 1623939100
transform 1 0 48024 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_522
timestamp 1623939100
transform 1 0 49128 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_534
timestamp 1623939100
transform 1 0 50232 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1229
timestamp 1623939100
transform 1 0 50968 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_543
timestamp 1623939100
transform 1 0 51060 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_555
timestamp 1623939100
transform 1 0 52164 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_567
timestamp 1623939100
transform 1 0 53268 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_579
timestamp 1623939100
transform 1 0 54372 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1230
timestamp 1623939100
transform 1 0 56212 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_591
timestamp 1623939100
transform 1 0 55476 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_600
timestamp 1623939100
transform 1 0 56304 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_612
timestamp 1623939100
transform 1 0 57408 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_624
timestamp 1623939100
transform 1 0 58512 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_636
timestamp 1623939100
transform 1 0 59616 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1231
timestamp 1623939100
transform 1 0 61456 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_648
timestamp 1623939100
transform 1 0 60720 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_657
timestamp 1623939100
transform 1 0 61548 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_669
timestamp 1623939100
transform 1 0 62652 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_681
timestamp 1623939100
transform 1 0 63756 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_693
timestamp 1623939100
transform 1 0 64860 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_705
timestamp 1623939100
transform 1 0 65964 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1232
timestamp 1623939100
transform 1 0 66700 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_714
timestamp 1623939100
transform 1 0 66792 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_726
timestamp 1623939100
transform 1 0 67896 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_738
timestamp 1623939100
transform 1 0 69000 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_750
timestamp 1623939100
transform 1 0 70104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _544_
timestamp 1623939100
transform 1 0 70380 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1233
timestamp 1623939100
transform 1 0 71944 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_762
timestamp 1623939100
transform 1 0 71208 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_771
timestamp 1623939100
transform 1 0 72036 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_783
timestamp 1623939100
transform 1 0 73140 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_795
timestamp 1623939100
transform 1 0 74244 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_807
timestamp 1623939100
transform 1 0 75348 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _430_
timestamp 1623939100
transform 1 0 77648 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1234
timestamp 1623939100
transform 1 0 77188 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_819
timestamp 1623939100
transform 1 0 76452 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_828
timestamp 1623939100
transform 1 0 77280 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_841
timestamp 1623939100
transform 1 0 78476 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_853
timestamp 1623939100
transform 1 0 79580 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_865
timestamp 1623939100
transform 1 0 80684 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1235
timestamp 1623939100
transform 1 0 82432 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_877
timestamp 1623939100
transform 1 0 81788 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_883
timestamp 1623939100
transform 1 0 82340 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_885
timestamp 1623939100
transform 1 0 82524 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_897
timestamp 1623939100
transform 1 0 83628 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_909
timestamp 1623939100
transform 1 0 84732 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_921
timestamp 1623939100
transform 1 0 85836 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_933
timestamp 1623939100
transform 1 0 86940 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1236
timestamp 1623939100
transform 1 0 87676 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_942
timestamp 1623939100
transform 1 0 87768 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_954
timestamp 1623939100
transform 1 0 88872 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_966
timestamp 1623939100
transform 1 0 89976 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_978
timestamp 1623939100
transform 1 0 91080 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1237
timestamp 1623939100
transform 1 0 92920 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_990
timestamp 1623939100
transform 1 0 92184 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_999
timestamp 1623939100
transform 1 0 93012 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _718_
timestamp 1623939100
transform -1 0 95128 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1623939100
transform -1 0 93380 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1022
timestamp 1623939100
transform 1 0 95128 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1034
timestamp 1623939100
transform 1 0 96232 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1623939100
transform -1 0 98808 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1238
timestamp 1623939100
transform 1 0 98164 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_1046
timestamp 1623939100
transform 1 0 97336 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1054
timestamp 1623939100
transform 1 0 98072 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_1056
timestamp 1623939100
transform 1 0 98256 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1623939100
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1623939100
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1623939100
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1623939100
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1623939100
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1623939100
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1257
timestamp 1623939100
transform 1 0 3772 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1623939100
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1623939100
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_27
timestamp 1623939100
transform 1 0 3588 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_30
timestamp 1623939100
transform 1 0 3864 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1239
timestamp 1623939100
transform 1 0 6348 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_51
timestamp 1623939100
transform 1 0 5796 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_58
timestamp 1623939100
transform 1 0 6440 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_42
timestamp 1623939100
transform 1 0 4968 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_54
timestamp 1623939100
transform 1 0 6072 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_70
timestamp 1623939100
transform 1 0 7544 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_82
timestamp 1623939100
transform 1 0 8648 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_66
timestamp 1623939100
transform 1 0 7176 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_78
timestamp 1623939100
transform 1 0 8280 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1258
timestamp 1623939100
transform 1 0 9016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_94
timestamp 1623939100
transform 1 0 9752 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_87
timestamp 1623939100
transform 1 0 9108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_99
timestamp 1623939100
transform 1 0 10212 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1240
timestamp 1623939100
transform 1 0 11592 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_106
timestamp 1623939100
transform 1 0 10856 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_115
timestamp 1623939100
transform 1 0 11684 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_111
timestamp 1623939100
transform 1 0 11316 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_123
timestamp 1623939100
transform 1 0 12420 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1259
timestamp 1623939100
transform 1 0 14260 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_127
timestamp 1623939100
transform 1 0 12788 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_139
timestamp 1623939100
transform 1 0 13892 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_135
timestamp 1623939100
transform 1 0 13524 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_144
timestamp 1623939100
transform 1 0 14352 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_151
timestamp 1623939100
transform 1 0 14996 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_163
timestamp 1623939100
transform 1 0 16100 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_156
timestamp 1623939100
transform 1 0 15456 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _555_
timestamp 1623939100
transform 1 0 17204 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1241
timestamp 1623939100
transform 1 0 16836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_172
timestamp 1623939100
transform 1 0 16928 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1623939100
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_168
timestamp 1623939100
transform 1 0 16560 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_174
timestamp 1623939100
transform 1 0 17112 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_178
timestamp 1623939100
transform 1 0 17480 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1260
timestamp 1623939100
transform 1 0 19504 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1623939100
transform 1 0 19136 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_208
timestamp 1623939100
transform 1 0 20240 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_190
timestamp 1623939100
transform 1 0 18584 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_198
timestamp 1623939100
transform 1 0 19320 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_201
timestamp 1623939100
transform 1 0 19596 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1242
timestamp 1623939100
transform 1 0 22080 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_220
timestamp 1623939100
transform 1 0 21344 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_229
timestamp 1623939100
transform 1 0 22172 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_213
timestamp 1623939100
transform 1 0 20700 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_225
timestamp 1623939100
transform 1 0 21804 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_241
timestamp 1623939100
transform 1 0 23276 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_237
timestamp 1623939100
transform 1 0 22908 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_249
timestamp 1623939100
transform 1 0 24012 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1261
timestamp 1623939100
transform 1 0 24748 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_253
timestamp 1623939100
transform 1 0 24380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_265
timestamp 1623939100
transform 1 0 25484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_258
timestamp 1623939100
transform 1 0 24840 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_270
timestamp 1623939100
transform 1 0 25944 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _676_
timestamp 1623939100
transform 1 0 27784 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1243
timestamp 1623939100
transform 1 0 27324 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_268
timestamp 1623939100
transform 1 0 27600 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_277
timestamp 1623939100
transform 1 0 26588 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_286
timestamp 1623939100
transform 1 0 27416 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_282
timestamp 1623939100
transform 1 0 27048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1623939100
transform 1 0 28060 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1623939100
transform 1 0 29164 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_294
timestamp 1623939100
transform 1 0 28152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_306
timestamp 1623939100
transform 1 0 29256 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1262
timestamp 1623939100
transform 1 0 29992 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1623939100
transform 1 0 30268 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_329
timestamp 1623939100
transform 1 0 31372 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_315
timestamp 1623939100
transform 1 0 30084 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_327
timestamp 1623939100
transform 1 0 31188 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1244
timestamp 1623939100
transform 1 0 32568 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_341
timestamp 1623939100
transform 1 0 32476 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_343
timestamp 1623939100
transform 1 0 32660 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_339
timestamp 1623939100
transform 1 0 32292 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_351
timestamp 1623939100
transform 1 0 33396 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _594_
timestamp 1623939100
transform 1 0 34592 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1263
timestamp 1623939100
transform 1 0 35236 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_305
timestamp 1623939100
transform 1 0 34408 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_355
timestamp 1623939100
transform 1 0 33764 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_361
timestamp 1623939100
transform 1 0 34316 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1623939100
transform 1 0 34868 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_363
timestamp 1623939100
transform 1 0 34500 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_372
timestamp 1623939100
transform 1 0 35328 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _677_
timestamp 1623939100
transform 1 0 36616 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_270
timestamp 1623939100
transform 1 0 36432 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_379
timestamp 1623939100
transform 1 0 35972 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_391
timestamp 1623939100
transform 1 0 37076 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1623939100
transform 1 0 36892 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _721_
timestamp 1623939100
transform 1 0 39376 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1245
timestamp 1623939100
transform 1 0 37812 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_400
timestamp 1623939100
transform 1 0 37904 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_412
timestamp 1623939100
transform 1 0 39008 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1623939100
transform 1 0 37996 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_413
timestamp 1623939100
transform 1 0 39100 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1264
timestamp 1623939100
transform 1 0 40480 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_433
timestamp 1623939100
transform 1 0 40940 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_425
timestamp 1623939100
transform 1 0 40204 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_429
timestamp 1623939100
transform 1 0 40572 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1246
timestamp 1623939100
transform 1 0 43056 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_445
timestamp 1623939100
transform 1 0 42044 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_453
timestamp 1623939100
transform 1 0 42780 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_457
timestamp 1623939100
transform 1 0 43148 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_441
timestamp 1623939100
transform 1 0 41676 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_453
timestamp 1623939100
transform 1 0 42780 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _371_
timestamp 1623939100
transform 1 0 43424 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_59_469
timestamp 1623939100
transform 1 0 44252 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_459
timestamp 1623939100
transform 1 0 43332 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_467
timestamp 1623939100
transform 1 0 44068 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_479
timestamp 1623939100
transform 1 0 45172 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _339_
timestamp 1623939100
transform 1 0 46736 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1265
timestamp 1623939100
transform 1 0 45724 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_481
timestamp 1623939100
transform 1 0 45356 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_493
timestamp 1623939100
transform 1 0 46460 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_486
timestamp 1623939100
transform 1 0 45816 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_494
timestamp 1623939100
transform 1 0 46552 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1247
timestamp 1623939100
transform 1 0 48300 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1623939100
transform 1 0 47564 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_514
timestamp 1623939100
transform 1 0 48392 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_504
timestamp 1623939100
transform 1 0 47472 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_516
timestamp 1623939100
transform 1 0 48576 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_526
timestamp 1623939100
transform 1 0 49496 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_538
timestamp 1623939100
transform 1 0 50600 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_528
timestamp 1623939100
transform 1 0 49680 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_540
timestamp 1623939100
transform 1 0 50784 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1266
timestamp 1623939100
transform 1 0 50968 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_550
timestamp 1623939100
transform 1 0 51704 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_562
timestamp 1623939100
transform 1 0 52808 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_543
timestamp 1623939100
transform 1 0 51060 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_555
timestamp 1623939100
transform 1 0 52164 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_4  _481_
timestamp 1623939100
transform 1 0 54096 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1248
timestamp 1623939100
transform 1 0 53544 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_571
timestamp 1623939100
transform 1 0 53636 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_583
timestamp 1623939100
transform 1 0 54740 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_567
timestamp 1623939100
transform 1 0 53268 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_575
timestamp 1623939100
transform 1 0 54004 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_581
timestamp 1623939100
transform 1 0 54556 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1267
timestamp 1623939100
transform 1 0 56212 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_595
timestamp 1623939100
transform 1 0 55844 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_593
timestamp 1623939100
transform 1 0 55660 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_600
timestamp 1623939100
transform 1 0 56304 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_607
timestamp 1623939100
transform 1 0 56948 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_619
timestamp 1623939100
transform 1 0 58052 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_612
timestamp 1623939100
transform 1 0 57408 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_624
timestamp 1623939100
transform 1 0 58512 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _354_
timestamp 1623939100
transform 1 0 59248 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1249
timestamp 1623939100
transform 1 0 58788 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_628
timestamp 1623939100
transform 1 0 58880 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_641
timestamp 1623939100
transform 1 0 60076 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_636
timestamp 1623939100
transform 1 0 59616 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _789_
timestamp 1623939100
transform 1 0 62008 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1268
timestamp 1623939100
transform 1 0 61456 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_125
timestamp 1623939100
transform 1 0 61824 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_653
timestamp 1623939100
transform 1 0 61180 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_665
timestamp 1623939100
transform 1 0 62284 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_648
timestamp 1623939100
transform 1 0 60720 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_657
timestamp 1623939100
transform 1 0 61548 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1250
timestamp 1623939100
transform 1 0 64032 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_677
timestamp 1623939100
transform 1 0 63388 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_683
timestamp 1623939100
transform 1 0 63940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_685
timestamp 1623939100
transform 1 0 64124 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_681
timestamp 1623939100
transform 1 0 63756 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_697
timestamp 1623939100
transform 1 0 65228 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_693
timestamp 1623939100
transform 1 0 64860 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_705
timestamp 1623939100
transform 1 0 65964 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_714
timestamp 1623939100
transform 1 0 66792 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_709
timestamp 1623939100
transform 1 0 66332 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_349
timestamp 1623939100
transform 1 0 67068 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1269
timestamp 1623939100
transform 1 0 66700 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_722
timestamp 1623939100
transform 1 0 67528 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_109
timestamp 1623939100
transform 1 0 67712 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_107
timestamp 1623939100
transform 1 0 67896 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _646_
timestamp 1623939100
transform 1 0 67252 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_722
timestamp 1623939100
transform 1 0 67528 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _421_
timestamp 1623939100
transform 1 0 68080 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1251
timestamp 1623939100
transform 1 0 69276 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_108
timestamp 1623939100
transform 1 0 69552 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_110
timestamp 1623939100
transform 1 0 69736 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_734
timestamp 1623939100
transform 1 0 68632 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_740
timestamp 1623939100
transform 1 0 69184 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_742
timestamp 1623939100
transform 1 0 69368 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_748
timestamp 1623939100
transform 1 0 69920 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1270
timestamp 1623939100
transform 1 0 71944 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_754
timestamp 1623939100
transform 1 0 70472 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_766
timestamp 1623939100
transform 1 0 71576 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_760
timestamp 1623939100
transform 1 0 71024 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_768
timestamp 1623939100
transform 1 0 71760 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _661_
timestamp 1623939100
transform 1 0 73784 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_364
timestamp 1623939100
transform 1 0 73600 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_778
timestamp 1623939100
transform 1 0 72680 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_786
timestamp 1623939100
transform 1 0 73416 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_771
timestamp 1623939100
transform 1 0 72036 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_783
timestamp 1623939100
transform 1 0 73140 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1252
timestamp 1623939100
transform 1 0 74520 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_793
timestamp 1623939100
transform 1 0 74060 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_797
timestamp 1623939100
transform 1 0 74428 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_799
timestamp 1623939100
transform 1 0 74612 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_811
timestamp 1623939100
transform 1 0 75716 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_795
timestamp 1623939100
transform 1 0 74244 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_807
timestamp 1623939100
transform 1 0 75348 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1271
timestamp 1623939100
transform 1 0 77188 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_823
timestamp 1623939100
transform 1 0 76820 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_819
timestamp 1623939100
transform 1 0 76452 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_828
timestamp 1623939100
transform 1 0 77280 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _288_
timestamp 1623939100
transform 1 0 78752 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_59_835
timestamp 1623939100
transform 1 0 77924 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_847
timestamp 1623939100
transform 1 0 79028 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_840
timestamp 1623939100
transform 1 0 78384 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_853
timestamp 1623939100
transform 1 0 79580 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _300_
timestamp 1623939100
transform 1 0 81604 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1253
timestamp 1623939100
transform 1 0 79764 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_856
timestamp 1623939100
transform 1 0 79856 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_868
timestamp 1623939100
transform 1 0 80960 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_874
timestamp 1623939100
transform 1 0 81512 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_865
timestamp 1623939100
transform 1 0 80684 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1272
timestamp 1623939100
transform 1 0 82432 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_884
timestamp 1623939100
transform 1 0 82432 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_877
timestamp 1623939100
transform 1 0 81788 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_883
timestamp 1623939100
transform 1 0 82340 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_885
timestamp 1623939100
transform 1 0 82524 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1254
timestamp 1623939100
transform 1 0 85008 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_896
timestamp 1623939100
transform 1 0 83536 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_908
timestamp 1623939100
transform 1 0 84640 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_913
timestamp 1623939100
transform 1 0 85100 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_897
timestamp 1623939100
transform 1 0 83628 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_909
timestamp 1623939100
transform 1 0 84732 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _452_
timestamp 1623939100
transform 1 0 86112 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_161
timestamp 1623939100
transform 1 0 85928 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_925
timestamp 1623939100
transform 1 0 86204 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_937
timestamp 1623939100
transform 1 0 87308 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_921
timestamp 1623939100
transform 1 0 85836 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_933
timestamp 1623939100
transform 1 0 86940 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1273
timestamp 1623939100
transform 1 0 87676 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_949
timestamp 1623939100
transform 1 0 88412 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_942
timestamp 1623939100
transform 1 0 87768 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_954
timestamp 1623939100
transform 1 0 88872 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1255
timestamp 1623939100
transform 1 0 90252 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_961
timestamp 1623939100
transform 1 0 89516 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_970
timestamp 1623939100
transform 1 0 90344 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_966
timestamp 1623939100
transform 1 0 89976 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_978
timestamp 1623939100
transform 1 0 91080 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1274
timestamp 1623939100
transform 1 0 92920 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_982
timestamp 1623939100
transform 1 0 91448 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_994
timestamp 1623939100
transform 1 0 92552 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_990
timestamp 1623939100
transform 1 0 92184 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_999
timestamp 1623939100
transform 1 0 93012 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _539_
timestamp 1623939100
transform 1 0 95036 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _566_
timestamp 1623939100
transform 1 0 94392 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_248
timestamp 1623939100
transform 1 0 94208 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1006
timestamp 1623939100
transform 1 0 93656 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1017
timestamp 1623939100
transform 1 0 94668 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_1011
timestamp 1623939100
transform 1 0 94116 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_1019
timestamp 1623939100
transform 1 0 94852 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1256
timestamp 1623939100
transform 1 0 95496 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1025
timestamp 1623939100
transform 1 0 95404 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1027
timestamp 1623939100
transform 1 0 95588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1039
timestamp 1623939100
transform 1 0 96692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1030
timestamp 1623939100
transform 1 0 95864 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1623939100
transform -1 0 98808 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1623939100
transform -1 0 98808 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1275
timestamp 1623939100
transform 1 0 98164 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1051
timestamp 1623939100
transform 1 0 97796 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1042
timestamp 1623939100
transform 1 0 96968 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1054
timestamp 1623939100
transform 1 0 98072 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_1056
timestamp 1623939100
transform 1 0 98256 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1623939100
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1623939100
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1623939100
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1623939100
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1623939100
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1276
timestamp 1623939100
transform 1 0 6348 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_51
timestamp 1623939100
transform 1 0 5796 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_58
timestamp 1623939100
transform 1 0 6440 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_70
timestamp 1623939100
transform 1 0 7544 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_82
timestamp 1623939100
transform 1 0 8648 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_94
timestamp 1623939100
transform 1 0 9752 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1277
timestamp 1623939100
transform 1 0 11592 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_106
timestamp 1623939100
transform 1 0 10856 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_115
timestamp 1623939100
transform 1 0 11684 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_127
timestamp 1623939100
transform 1 0 12788 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_139
timestamp 1623939100
transform 1 0 13892 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_151
timestamp 1623939100
transform 1 0 14996 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_163
timestamp 1623939100
transform 1 0 16100 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1278
timestamp 1623939100
transform 1 0 16836 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_172
timestamp 1623939100
transform 1 0 16928 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_184
timestamp 1623939100
transform 1 0 18032 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _674_
timestamp 1623939100
transform 1 0 18952 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_264
timestamp 1623939100
transform 1 0 18768 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_197
timestamp 1623939100
transform 1 0 19228 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1279
timestamp 1623939100
transform 1 0 22080 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_209
timestamp 1623939100
transform 1 0 20332 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_221
timestamp 1623939100
transform 1 0 21436 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_227
timestamp 1623939100
transform 1 0 21988 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_229
timestamp 1623939100
transform 1 0 22172 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_241
timestamp 1623939100
transform 1 0 23276 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_249
timestamp 1623939100
transform 1 0 24012 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_4  _414_
timestamp 1623939100
transform 1 0 24196 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_61_265
timestamp 1623939100
transform 1 0 25484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1280
timestamp 1623939100
transform 1 0 27324 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_277
timestamp 1623939100
transform 1 0 26588 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_286
timestamp 1623939100
transform 1 0 27416 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_298
timestamp 1623939100
transform 1 0 28520 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_310
timestamp 1623939100
transform 1 0 29624 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_322
timestamp 1623939100
transform 1 0 30728 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1281
timestamp 1623939100
transform 1 0 32568 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_334
timestamp 1623939100
transform 1 0 31832 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_343
timestamp 1623939100
transform 1 0 32660 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_355
timestamp 1623939100
transform 1 0 33764 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1623939100
transform 1 0 34868 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1623939100
transform 1 0 35972 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_391
timestamp 1623939100
transform 1 0 37076 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1282
timestamp 1623939100
transform 1 0 37812 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_93
timestamp 1623939100
transform 1 0 39376 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_400
timestamp 1623939100
transform 1 0 37904 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_412
timestamp 1623939100
transform 1 0 39008 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _752_
timestamp 1623939100
transform 1 0 39560 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_61_437
timestamp 1623939100
transform 1 0 41308 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1283
timestamp 1623939100
transform 1 0 43056 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_449
timestamp 1623939100
transform 1 0 42412 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_455
timestamp 1623939100
transform 1 0 42964 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_457
timestamp 1623939100
transform 1 0 43148 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_469
timestamp 1623939100
transform 1 0 44252 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_481
timestamp 1623939100
transform 1 0 45356 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_493
timestamp 1623939100
transform 1 0 46460 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1284
timestamp 1623939100
transform 1 0 48300 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1623939100
transform 1 0 47564 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_514
timestamp 1623939100
transform 1 0 48392 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_526
timestamp 1623939100
transform 1 0 49496 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_538
timestamp 1623939100
transform 1 0 50600 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_550
timestamp 1623939100
transform 1 0 51704 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_562
timestamp 1623939100
transform 1 0 52808 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1285
timestamp 1623939100
transform 1 0 53544 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_571
timestamp 1623939100
transform 1 0 53636 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_583
timestamp 1623939100
transform 1 0 54740 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _714_
timestamp 1623939100
transform 1 0 55660 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_61_591
timestamp 1623939100
transform 1 0 55476 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_612
timestamp 1623939100
transform 1 0 57408 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_624
timestamp 1623939100
transform 1 0 58512 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1286
timestamp 1623939100
transform 1 0 58788 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_628
timestamp 1623939100
transform 1 0 58880 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_640
timestamp 1623939100
transform 1 0 59984 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_652
timestamp 1623939100
transform 1 0 61088 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_664
timestamp 1623939100
transform 1 0 62192 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1287
timestamp 1623939100
transform 1 0 64032 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_676
timestamp 1623939100
transform 1 0 63296 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_685
timestamp 1623939100
transform 1 0 64124 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_697
timestamp 1623939100
transform 1 0 65228 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_709
timestamp 1623939100
transform 1 0 66332 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_721
timestamp 1623939100
transform 1 0 67436 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1288
timestamp 1623939100
transform 1 0 69276 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_733
timestamp 1623939100
transform 1 0 68540 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_742
timestamp 1623939100
transform 1 0 69368 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_754
timestamp 1623939100
transform 1 0 70472 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_766
timestamp 1623939100
transform 1 0 71576 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_778
timestamp 1623939100
transform 1 0 72680 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_790
timestamp 1623939100
transform 1 0 73784 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1289
timestamp 1623939100
transform 1 0 74520 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_799
timestamp 1623939100
transform 1 0 74612 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_811
timestamp 1623939100
transform 1 0 75716 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_823
timestamp 1623939100
transform 1 0 76820 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_835
timestamp 1623939100
transform 1 0 77924 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_847
timestamp 1623939100
transform 1 0 79028 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1290
timestamp 1623939100
transform 1 0 79764 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_856
timestamp 1623939100
transform 1 0 79856 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_868
timestamp 1623939100
transform 1 0 80960 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _441_
timestamp 1623939100
transform 1 0 81880 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_61_876
timestamp 1623939100
transform 1 0 81696 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_887
timestamp 1623939100
transform 1 0 82708 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1291
timestamp 1623939100
transform 1 0 85008 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_899
timestamp 1623939100
transform 1 0 83812 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_911
timestamp 1623939100
transform 1 0 84916 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_913
timestamp 1623939100
transform 1 0 85100 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_925
timestamp 1623939100
transform 1 0 86204 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_937
timestamp 1623939100
transform 1 0 87308 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_949
timestamp 1623939100
transform 1 0 88412 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1292
timestamp 1623939100
transform 1 0 90252 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_961
timestamp 1623939100
transform 1 0 89516 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_970
timestamp 1623939100
transform 1 0 90344 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_982
timestamp 1623939100
transform 1 0 91448 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_994
timestamp 1623939100
transform 1 0 92552 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1006
timestamp 1623939100
transform 1 0 93656 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1018
timestamp 1623939100
transform 1 0 94760 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1293
timestamp 1623939100
transform 1 0 95496 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1027
timestamp 1623939100
transform 1 0 95588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1039
timestamp 1623939100
transform 1 0 96692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1623939100
transform -1 0 98808 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1051
timestamp 1623939100
transform 1 0 97796 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1623939100
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1623939100
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1623939100
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1294
timestamp 1623939100
transform 1 0 3772 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_27
timestamp 1623939100
transform 1 0 3588 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_30
timestamp 1623939100
transform 1 0 3864 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _449_
timestamp 1623939100
transform 1 0 5244 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_62_42
timestamp 1623939100
transform 1 0 4968 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_61
timestamp 1623939100
transform 1 0 6716 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_73
timestamp 1623939100
transform 1 0 7820 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1295
timestamp 1623939100
transform 1 0 9016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_85
timestamp 1623939100
transform 1 0 8924 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_87
timestamp 1623939100
transform 1 0 9108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_99
timestamp 1623939100
transform 1 0 10212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_111
timestamp 1623939100
transform 1 0 11316 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_123
timestamp 1623939100
transform 1 0 12420 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _495_
timestamp 1623939100
transform 1 0 12880 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1296
timestamp 1623939100
transform 1 0 14260 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_127
timestamp 1623939100
transform 1 0 12788 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_137
timestamp 1623939100
transform 1 0 13708 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_144
timestamp 1623939100
transform 1 0 14352 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_156
timestamp 1623939100
transform 1 0 15456 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_356
timestamp 1623939100
transform 1 0 18308 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_168
timestamp 1623939100
transform 1 0 16560 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_180
timestamp 1623939100
transform 1 0 17664 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_186
timestamp 1623939100
transform 1 0 18216 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _655_
timestamp 1623939100
transform 1 0 18492 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1297
timestamp 1623939100
transform 1 0 19504 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_192
timestamp 1623939100
transform 1 0 18768 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_201
timestamp 1623939100
transform 1 0 19596 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_213
timestamp 1623939100
transform 1 0 20700 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_225
timestamp 1623939100
transform 1 0 21804 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_237
timestamp 1623939100
transform 1 0 22908 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_249
timestamp 1623939100
transform 1 0 24012 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1298
timestamp 1623939100
transform 1 0 24748 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_258
timestamp 1623939100
transform 1 0 24840 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_270
timestamp 1623939100
transform 1 0 25944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_4  _458_
timestamp 1623939100
transform 1 0 27416 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_62_282
timestamp 1623939100
transform 1 0 27048 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_302
timestamp 1623939100
transform 1 0 28888 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1299
timestamp 1623939100
transform 1 0 29992 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_315
timestamp 1623939100
transform 1 0 30084 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_327
timestamp 1623939100
transform 1 0 31188 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_339
timestamp 1623939100
transform 1 0 32292 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_351
timestamp 1623939100
transform 1 0 33396 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1300
timestamp 1623939100
transform 1 0 35236 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_363
timestamp 1623939100
transform 1 0 34500 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_372
timestamp 1623939100
transform 1 0 35328 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _694_
timestamp 1623939100
transform 1 0 37260 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_289
timestamp 1623939100
transform 1 0 37076 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_384
timestamp 1623939100
transform 1 0 36432 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_390
timestamp 1623939100
transform 1 0 36984 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_396
timestamp 1623939100
transform 1 0 37536 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_408
timestamp 1623939100
transform 1 0 38640 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1301
timestamp 1623939100
transform 1 0 40480 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_420
timestamp 1623939100
transform 1 0 39744 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_429
timestamp 1623939100
transform 1 0 40572 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_441
timestamp 1623939100
transform 1 0 41676 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_453
timestamp 1623939100
transform 1 0 42780 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_465
timestamp 1623939100
transform 1 0 43884 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_477
timestamp 1623939100
transform 1 0 44988 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1302
timestamp 1623939100
transform 1 0 45724 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1623939100
transform 1 0 47012 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_486
timestamp 1623939100
transform 1 0 45816 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_498
timestamp 1623939100
transform 1 0 46920 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _728_
timestamp 1623939100
transform 1 0 47196 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_520
timestamp 1623939100
transform 1 0 48944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_532
timestamp 1623939100
transform 1 0 50048 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_540
timestamp 1623939100
transform 1 0 50784 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_6  _459_
timestamp 1623939100
transform 1 0 52072 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1303
timestamp 1623939100
transform 1 0 50968 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_543
timestamp 1623939100
transform 1 0 51060 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_551
timestamp 1623939100
transform 1 0 51796 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_563
timestamp 1623939100
transform 1 0 52900 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_575
timestamp 1623939100
transform 1 0 54004 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_583
timestamp 1623939100
transform 1 0 54740 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _457_
timestamp 1623939100
transform 1 0 54832 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1304
timestamp 1623939100
transform 1 0 56212 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_593
timestamp 1623939100
transform 1 0 55660 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_600
timestamp 1623939100
transform 1 0 56304 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_612
timestamp 1623939100
transform 1 0 57408 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_624
timestamp 1623939100
transform 1 0 58512 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_636
timestamp 1623939100
transform 1 0 59616 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1305
timestamp 1623939100
transform 1 0 61456 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_648
timestamp 1623939100
transform 1 0 60720 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_657
timestamp 1623939100
transform 1 0 61548 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _730_
timestamp 1623939100
transform 1 0 63112 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_62_669
timestamp 1623939100
transform 1 0 62652 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_673
timestamp 1623939100
transform 1 0 63020 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output422
timestamp 1623939100
transform 1 0 65228 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_693
timestamp 1623939100
transform 1 0 64860 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_701
timestamp 1623939100
transform 1 0 65596 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1306
timestamp 1623939100
transform 1 0 66700 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_714
timestamp 1623939100
transform 1 0 66792 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_726
timestamp 1623939100
transform 1 0 67896 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_738
timestamp 1623939100
transform 1 0 69000 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_750
timestamp 1623939100
transform 1 0 70104 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1307
timestamp 1623939100
transform 1 0 71944 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_762
timestamp 1623939100
transform 1 0 71208 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _543_
timestamp 1623939100
transform 1 0 73876 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_771
timestamp 1623939100
transform 1 0 72036 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_783
timestamp 1623939100
transform 1 0 73140 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_800
timestamp 1623939100
transform 1 0 74704 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_812
timestamp 1623939100
transform 1 0 75808 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1308
timestamp 1623939100
transform 1 0 77188 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_824
timestamp 1623939100
transform 1 0 76912 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_828
timestamp 1623939100
transform 1 0 77280 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_840
timestamp 1623939100
transform 1 0 78384 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_852
timestamp 1623939100
transform 1 0 79488 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_864
timestamp 1623939100
transform 1 0 80592 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1309
timestamp 1623939100
transform 1 0 82432 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_876
timestamp 1623939100
transform 1 0 81696 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_885
timestamp 1623939100
transform 1 0 82524 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_897
timestamp 1623939100
transform 1 0 83628 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_909
timestamp 1623939100
transform 1 0 84732 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_921
timestamp 1623939100
transform 1 0 85836 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_933
timestamp 1623939100
transform 1 0 86940 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1310
timestamp 1623939100
transform 1 0 87676 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_942
timestamp 1623939100
transform 1 0 87768 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_954
timestamp 1623939100
transform 1 0 88872 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_966
timestamp 1623939100
transform 1 0 89976 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_978
timestamp 1623939100
transform 1 0 91080 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1311
timestamp 1623939100
transform 1 0 92920 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_990
timestamp 1623939100
transform 1 0 92184 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_999
timestamp 1623939100
transform 1 0 93012 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _475_
timestamp 1623939100
transform 1 0 93380 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1623939100
transform 1 0 95036 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1012
timestamp 1623939100
transform 1 0 94208 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1020
timestamp 1623939100
transform 1 0 94944 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1024
timestamp 1623939100
transform 1 0 95312 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1036
timestamp 1623939100
transform 1 0 96416 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1623939100
transform -1 0 98808 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1312
timestamp 1623939100
transform 1 0 98164 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1623939100
transform 1 0 97520 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1051
timestamp 1623939100
transform 1 0 97796 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_1056
timestamp 1623939100
transform 1 0 98256 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _708_
timestamp 1623939100
transform 1 0 2944 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1623939100
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output406
timestamp 1623939100
transform -1 0 2484 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_227
timestamp 1623939100
transform -1 0 2116 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_3
timestamp 1623939100
transform 1 0 1380 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1623939100
transform 1 0 2484 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_19
timestamp 1623939100
transform 1 0 2852 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1623939100
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1313
timestamp 1623939100
transform 1 0 6348 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_51
timestamp 1623939100
transform 1 0 5796 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_58
timestamp 1623939100
transform 1 0 6440 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1623939100
transform 1 0 8188 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output428
timestamp 1623939100
transform 1 0 7360 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_66
timestamp 1623939100
transform 1 0 7176 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_72
timestamp 1623939100
transform 1 0 7728 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_76
timestamp 1623939100
transform 1 0 8096 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_80
timestamp 1623939100
transform 1 0 8464 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output437
timestamp 1623939100
transform 1 0 9936 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_92
timestamp 1623939100
transform 1 0 9568 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_100
timestamp 1623939100
transform 1 0 10304 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1314
timestamp 1623939100
transform 1 0 11592 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output438
timestamp 1623939100
transform 1 0 12604 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_112
timestamp 1623939100
transform 1 0 11408 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_115
timestamp 1623939100
transform 1 0 11684 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_123
timestamp 1623939100
transform 1 0 12420 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_129
timestamp 1623939100
transform 1 0 12972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_141
timestamp 1623939100
transform 1 0 14076 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output439
timestamp 1623939100
transform 1 0 15272 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_153
timestamp 1623939100
transform 1 0 15180 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_158
timestamp 1623939100
transform 1 0 15640 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1315
timestamp 1623939100
transform 1 0 16836 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output440
timestamp 1623939100
transform -1 0 18216 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_244
timestamp 1623939100
transform -1 0 17848 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_170
timestamp 1623939100
transform 1 0 16744 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_172
timestamp 1623939100
transform 1 0 16928 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_186
timestamp 1623939100
transform 1 0 18216 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _480_
timestamp 1623939100
transform -1 0 19596 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_153
timestamp 1623939100
transform -1 0 18768 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_201
timestamp 1623939100
transform 1 0 19596 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1316
timestamp 1623939100
transform 1 0 22080 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output441
timestamp 1623939100
transform 1 0 20516 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_209
timestamp 1623939100
transform 1 0 20332 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_215
timestamp 1623939100
transform 1 0 20884 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_227
timestamp 1623939100
transform 1 0 21988 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_229
timestamp 1623939100
transform 1 0 22172 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_241
timestamp 1623939100
transform 1 0 23276 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_253
timestamp 1623939100
transform 1 0 24380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_265
timestamp 1623939100
transform 1 0 25484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1317
timestamp 1623939100
transform 1 0 27324 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1623939100
transform 1 0 26680 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_277
timestamp 1623939100
transform 1 0 26588 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_281
timestamp 1623939100
transform 1 0 26956 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_286
timestamp 1623939100
transform 1 0 27416 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _297_
timestamp 1623939100
transform 1 0 28520 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1623939100
transform 1 0 29716 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_307
timestamp 1623939100
transform 1 0 29348 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _666_
timestamp 1623939100
transform 1 0 31464 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_373
timestamp 1623939100
transform 1 0 31280 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_314
timestamp 1623939100
transform 1 0 29992 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_326
timestamp 1623939100
transform 1 0 31096 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_333
timestamp 1623939100
transform 1 0 31740 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1318
timestamp 1623939100
transform 1 0 32568 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output409
timestamp 1623939100
transform 1 0 33672 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_341
timestamp 1623939100
transform 1 0 32476 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_343
timestamp 1623939100
transform 1 0 32660 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_351
timestamp 1623939100
transform 1 0 33396 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_358
timestamp 1623939100
transform 1 0 34040 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_370
timestamp 1623939100
transform 1 0 35144 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output410
timestamp 1623939100
transform 1 0 36248 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_386
timestamp 1623939100
transform 1 0 36616 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1319
timestamp 1623939100
transform 1 0 37812 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_398
timestamp 1623939100
transform 1 0 37720 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_400
timestamp 1623939100
transform 1 0 37904 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_412
timestamp 1623939100
transform 1 0 39008 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_424
timestamp 1623939100
transform 1 0 40112 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_436
timestamp 1623939100
transform 1 0 41216 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1320
timestamp 1623939100
transform 1 0 43056 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1623939100
transform 1 0 42412 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_448
timestamp 1623939100
transform 1 0 42320 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_452
timestamp 1623939100
transform 1 0 42688 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_457
timestamp 1623939100
transform 1 0 43148 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _754_
timestamp 1623939100
transform 1 0 43516 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_2  output414
timestamp 1623939100
transform 1 0 46828 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_480
timestamp 1623939100
transform 1 0 45264 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_492
timestamp 1623939100
transform 1 0 46368 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_496
timestamp 1623939100
transform 1 0 46736 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1321
timestamp 1623939100
transform 1 0 48300 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_501
timestamp 1623939100
transform 1 0 47196 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_514
timestamp 1623939100
transform 1 0 48392 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_526
timestamp 1623939100
transform 1 0 49496 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_538
timestamp 1623939100
transform 1 0 50600 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_550
timestamp 1623939100
transform 1 0 51704 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_562
timestamp 1623939100
transform 1 0 52808 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1322
timestamp 1623939100
transform 1 0 53544 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output418
timestamp 1623939100
transform 1 0 54740 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_571
timestamp 1623939100
transform 1 0 53636 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _607_
timestamp 1623939100
transform -1 0 55752 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1623939100
transform 1 0 56120 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_313
timestamp 1623939100
transform -1 0 55476 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_587
timestamp 1623939100
transform 1 0 55108 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_594
timestamp 1623939100
transform 1 0 55752 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_601
timestamp 1623939100
transform 1 0 56396 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output419
timestamp 1623939100
transform 1 0 57316 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_609
timestamp 1623939100
transform 1 0 57132 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_615
timestamp 1623939100
transform 1 0 57684 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1323
timestamp 1623939100
transform 1 0 58788 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output420
timestamp 1623939100
transform 1 0 59984 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_628
timestamp 1623939100
transform 1 0 58880 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_644
timestamp 1623939100
transform 1 0 60352 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_656
timestamp 1623939100
transform 1 0 61456 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1324
timestamp 1623939100
transform 1 0 64032 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output421
timestamp 1623939100
transform 1 0 62560 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_672
timestamp 1623939100
transform 1 0 62928 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_685
timestamp 1623939100
transform 1 0 64124 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _451_
timestamp 1623939100
transform 1 0 65320 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_63_697
timestamp 1623939100
transform 1 0 65228 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_707
timestamp 1623939100
transform 1 0 66148 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output423
timestamp 1623939100
transform 1 0 67896 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_719
timestamp 1623939100
transform 1 0 67252 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_725
timestamp 1623939100
transform 1 0 67804 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _599_
timestamp 1623939100
transform -1 0 68908 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1325
timestamp 1623939100
transform 1 0 69276 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_307
timestamp 1623939100
transform -1 0 68632 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_730
timestamp 1623939100
transform 1 0 68264 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_737
timestamp 1623939100
transform 1 0 68908 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_742
timestamp 1623939100
transform 1 0 69368 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output424
timestamp 1623939100
transform 1 0 70472 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_758
timestamp 1623939100
transform 1 0 70840 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_770
timestamp 1623939100
transform 1 0 71944 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _392_
timestamp 1623939100
transform 1 0 73508 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output425
timestamp 1623939100
transform 1 0 72772 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_778
timestamp 1623939100
transform 1 0 72680 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_783
timestamp 1623939100
transform 1 0 73140 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1326
timestamp 1623939100
transform 1 0 74520 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output426
timestamp 1623939100
transform 1 0 75808 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_793
timestamp 1623939100
transform 1 0 74060 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_797
timestamp 1623939100
transform 1 0 74428 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_799
timestamp 1623939100
transform 1 0 74612 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_811
timestamp 1623939100
transform 1 0 75716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_816
timestamp 1623939100
transform 1 0 76176 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_828
timestamp 1623939100
transform 1 0 77280 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1623939100
transform 1 0 79120 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output427
timestamp 1623939100
transform 1 0 78384 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_844
timestamp 1623939100
transform 1 0 78752 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_851
timestamp 1623939100
transform 1 0 79396 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1327
timestamp 1623939100
transform 1 0 79764 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_856
timestamp 1623939100
transform 1 0 79856 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_868
timestamp 1623939100
transform 1 0 80960 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_880
timestamp 1623939100
transform 1 0 82064 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_892
timestamp 1623939100
transform 1 0 83168 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1328
timestamp 1623939100
transform 1 0 85008 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1623939100
transform 1 0 84364 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_904
timestamp 1623939100
transform 1 0 84272 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_908
timestamp 1623939100
transform 1 0 84640 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_913
timestamp 1623939100
transform 1 0 85100 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1623939100
transform 1 0 87124 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_925
timestamp 1623939100
transform 1 0 86204 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_933
timestamp 1623939100
transform 1 0 86940 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_938
timestamp 1623939100
transform 1 0 87400 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_950
timestamp 1623939100
transform 1 0 88504 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1329
timestamp 1623939100
transform 1 0 90252 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1623939100
transform 1 0 89608 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_965
timestamp 1623939100
transform 1 0 89884 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_970
timestamp 1623939100
transform 1 0 90344 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1623939100
transform 1 0 92460 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_982
timestamp 1623939100
transform 1 0 91448 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_990
timestamp 1623939100
transform 1 0 92184 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_996
timestamp 1623939100
transform 1 0 92736 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output434
timestamp 1623939100
transform -1 0 94576 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_238
timestamp 1623939100
transform -1 0 94208 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1008
timestamp 1623939100
transform 1 0 93840 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1016
timestamp 1623939100
transform 1 0 94576 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1330
timestamp 1623939100
transform 1 0 95496 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output435
timestamp 1623939100
transform -1 0 97152 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_239
timestamp 1623939100
transform -1 0 96784 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1024
timestamp 1623939100
transform 1 0 95312 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1027
timestamp 1623939100
transform 1 0 95588 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_1035
timestamp 1623939100
transform 1 0 96324 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1623939100
transform -1 0 98808 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output436
timestamp 1623939100
transform 1 0 97796 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_241
timestamp 1623939100
transform 1 0 97612 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_242
timestamp 1623939100
transform 1 0 98164 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1044
timestamp 1623939100
transform 1 0 97152 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1048
timestamp 1623939100
transform 1 0 97520 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1057
timestamp 1623939100
transform 1 0 98348 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1623939100
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1623939100
transform 1 0 1748 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1623939100
transform 1 0 2944 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_180
timestamp 1623939100
transform 1 0 1564 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_181
timestamp 1623939100
transform 1 0 2300 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1623939100
transform 1 0 1380 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1623939100
transform 1 0 2484 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_19
timestamp 1623939100
transform 1 0 2852 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1331
timestamp 1623939100
transform 1 0 3772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output368
timestamp 1623939100
transform 1 0 4232 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1623939100
transform 1 0 3312 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_28
timestamp 1623939100
transform 1 0 3680 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_30
timestamp 1623939100
transform 1 0 3864 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_38
timestamp 1623939100
transform 1 0 4600 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1332
timestamp 1623939100
transform 1 0 6440 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  input23
timestamp 1623939100
transform 1 0 5244 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_64_44
timestamp 1623939100
transform 1 0 5152 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_54
timestamp 1623939100
transform 1 0 6072 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_59
timestamp 1623939100
transform 1 0 6532 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output379
timestamp 1623939100
transform 1 0 6900 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output390
timestamp 1623939100
transform 1 0 7636 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output417
timestamp 1623939100
transform 1 0 8372 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_67
timestamp 1623939100
transform 1 0 7268 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_75
timestamp 1623939100
transform 1 0 8004 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_83
timestamp 1623939100
transform 1 0 8740 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1333
timestamp 1623939100
transform 1 0 9108 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output399
timestamp 1623939100
transform -1 0 9936 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_222
timestamp 1623939100
transform -1 0 9568 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_88
timestamp 1623939100
transform 1 0 9200 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_96
timestamp 1623939100
transform 1 0 9936 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_104
timestamp 1623939100
transform 1 0 10672 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1334
timestamp 1623939100
transform 1 0 11776 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input33
timestamp 1623939100
transform 1 0 10856 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output400
timestamp 1623939100
transform 1 0 12236 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_110
timestamp 1623939100
transform 1 0 11224 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_117
timestamp 1623939100
transform 1 0 11868 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_125
timestamp 1623939100
transform 1 0 12604 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1335
timestamp 1623939100
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input34
timestamp 1623939100
transform 1 0 13524 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_133
timestamp 1623939100
transform 1 0 13340 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1623939100
transform 1 0 14076 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input35
timestamp 1623939100
transform 1 0 16100 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output401
timestamp 1623939100
transform -1 0 15272 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_224
timestamp 1623939100
transform -1 0 14904 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_146
timestamp 1623939100
transform 1 0 14536 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_154
timestamp 1623939100
transform 1 0 15272 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_162
timestamp 1623939100
transform 1 0 16008 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1336
timestamp 1623939100
transform 1 0 17112 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output402
timestamp 1623939100
transform 1 0 17572 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_169
timestamp 1623939100
transform 1 0 16652 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_173
timestamp 1623939100
transform 1 0 17020 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_175
timestamp 1623939100
transform 1 0 17204 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_183
timestamp 1623939100
transform 1 0 17940 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1337
timestamp 1623939100
transform 1 0 19780 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input36
timestamp 1623939100
transform 1 0 18768 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output403
timestamp 1623939100
transform 1 0 20240 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_191
timestamp 1623939100
transform 1 0 18676 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_198
timestamp 1623939100
transform 1 0 19320 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_202
timestamp 1623939100
transform 1 0 19688 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_204
timestamp 1623939100
transform 1 0 19872 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1623939100
transform 1 0 21344 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_212
timestamp 1623939100
transform 1 0 20608 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_224
timestamp 1623939100
transform 1 0 21712 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1338
timestamp 1623939100
transform 1 0 22448 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623939100
transform 1 0 23828 0 -1 37536
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  output404
timestamp 1623939100
transform 1 0 22908 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_233
timestamp 1623939100
transform 1 0 22540 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_241
timestamp 1623939100
transform 1 0 23276 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1339
timestamp 1623939100
transform 1 0 25116 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output405
timestamp 1623939100
transform 1 0 25576 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_257
timestamp 1623939100
transform 1 0 24748 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_262
timestamp 1623939100
transform 1 0 25208 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_270
timestamp 1623939100
transform 1 0 25944 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1340
timestamp 1623939100
transform 1 0 27784 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output442
timestamp 1623939100
transform -1 0 26680 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output443
timestamp 1623939100
transform 1 0 27048 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_247
timestamp 1623939100
transform -1 0 26312 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_278
timestamp 1623939100
transform 1 0 26680 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1623939100
transform 1 0 27416 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_291
timestamp 1623939100
transform 1 0 27876 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output369
timestamp 1623939100
transform 1 0 28244 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output407
timestamp 1623939100
transform 1 0 28980 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output408
timestamp 1623939100
transform 1 0 29716 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_299
timestamp 1623939100
transform 1 0 28612 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_307
timestamp 1623939100
transform 1 0 29348 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1341
timestamp 1623939100
transform 1 0 30452 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output370
timestamp 1623939100
transform 1 0 30912 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1623939100
transform 1 0 30084 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_320
timestamp 1623939100
transform 1 0 30544 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_328
timestamp 1623939100
transform 1 0 31280 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1342
timestamp 1623939100
transform 1 0 33120 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1623939100
transform 1 0 31924 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output371
timestamp 1623939100
transform 1 0 33580 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_334
timestamp 1623939100
transform 1 0 31832 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_339
timestamp 1623939100
transform 1 0 32292 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_347
timestamp 1623939100
transform 1 0 33028 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_349
timestamp 1623939100
transform 1 0 33212 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1623939100
transform 1 0 34500 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1623939100
transform 1 0 33948 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_367
timestamp 1623939100
transform 1 0 34868 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_375
timestamp 1623939100
transform 1 0 35604 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1343
timestamp 1623939100
transform 1 0 35788 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1623939100
transform 1 0 37168 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output372
timestamp 1623939100
transform 1 0 36248 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_378
timestamp 1623939100
transform 1 0 35880 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_386
timestamp 1623939100
transform 1 0 36616 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1344
timestamp 1623939100
transform 1 0 38456 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output373
timestamp 1623939100
transform 1 0 38916 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_396
timestamp 1623939100
transform 1 0 37536 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_404
timestamp 1623939100
transform 1 0 38272 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_407
timestamp 1623939100
transform 1 0 38548 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_415
timestamp 1623939100
transform 1 0 39284 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1345
timestamp 1623939100
transform 1 0 41124 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1623939100
transform 1 0 39836 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_425
timestamp 1623939100
transform 1 0 40204 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_433
timestamp 1623939100
transform 1 0 40940 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_436
timestamp 1623939100
transform 1 0 41216 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output374
timestamp 1623939100
transform 1 0 41584 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output375
timestamp 1623939100
transform 1 0 43056 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output411
timestamp 1623939100
transform 1 0 42320 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_444
timestamp 1623939100
transform 1 0 41952 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_452
timestamp 1623939100
transform 1 0 42688 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1346
timestamp 1623939100
transform 1 0 43792 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1623939100
transform 1 0 45080 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output412
timestamp 1623939100
transform 1 0 44252 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_460
timestamp 1623939100
transform 1 0 43424 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_465
timestamp 1623939100
transform 1 0 43884 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_473
timestamp 1623939100
transform 1 0 44620 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_477
timestamp 1623939100
transform 1 0 44988 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1347
timestamp 1623939100
transform 1 0 46460 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output376
timestamp 1623939100
transform 1 0 46920 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_482
timestamp 1623939100
transform 1 0 45448 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_490
timestamp 1623939100
transform 1 0 46184 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_494
timestamp 1623939100
transform 1 0 46552 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1623939100
transform 1 0 47656 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output377
timestamp 1623939100
transform 1 0 48392 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_502
timestamp 1623939100
transform 1 0 47288 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_510
timestamp 1623939100
transform 1 0 48024 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_518
timestamp 1623939100
transform 1 0 48760 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1348
timestamp 1623939100
transform 1 0 49128 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1623939100
transform 1 0 50324 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output413
timestamp 1623939100
transform 1 0 49588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_523
timestamp 1623939100
transform 1 0 49220 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_531
timestamp 1623939100
transform 1 0 49956 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_539
timestamp 1623939100
transform 1 0 50692 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1349
timestamp 1623939100
transform 1 0 51796 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output378
timestamp 1623939100
transform 1 0 51060 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output415
timestamp 1623939100
transform 1 0 52256 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_547
timestamp 1623939100
transform 1 0 51428 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_552
timestamp 1623939100
transform 1 0 51888 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_560
timestamp 1623939100
transform 1 0 52624 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1350
timestamp 1623939100
transform 1 0 54464 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input13
timestamp 1623939100
transform 1 0 52992 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_570
timestamp 1623939100
transform 1 0 53544 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_578
timestamp 1623939100
transform 1 0 54280 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_581
timestamp 1623939100
transform 1 0 54556 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output380
timestamp 1623939100
transform 1 0 54924 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output381
timestamp 1623939100
transform 1 0 56396 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output416
timestamp 1623939100
transform 1 0 55660 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_589
timestamp 1623939100
transform 1 0 55292 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_597
timestamp 1623939100
transform 1 0 56028 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _429_
timestamp 1623939100
transform 1 0 58328 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1351
timestamp 1623939100
transform 1 0 57132 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1623939100
transform 1 0 57592 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_605
timestamp 1623939100
transform 1 0 56764 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_610
timestamp 1623939100
transform 1 0 57224 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_618
timestamp 1623939100
transform 1 0 57960 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1352
timestamp 1623939100
transform 1 0 59800 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_631
timestamp 1623939100
transform 1 0 59156 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_637
timestamp 1623939100
transform 1 0 59708 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_639
timestamp 1623939100
transform 1 0 59892 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1623939100
transform 1 0 60812 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output382
timestamp 1623939100
transform 1 0 61548 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_647
timestamp 1623939100
transform 1 0 60628 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_653
timestamp 1623939100
transform 1 0 61180 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_661
timestamp 1623939100
transform 1 0 61916 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1353
timestamp 1623939100
transform 1 0 62468 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1623939100
transform 1 0 63480 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output383
timestamp 1623939100
transform 1 0 64216 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_668
timestamp 1623939100
transform 1 0 62560 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_676
timestamp 1623939100
transform 1 0 63296 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_682
timestamp 1623939100
transform 1 0 63848 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1354
timestamp 1623939100
transform 1 0 65136 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1623939100
transform 1 0 66148 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_690
timestamp 1623939100
transform 1 0 64584 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_697
timestamp 1623939100
transform 1 0 65228 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_705
timestamp 1623939100
transform 1 0 65964 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1355
timestamp 1623939100
transform 1 0 67804 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output384
timestamp 1623939100
transform 1 0 66884 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_711
timestamp 1623939100
transform 1 0 66516 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_719
timestamp 1623939100
transform 1 0 67252 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_726
timestamp 1623939100
transform 1 0 67896 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1623939100
transform 1 0 68724 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output385
timestamp 1623939100
transform 1 0 69460 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_734
timestamp 1623939100
transform 1 0 68632 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_739
timestamp 1623939100
transform 1 0 69092 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_747
timestamp 1623939100
transform 1 0 69828 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1356
timestamp 1623939100
transform 1 0 70472 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1623939100
transform 1 0 71392 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_753
timestamp 1623939100
transform 1 0 70380 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_755
timestamp 1623939100
transform 1 0 70564 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_763
timestamp 1623939100
transform 1 0 71300 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_768
timestamp 1623939100
transform 1 0 71760 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1357
timestamp 1623939100
transform 1 0 73140 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output386
timestamp 1623939100
transform 1 0 72128 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_776
timestamp 1623939100
transform 1 0 72496 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_782
timestamp 1623939100
transform 1 0 73048 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_784
timestamp 1623939100
transform 1 0 73232 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1358
timestamp 1623939100
transform 1 0 75808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1623939100
transform 1 0 73968 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output387
timestamp 1623939100
transform 1 0 74704 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_796
timestamp 1623939100
transform 1 0 74336 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_804
timestamp 1623939100
transform 1 0 75072 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1623939100
transform 1 0 76636 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output388
timestamp 1623939100
transform 1 0 77372 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_813
timestamp 1623939100
transform 1 0 75900 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_825
timestamp 1623939100
transform 1 0 77004 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_833
timestamp 1623939100
transform 1 0 77740 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1359
timestamp 1623939100
transform 1 0 78476 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output389
timestamp 1623939100
transform 1 0 78936 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_842
timestamp 1623939100
transform 1 0 78568 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_850
timestamp 1623939100
transform 1 0 79304 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1360
timestamp 1623939100
transform 1 0 81144 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output391
timestamp 1623939100
transform 1 0 80132 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_858
timestamp 1623939100
transform 1 0 80040 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_863
timestamp 1623939100
transform 1 0 80500 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_869
timestamp 1623939100
transform 1 0 81052 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_871
timestamp 1623939100
transform 1 0 81236 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1623939100
transform 1 0 81880 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output392
timestamp 1623939100
transform 1 0 82800 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_877
timestamp 1623939100
transform 1 0 81788 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_882
timestamp 1623939100
transform 1 0 82248 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_892
timestamp 1623939100
transform 1 0 83168 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1361
timestamp 1623939100
transform 1 0 83812 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output393
timestamp 1623939100
transform -1 0 85744 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output429
timestamp 1623939100
transform 1 0 84272 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_212
timestamp 1623939100
transform -1 0 85376 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_898
timestamp 1623939100
transform 1 0 83720 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_900
timestamp 1623939100
transform 1 0 83904 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_908
timestamp 1623939100
transform 1 0 84640 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1362
timestamp 1623939100
transform 1 0 86480 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output430
timestamp 1623939100
transform 1 0 86940 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_920
timestamp 1623939100
transform 1 0 85744 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_929
timestamp 1623939100
transform 1 0 86572 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_937
timestamp 1623939100
transform 1 0 87308 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1363
timestamp 1623939100
transform 1 0 89148 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output394
timestamp 1623939100
transform -1 0 88412 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_213
timestamp 1623939100
transform -1 0 88044 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_949
timestamp 1623939100
transform 1 0 88412 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_958
timestamp 1623939100
transform 1 0 89240 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output395
timestamp 1623939100
transform -1 0 91080 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output431
timestamp 1623939100
transform -1 0 89976 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_215
timestamp 1623939100
transform -1 0 90712 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_216
timestamp 1623939100
transform -1 0 91264 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_234
timestamp 1623939100
transform -1 0 89608 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_966
timestamp 1623939100
transform 1 0 89976 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1364
timestamp 1623939100
transform 1 0 91816 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output432
timestamp 1623939100
transform -1 0 92644 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_218
timestamp 1623939100
transform -1 0 93288 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_236
timestamp 1623939100
transform -1 0 92276 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_237
timestamp 1623939100
transform -1 0 92828 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_980
timestamp 1623939100
transform 1 0 91264 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_987
timestamp 1623939100
transform 1 0 91908 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_997
timestamp 1623939100
transform 1 0 92828 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1365
timestamp 1623939100
transform 1 0 94484 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output396
timestamp 1623939100
transform -1 0 93656 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output433
timestamp 1623939100
transform 1 0 94944 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_1006
timestamp 1623939100
transform 1 0 93656 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1014
timestamp 1623939100
transform 1 0 94392 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1016
timestamp 1623939100
transform 1 0 94576 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output397
timestamp 1623939100
transform 1 0 95956 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1024
timestamp 1623939100
transform 1 0 95312 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1030
timestamp 1623939100
transform 1 0 95864 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_1035
timestamp 1623939100
transform 1 0 96324 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1623939100
transform -1 0 98808 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1366
timestamp 1623939100
transform 1 0 97152 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output398
timestamp 1623939100
transform 1 0 97796 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_220
timestamp 1623939100
transform 1 0 97612 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_221
timestamp 1623939100
transform 1 0 98164 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1043
timestamp 1623939100
transform 1 0 97060 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1045
timestamp 1623939100
transform 1 0 97244 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1057
timestamp 1623939100
transform 1 0 98348 0 -1 37536
box -38 -48 222 592
<< labels >>
rlabel metal2 s 386 39200 442 40000 6 io_in[0]
port 0 nsew signal input
rlabel metal2 s 26698 39200 26754 40000 6 io_in[10]
port 1 nsew signal input
rlabel metal2 s 29274 39200 29330 40000 6 io_in[11]
port 2 nsew signal input
rlabel metal2 s 31942 39200 31998 40000 6 io_in[12]
port 3 nsew signal input
rlabel metal2 s 34518 39200 34574 40000 6 io_in[13]
port 4 nsew signal input
rlabel metal2 s 37186 39200 37242 40000 6 io_in[14]
port 5 nsew signal input
rlabel metal2 s 39854 39200 39910 40000 6 io_in[15]
port 6 nsew signal input
rlabel metal2 s 42430 39200 42486 40000 6 io_in[16]
port 7 nsew signal input
rlabel metal2 s 45098 39200 45154 40000 6 io_in[17]
port 8 nsew signal input
rlabel metal2 s 47674 39200 47730 40000 6 io_in[18]
port 9 nsew signal input
rlabel metal2 s 50342 39200 50398 40000 6 io_in[19]
port 10 nsew signal input
rlabel metal2 s 2962 39200 3018 40000 6 io_in[1]
port 11 nsew signal input
rlabel metal2 s 53010 39200 53066 40000 6 io_in[20]
port 12 nsew signal input
rlabel metal2 s 55586 39200 55642 40000 6 io_in[21]
port 13 nsew signal input
rlabel metal2 s 58254 39200 58310 40000 6 io_in[22]
port 14 nsew signal input
rlabel metal2 s 60830 39200 60886 40000 6 io_in[23]
port 15 nsew signal input
rlabel metal2 s 63498 39200 63554 40000 6 io_in[24]
port 16 nsew signal input
rlabel metal2 s 66166 39200 66222 40000 6 io_in[25]
port 17 nsew signal input
rlabel metal2 s 68742 39200 68798 40000 6 io_in[26]
port 18 nsew signal input
rlabel metal2 s 71410 39200 71466 40000 6 io_in[27]
port 19 nsew signal input
rlabel metal2 s 73986 39200 74042 40000 6 io_in[28]
port 20 nsew signal input
rlabel metal2 s 76654 39200 76710 40000 6 io_in[29]
port 21 nsew signal input
rlabel metal2 s 5630 39200 5686 40000 6 io_in[2]
port 22 nsew signal input
rlabel metal2 s 79322 39200 79378 40000 6 io_in[30]
port 23 nsew signal input
rlabel metal2 s 81898 39200 81954 40000 6 io_in[31]
port 24 nsew signal input
rlabel metal2 s 84566 39200 84622 40000 6 io_in[32]
port 25 nsew signal input
rlabel metal2 s 87142 39200 87198 40000 6 io_in[33]
port 26 nsew signal input
rlabel metal2 s 89810 39200 89866 40000 6 io_in[34]
port 27 nsew signal input
rlabel metal2 s 92478 39200 92534 40000 6 io_in[35]
port 28 nsew signal input
rlabel metal2 s 95054 39200 95110 40000 6 io_in[36]
port 29 nsew signal input
rlabel metal2 s 97722 39200 97778 40000 6 io_in[37]
port 30 nsew signal input
rlabel metal2 s 8206 39200 8262 40000 6 io_in[3]
port 31 nsew signal input
rlabel metal2 s 10874 39200 10930 40000 6 io_in[4]
port 32 nsew signal input
rlabel metal2 s 13542 39200 13598 40000 6 io_in[5]
port 33 nsew signal input
rlabel metal2 s 16118 39200 16174 40000 6 io_in[6]
port 34 nsew signal input
rlabel metal2 s 18786 39200 18842 40000 6 io_in[7]
port 35 nsew signal input
rlabel metal2 s 21362 39200 21418 40000 6 io_in[8]
port 36 nsew signal input
rlabel metal2 s 24030 39200 24086 40000 6 io_in[9]
port 37 nsew signal input
rlabel metal2 s 1214 39200 1270 40000 6 io_oeb[0]
port 38 nsew signal tristate
rlabel metal2 s 27526 39200 27582 40000 6 io_oeb[10]
port 39 nsew signal tristate
rlabel metal2 s 30194 39200 30250 40000 6 io_oeb[11]
port 40 nsew signal tristate
rlabel metal2 s 32770 39200 32826 40000 6 io_oeb[12]
port 41 nsew signal tristate
rlabel metal2 s 35438 39200 35494 40000 6 io_oeb[13]
port 42 nsew signal tristate
rlabel metal2 s 38106 39200 38162 40000 6 io_oeb[14]
port 43 nsew signal tristate
rlabel metal2 s 40682 39200 40738 40000 6 io_oeb[15]
port 44 nsew signal tristate
rlabel metal2 s 43350 39200 43406 40000 6 io_oeb[16]
port 45 nsew signal tristate
rlabel metal2 s 45926 39200 45982 40000 6 io_oeb[17]
port 46 nsew signal tristate
rlabel metal2 s 48594 39200 48650 40000 6 io_oeb[18]
port 47 nsew signal tristate
rlabel metal2 s 51262 39200 51318 40000 6 io_oeb[19]
port 48 nsew signal tristate
rlabel metal2 s 3882 39200 3938 40000 6 io_oeb[1]
port 49 nsew signal tristate
rlabel metal2 s 53838 39200 53894 40000 6 io_oeb[20]
port 50 nsew signal tristate
rlabel metal2 s 56506 39200 56562 40000 6 io_oeb[21]
port 51 nsew signal tristate
rlabel metal2 s 59082 39200 59138 40000 6 io_oeb[22]
port 52 nsew signal tristate
rlabel metal2 s 61750 39200 61806 40000 6 io_oeb[23]
port 53 nsew signal tristate
rlabel metal2 s 64418 39200 64474 40000 6 io_oeb[24]
port 54 nsew signal tristate
rlabel metal2 s 66994 39200 67050 40000 6 io_oeb[25]
port 55 nsew signal tristate
rlabel metal2 s 69662 39200 69718 40000 6 io_oeb[26]
port 56 nsew signal tristate
rlabel metal2 s 72238 39200 72294 40000 6 io_oeb[27]
port 57 nsew signal tristate
rlabel metal2 s 74906 39200 74962 40000 6 io_oeb[28]
port 58 nsew signal tristate
rlabel metal2 s 77574 39200 77630 40000 6 io_oeb[29]
port 59 nsew signal tristate
rlabel metal2 s 6458 39200 6514 40000 6 io_oeb[2]
port 60 nsew signal tristate
rlabel metal2 s 80150 39200 80206 40000 6 io_oeb[30]
port 61 nsew signal tristate
rlabel metal2 s 82818 39200 82874 40000 6 io_oeb[31]
port 62 nsew signal tristate
rlabel metal2 s 85394 39200 85450 40000 6 io_oeb[32]
port 63 nsew signal tristate
rlabel metal2 s 88062 39200 88118 40000 6 io_oeb[33]
port 64 nsew signal tristate
rlabel metal2 s 90730 39200 90786 40000 6 io_oeb[34]
port 65 nsew signal tristate
rlabel metal2 s 93306 39200 93362 40000 6 io_oeb[35]
port 66 nsew signal tristate
rlabel metal2 s 95974 39200 96030 40000 6 io_oeb[36]
port 67 nsew signal tristate
rlabel metal2 s 98550 39200 98606 40000 6 io_oeb[37]
port 68 nsew signal tristate
rlabel metal2 s 9126 39200 9182 40000 6 io_oeb[3]
port 69 nsew signal tristate
rlabel metal2 s 11702 39200 11758 40000 6 io_oeb[4]
port 70 nsew signal tristate
rlabel metal2 s 14370 39200 14426 40000 6 io_oeb[5]
port 71 nsew signal tristate
rlabel metal2 s 17038 39200 17094 40000 6 io_oeb[6]
port 72 nsew signal tristate
rlabel metal2 s 19614 39200 19670 40000 6 io_oeb[7]
port 73 nsew signal tristate
rlabel metal2 s 22282 39200 22338 40000 6 io_oeb[8]
port 74 nsew signal tristate
rlabel metal2 s 24858 39200 24914 40000 6 io_oeb[9]
port 75 nsew signal tristate
rlabel metal2 s 2134 39200 2190 40000 6 io_out[0]
port 76 nsew signal tristate
rlabel metal2 s 28446 39200 28502 40000 6 io_out[10]
port 77 nsew signal tristate
rlabel metal2 s 31022 39200 31078 40000 6 io_out[11]
port 78 nsew signal tristate
rlabel metal2 s 33690 39200 33746 40000 6 io_out[12]
port 79 nsew signal tristate
rlabel metal2 s 36266 39200 36322 40000 6 io_out[13]
port 80 nsew signal tristate
rlabel metal2 s 38934 39200 38990 40000 6 io_out[14]
port 81 nsew signal tristate
rlabel metal2 s 41602 39200 41658 40000 6 io_out[15]
port 82 nsew signal tristate
rlabel metal2 s 44178 39200 44234 40000 6 io_out[16]
port 83 nsew signal tristate
rlabel metal2 s 46846 39200 46902 40000 6 io_out[17]
port 84 nsew signal tristate
rlabel metal2 s 49422 39200 49478 40000 6 io_out[18]
port 85 nsew signal tristate
rlabel metal2 s 52090 39200 52146 40000 6 io_out[19]
port 86 nsew signal tristate
rlabel metal2 s 4710 39200 4766 40000 6 io_out[1]
port 87 nsew signal tristate
rlabel metal2 s 54758 39200 54814 40000 6 io_out[20]
port 88 nsew signal tristate
rlabel metal2 s 57334 39200 57390 40000 6 io_out[21]
port 89 nsew signal tristate
rlabel metal2 s 60002 39200 60058 40000 6 io_out[22]
port 90 nsew signal tristate
rlabel metal2 s 62578 39200 62634 40000 6 io_out[23]
port 91 nsew signal tristate
rlabel metal2 s 65246 39200 65302 40000 6 io_out[24]
port 92 nsew signal tristate
rlabel metal2 s 67914 39200 67970 40000 6 io_out[25]
port 93 nsew signal tristate
rlabel metal2 s 70490 39200 70546 40000 6 io_out[26]
port 94 nsew signal tristate
rlabel metal2 s 73158 39200 73214 40000 6 io_out[27]
port 95 nsew signal tristate
rlabel metal2 s 75826 39200 75882 40000 6 io_out[28]
port 96 nsew signal tristate
rlabel metal2 s 78402 39200 78458 40000 6 io_out[29]
port 97 nsew signal tristate
rlabel metal2 s 7378 39200 7434 40000 6 io_out[2]
port 98 nsew signal tristate
rlabel metal2 s 81070 39200 81126 40000 6 io_out[30]
port 99 nsew signal tristate
rlabel metal2 s 83646 39200 83702 40000 6 io_out[31]
port 100 nsew signal tristate
rlabel metal2 s 86314 39200 86370 40000 6 io_out[32]
port 101 nsew signal tristate
rlabel metal2 s 88982 39200 89038 40000 6 io_out[33]
port 102 nsew signal tristate
rlabel metal2 s 91558 39200 91614 40000 6 io_out[34]
port 103 nsew signal tristate
rlabel metal2 s 94226 39200 94282 40000 6 io_out[35]
port 104 nsew signal tristate
rlabel metal2 s 96802 39200 96858 40000 6 io_out[36]
port 105 nsew signal tristate
rlabel metal2 s 99470 39200 99526 40000 6 io_out[37]
port 106 nsew signal tristate
rlabel metal2 s 9954 39200 10010 40000 6 io_out[3]
port 107 nsew signal tristate
rlabel metal2 s 12622 39200 12678 40000 6 io_out[4]
port 108 nsew signal tristate
rlabel metal2 s 15290 39200 15346 40000 6 io_out[5]
port 109 nsew signal tristate
rlabel metal2 s 17866 39200 17922 40000 6 io_out[6]
port 110 nsew signal tristate
rlabel metal2 s 20534 39200 20590 40000 6 io_out[7]
port 111 nsew signal tristate
rlabel metal2 s 23110 39200 23166 40000 6 io_out[8]
port 112 nsew signal tristate
rlabel metal2 s 25778 39200 25834 40000 6 io_out[9]
port 113 nsew signal tristate
rlabel metal2 s 99654 0 99710 800 6 irq[0]
port 114 nsew signal tristate
rlabel metal2 s 99838 0 99894 800 6 irq[1]
port 115 nsew signal tristate
rlabel metal3 s 99200 20000 100000 20120 6 irq[2]
port 116 nsew signal tristate
rlabel metal2 s 21638 0 21694 800 6 la_data_in[0]
port 117 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[100]
port 118 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_data_in[101]
port 119 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[102]
port 120 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[103]
port 121 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[104]
port 122 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_data_in[105]
port 123 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[106]
port 124 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[107]
port 125 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[108]
port 126 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[109]
port 127 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[10]
port 128 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[110]
port 129 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_data_in[111]
port 130 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[112]
port 131 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[113]
port 132 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[114]
port 133 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[115]
port 134 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[116]
port 135 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[117]
port 136 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[118]
port 137 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[119]
port 138 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_in[11]
port 139 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[120]
port 140 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[121]
port 141 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[122]
port 142 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[123]
port 143 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[124]
port 144 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[125]
port 145 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[126]
port 146 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[127]
port 147 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in[12]
port 148 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[13]
port 149 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[14]
port 150 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in[15]
port 151 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_data_in[16]
port 152 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[17]
port 153 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[18]
port 154 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_data_in[19]
port 155 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[1]
port 156 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_data_in[20]
port 157 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[21]
port 158 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[22]
port 159 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_data_in[23]
port 160 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[24]
port 161 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[25]
port 162 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_in[26]
port 163 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[27]
port 164 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_data_in[28]
port 165 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[29]
port 166 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_data_in[2]
port 167 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[30]
port 168 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[31]
port 169 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[32]
port 170 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[33]
port 171 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[34]
port 172 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_data_in[35]
port 173 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[36]
port 174 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[37]
port 175 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[38]
port 176 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[39]
port 177 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[3]
port 178 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[40]
port 179 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[41]
port 180 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[42]
port 181 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[43]
port 182 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_data_in[44]
port 183 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[45]
port 184 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[46]
port 185 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[47]
port 186 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_data_in[48]
port 187 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[49]
port 188 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[4]
port 189 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_data_in[50]
port 190 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[51]
port 191 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[52]
port 192 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[53]
port 193 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[54]
port 194 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[55]
port 195 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[56]
port 196 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[57]
port 197 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[58]
port 198 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[59]
port 199 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 la_data_in[5]
port 200 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_data_in[60]
port 201 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[61]
port 202 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[62]
port 203 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[63]
port 204 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[64]
port 205 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[65]
port 206 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[66]
port 207 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_data_in[67]
port 208 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[68]
port 209 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[69]
port 210 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[6]
port 211 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[70]
port 212 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[71]
port 213 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_data_in[72]
port 214 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[73]
port 215 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[74]
port 216 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[75]
port 217 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[76]
port 218 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[77]
port 219 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[78]
port 220 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[79]
port 221 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[7]
port 222 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[80]
port 223 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[81]
port 224 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[82]
port 225 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[83]
port 226 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[84]
port 227 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[85]
port 228 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[86]
port 229 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[87]
port 230 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[88]
port 231 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[89]
port 232 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_data_in[8]
port 233 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[90]
port 234 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[91]
port 235 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[92]
port 236 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[93]
port 237 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[94]
port 238 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[95]
port 239 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[96]
port 240 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[97]
port 241 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[98]
port 242 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[99]
port 243 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[9]
port 244 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_out[0]
port 245 nsew signal tristate
rlabel metal2 s 82818 0 82874 800 6 la_data_out[100]
port 246 nsew signal tristate
rlabel metal2 s 83370 0 83426 800 6 la_data_out[101]
port 247 nsew signal tristate
rlabel metal2 s 84014 0 84070 800 6 la_data_out[102]
port 248 nsew signal tristate
rlabel metal2 s 84658 0 84714 800 6 la_data_out[103]
port 249 nsew signal tristate
rlabel metal2 s 85210 0 85266 800 6 la_data_out[104]
port 250 nsew signal tristate
rlabel metal2 s 85854 0 85910 800 6 la_data_out[105]
port 251 nsew signal tristate
rlabel metal2 s 86406 0 86462 800 6 la_data_out[106]
port 252 nsew signal tristate
rlabel metal2 s 87050 0 87106 800 6 la_data_out[107]
port 253 nsew signal tristate
rlabel metal2 s 87694 0 87750 800 6 la_data_out[108]
port 254 nsew signal tristate
rlabel metal2 s 88246 0 88302 800 6 la_data_out[109]
port 255 nsew signal tristate
rlabel metal2 s 27894 0 27950 800 6 la_data_out[10]
port 256 nsew signal tristate
rlabel metal2 s 88890 0 88946 800 6 la_data_out[110]
port 257 nsew signal tristate
rlabel metal2 s 89534 0 89590 800 6 la_data_out[111]
port 258 nsew signal tristate
rlabel metal2 s 90086 0 90142 800 6 la_data_out[112]
port 259 nsew signal tristate
rlabel metal2 s 90730 0 90786 800 6 la_data_out[113]
port 260 nsew signal tristate
rlabel metal2 s 91282 0 91338 800 6 la_data_out[114]
port 261 nsew signal tristate
rlabel metal2 s 91926 0 91982 800 6 la_data_out[115]
port 262 nsew signal tristate
rlabel metal2 s 92570 0 92626 800 6 la_data_out[116]
port 263 nsew signal tristate
rlabel metal2 s 93122 0 93178 800 6 la_data_out[117]
port 264 nsew signal tristate
rlabel metal2 s 93766 0 93822 800 6 la_data_out[118]
port 265 nsew signal tristate
rlabel metal2 s 94410 0 94466 800 6 la_data_out[119]
port 266 nsew signal tristate
rlabel metal2 s 28538 0 28594 800 6 la_data_out[11]
port 267 nsew signal tristate
rlabel metal2 s 94962 0 95018 800 6 la_data_out[120]
port 268 nsew signal tristate
rlabel metal2 s 95606 0 95662 800 6 la_data_out[121]
port 269 nsew signal tristate
rlabel metal2 s 96250 0 96306 800 6 la_data_out[122]
port 270 nsew signal tristate
rlabel metal2 s 96802 0 96858 800 6 la_data_out[123]
port 271 nsew signal tristate
rlabel metal2 s 97446 0 97502 800 6 la_data_out[124]
port 272 nsew signal tristate
rlabel metal2 s 97998 0 98054 800 6 la_data_out[125]
port 273 nsew signal tristate
rlabel metal2 s 98642 0 98698 800 6 la_data_out[126]
port 274 nsew signal tristate
rlabel metal2 s 99286 0 99342 800 6 la_data_out[127]
port 275 nsew signal tristate
rlabel metal2 s 29090 0 29146 800 6 la_data_out[12]
port 276 nsew signal tristate
rlabel metal2 s 29734 0 29790 800 6 la_data_out[13]
port 277 nsew signal tristate
rlabel metal2 s 30378 0 30434 800 6 la_data_out[14]
port 278 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 la_data_out[15]
port 279 nsew signal tristate
rlabel metal2 s 31574 0 31630 800 6 la_data_out[16]
port 280 nsew signal tristate
rlabel metal2 s 32218 0 32274 800 6 la_data_out[17]
port 281 nsew signal tristate
rlabel metal2 s 32770 0 32826 800 6 la_data_out[18]
port 282 nsew signal tristate
rlabel metal2 s 33414 0 33470 800 6 la_data_out[19]
port 283 nsew signal tristate
rlabel metal2 s 22466 0 22522 800 6 la_data_out[1]
port 284 nsew signal tristate
rlabel metal2 s 33966 0 34022 800 6 la_data_out[20]
port 285 nsew signal tristate
rlabel metal2 s 34610 0 34666 800 6 la_data_out[21]
port 286 nsew signal tristate
rlabel metal2 s 35254 0 35310 800 6 la_data_out[22]
port 287 nsew signal tristate
rlabel metal2 s 35806 0 35862 800 6 la_data_out[23]
port 288 nsew signal tristate
rlabel metal2 s 36450 0 36506 800 6 la_data_out[24]
port 289 nsew signal tristate
rlabel metal2 s 37094 0 37150 800 6 la_data_out[25]
port 290 nsew signal tristate
rlabel metal2 s 37646 0 37702 800 6 la_data_out[26]
port 291 nsew signal tristate
rlabel metal2 s 38290 0 38346 800 6 la_data_out[27]
port 292 nsew signal tristate
rlabel metal2 s 38842 0 38898 800 6 la_data_out[28]
port 293 nsew signal tristate
rlabel metal2 s 39486 0 39542 800 6 la_data_out[29]
port 294 nsew signal tristate
rlabel metal2 s 23018 0 23074 800 6 la_data_out[2]
port 295 nsew signal tristate
rlabel metal2 s 40130 0 40186 800 6 la_data_out[30]
port 296 nsew signal tristate
rlabel metal2 s 40682 0 40738 800 6 la_data_out[31]
port 297 nsew signal tristate
rlabel metal2 s 41326 0 41382 800 6 la_data_out[32]
port 298 nsew signal tristate
rlabel metal2 s 41970 0 42026 800 6 la_data_out[33]
port 299 nsew signal tristate
rlabel metal2 s 42522 0 42578 800 6 la_data_out[34]
port 300 nsew signal tristate
rlabel metal2 s 43166 0 43222 800 6 la_data_out[35]
port 301 nsew signal tristate
rlabel metal2 s 43810 0 43866 800 6 la_data_out[36]
port 302 nsew signal tristate
rlabel metal2 s 44362 0 44418 800 6 la_data_out[37]
port 303 nsew signal tristate
rlabel metal2 s 45006 0 45062 800 6 la_data_out[38]
port 304 nsew signal tristate
rlabel metal2 s 45558 0 45614 800 6 la_data_out[39]
port 305 nsew signal tristate
rlabel metal2 s 23662 0 23718 800 6 la_data_out[3]
port 306 nsew signal tristate
rlabel metal2 s 46202 0 46258 800 6 la_data_out[40]
port 307 nsew signal tristate
rlabel metal2 s 46846 0 46902 800 6 la_data_out[41]
port 308 nsew signal tristate
rlabel metal2 s 47398 0 47454 800 6 la_data_out[42]
port 309 nsew signal tristate
rlabel metal2 s 48042 0 48098 800 6 la_data_out[43]
port 310 nsew signal tristate
rlabel metal2 s 48686 0 48742 800 6 la_data_out[44]
port 311 nsew signal tristate
rlabel metal2 s 49238 0 49294 800 6 la_data_out[45]
port 312 nsew signal tristate
rlabel metal2 s 49882 0 49938 800 6 la_data_out[46]
port 313 nsew signal tristate
rlabel metal2 s 50434 0 50490 800 6 la_data_out[47]
port 314 nsew signal tristate
rlabel metal2 s 51078 0 51134 800 6 la_data_out[48]
port 315 nsew signal tristate
rlabel metal2 s 51722 0 51778 800 6 la_data_out[49]
port 316 nsew signal tristate
rlabel metal2 s 24214 0 24270 800 6 la_data_out[4]
port 317 nsew signal tristate
rlabel metal2 s 52274 0 52330 800 6 la_data_out[50]
port 318 nsew signal tristate
rlabel metal2 s 52918 0 52974 800 6 la_data_out[51]
port 319 nsew signal tristate
rlabel metal2 s 53562 0 53618 800 6 la_data_out[52]
port 320 nsew signal tristate
rlabel metal2 s 54114 0 54170 800 6 la_data_out[53]
port 321 nsew signal tristate
rlabel metal2 s 54758 0 54814 800 6 la_data_out[54]
port 322 nsew signal tristate
rlabel metal2 s 55310 0 55366 800 6 la_data_out[55]
port 323 nsew signal tristate
rlabel metal2 s 55954 0 56010 800 6 la_data_out[56]
port 324 nsew signal tristate
rlabel metal2 s 56598 0 56654 800 6 la_data_out[57]
port 325 nsew signal tristate
rlabel metal2 s 57150 0 57206 800 6 la_data_out[58]
port 326 nsew signal tristate
rlabel metal2 s 57794 0 57850 800 6 la_data_out[59]
port 327 nsew signal tristate
rlabel metal2 s 24858 0 24914 800 6 la_data_out[5]
port 328 nsew signal tristate
rlabel metal2 s 58438 0 58494 800 6 la_data_out[60]
port 329 nsew signal tristate
rlabel metal2 s 58990 0 59046 800 6 la_data_out[61]
port 330 nsew signal tristate
rlabel metal2 s 59634 0 59690 800 6 la_data_out[62]
port 331 nsew signal tristate
rlabel metal2 s 60186 0 60242 800 6 la_data_out[63]
port 332 nsew signal tristate
rlabel metal2 s 60830 0 60886 800 6 la_data_out[64]
port 333 nsew signal tristate
rlabel metal2 s 61474 0 61530 800 6 la_data_out[65]
port 334 nsew signal tristate
rlabel metal2 s 62026 0 62082 800 6 la_data_out[66]
port 335 nsew signal tristate
rlabel metal2 s 62670 0 62726 800 6 la_data_out[67]
port 336 nsew signal tristate
rlabel metal2 s 63314 0 63370 800 6 la_data_out[68]
port 337 nsew signal tristate
rlabel metal2 s 63866 0 63922 800 6 la_data_out[69]
port 338 nsew signal tristate
rlabel metal2 s 25502 0 25558 800 6 la_data_out[6]
port 339 nsew signal tristate
rlabel metal2 s 64510 0 64566 800 6 la_data_out[70]
port 340 nsew signal tristate
rlabel metal2 s 65062 0 65118 800 6 la_data_out[71]
port 341 nsew signal tristate
rlabel metal2 s 65706 0 65762 800 6 la_data_out[72]
port 342 nsew signal tristate
rlabel metal2 s 66350 0 66406 800 6 la_data_out[73]
port 343 nsew signal tristate
rlabel metal2 s 66902 0 66958 800 6 la_data_out[74]
port 344 nsew signal tristate
rlabel metal2 s 67546 0 67602 800 6 la_data_out[75]
port 345 nsew signal tristate
rlabel metal2 s 68190 0 68246 800 6 la_data_out[76]
port 346 nsew signal tristate
rlabel metal2 s 68742 0 68798 800 6 la_data_out[77]
port 347 nsew signal tristate
rlabel metal2 s 69386 0 69442 800 6 la_data_out[78]
port 348 nsew signal tristate
rlabel metal2 s 70030 0 70086 800 6 la_data_out[79]
port 349 nsew signal tristate
rlabel metal2 s 26054 0 26110 800 6 la_data_out[7]
port 350 nsew signal tristate
rlabel metal2 s 70582 0 70638 800 6 la_data_out[80]
port 351 nsew signal tristate
rlabel metal2 s 71226 0 71282 800 6 la_data_out[81]
port 352 nsew signal tristate
rlabel metal2 s 71778 0 71834 800 6 la_data_out[82]
port 353 nsew signal tristate
rlabel metal2 s 72422 0 72478 800 6 la_data_out[83]
port 354 nsew signal tristate
rlabel metal2 s 73066 0 73122 800 6 la_data_out[84]
port 355 nsew signal tristate
rlabel metal2 s 73618 0 73674 800 6 la_data_out[85]
port 356 nsew signal tristate
rlabel metal2 s 74262 0 74318 800 6 la_data_out[86]
port 357 nsew signal tristate
rlabel metal2 s 74906 0 74962 800 6 la_data_out[87]
port 358 nsew signal tristate
rlabel metal2 s 75458 0 75514 800 6 la_data_out[88]
port 359 nsew signal tristate
rlabel metal2 s 76102 0 76158 800 6 la_data_out[89]
port 360 nsew signal tristate
rlabel metal2 s 26698 0 26754 800 6 la_data_out[8]
port 361 nsew signal tristate
rlabel metal2 s 76654 0 76710 800 6 la_data_out[90]
port 362 nsew signal tristate
rlabel metal2 s 77298 0 77354 800 6 la_data_out[91]
port 363 nsew signal tristate
rlabel metal2 s 77942 0 77998 800 6 la_data_out[92]
port 364 nsew signal tristate
rlabel metal2 s 78494 0 78550 800 6 la_data_out[93]
port 365 nsew signal tristate
rlabel metal2 s 79138 0 79194 800 6 la_data_out[94]
port 366 nsew signal tristate
rlabel metal2 s 79782 0 79838 800 6 la_data_out[95]
port 367 nsew signal tristate
rlabel metal2 s 80334 0 80390 800 6 la_data_out[96]
port 368 nsew signal tristate
rlabel metal2 s 80978 0 81034 800 6 la_data_out[97]
port 369 nsew signal tristate
rlabel metal2 s 81530 0 81586 800 6 la_data_out[98]
port 370 nsew signal tristate
rlabel metal2 s 82174 0 82230 800 6 la_data_out[99]
port 371 nsew signal tristate
rlabel metal2 s 27342 0 27398 800 6 la_data_out[9]
port 372 nsew signal tristate
rlabel metal2 s 22006 0 22062 800 6 la_oenb[0]
port 373 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[100]
port 374 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[101]
port 375 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[102]
port 376 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_oenb[103]
port 377 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[104]
port 378 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[105]
port 379 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[106]
port 380 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[107]
port 381 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[108]
port 382 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[109]
port 383 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[10]
port 384 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oenb[110]
port 385 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[111]
port 386 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[112]
port 387 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[113]
port 388 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[114]
port 389 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[115]
port 390 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[116]
port 391 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[117]
port 392 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[118]
port 393 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[119]
port 394 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[11]
port 395 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[120]
port 396 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[121]
port 397 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[122]
port 398 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[123]
port 399 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[124]
port 400 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_oenb[125]
port 401 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[126]
port 402 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[127]
port 403 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[12]
port 404 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[13]
port 405 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_oenb[14]
port 406 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_oenb[15]
port 407 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_oenb[16]
port 408 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_oenb[17]
port 409 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[18]
port 410 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_oenb[19]
port 411 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_oenb[1]
port 412 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_oenb[20]
port 413 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_oenb[21]
port 414 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_oenb[22]
port 415 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[23]
port 416 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_oenb[24]
port 417 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_oenb[25]
port 418 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[26]
port 419 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_oenb[27]
port 420 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[28]
port 421 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_oenb[29]
port 422 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 la_oenb[2]
port 423 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_oenb[30]
port 424 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[31]
port 425 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_oenb[32]
port 426 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_oenb[33]
port 427 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[34]
port 428 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[35]
port 429 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[36]
port 430 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[37]
port 431 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[38]
port 432 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[39]
port 433 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_oenb[3]
port 434 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[40]
port 435 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[41]
port 436 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[42]
port 437 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[43]
port 438 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[44]
port 439 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_oenb[45]
port 440 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_oenb[46]
port 441 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[47]
port 442 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[48]
port 443 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[49]
port 444 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_oenb[4]
port 445 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[50]
port 446 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[51]
port 447 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[52]
port 448 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_oenb[53]
port 449 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[54]
port 450 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[55]
port 451 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[56]
port 452 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[57]
port 453 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[58]
port 454 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_oenb[59]
port 455 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_oenb[5]
port 456 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[60]
port 457 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[61]
port 458 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[62]
port 459 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[63]
port 460 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[64]
port 461 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[65]
port 462 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oenb[66]
port 463 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[67]
port 464 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[68]
port 465 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_oenb[69]
port 466 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_oenb[6]
port 467 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[70]
port 468 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oenb[71]
port 469 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[72]
port 470 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[73]
port 471 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[74]
port 472 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[75]
port 473 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[76]
port 474 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[77]
port 475 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oenb[78]
port 476 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[79]
port 477 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[7]
port 478 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[80]
port 479 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[81]
port 480 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[82]
port 481 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_oenb[83]
port 482 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oenb[84]
port 483 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[85]
port 484 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_oenb[86]
port 485 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[87]
port 486 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[88]
port 487 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[89]
port 488 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_oenb[8]
port 489 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[90]
port 490 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_oenb[91]
port 491 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[92]
port 492 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[93]
port 493 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[94]
port 494 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[95]
port 495 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[96]
port 496 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_oenb[97]
port 497 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[98]
port 498 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[99]
port 499 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[9]
port 500 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 user_clock2
port 501 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 504 nsew signal tristate
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 570 nsew signal tristate
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[10]
port 571 nsew signal tristate
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[11]
port 572 nsew signal tristate
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[12]
port 573 nsew signal tristate
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[13]
port 574 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[14]
port 575 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[15]
port 576 nsew signal tristate
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[16]
port 577 nsew signal tristate
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[17]
port 578 nsew signal tristate
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[18]
port 579 nsew signal tristate
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[19]
port 580 nsew signal tristate
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[1]
port 581 nsew signal tristate
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[20]
port 582 nsew signal tristate
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[21]
port 583 nsew signal tristate
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[22]
port 584 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[23]
port 585 nsew signal tristate
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[24]
port 586 nsew signal tristate
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[25]
port 587 nsew signal tristate
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[26]
port 588 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[27]
port 589 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[28]
port 590 nsew signal tristate
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[29]
port 591 nsew signal tristate
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[2]
port 592 nsew signal tristate
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[30]
port 593 nsew signal tristate
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[31]
port 594 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[3]
port 595 nsew signal tristate
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[4]
port 596 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[5]
port 597 nsew signal tristate
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[6]
port 598 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[7]
port 599 nsew signal tristate
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[8]
port 600 nsew signal tristate
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[9]
port 601 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 96368 2128 96688 37584 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 81008 2128 81328 37584 6 vssd1
port 612 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 613 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 97028 2176 97348 37536 6 vccd2
port 615 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 37536 6 vccd2
port 616 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 37536 6 vccd2
port 617 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 37536 6 vccd2
port 618 nsew power bidirectional
rlabel metal4 s 81668 2176 81988 37536 6 vssd2
port 619 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 37536 6 vssd2
port 620 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 37536 6 vssd2
port 621 nsew ground bidirectional
rlabel metal4 s 97688 2176 98008 37536 6 vdda1
port 622 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 37536 6 vdda1
port 623 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 37536 6 vdda1
port 624 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 37536 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 82328 2176 82648 37536 6 vssa1
port 626 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 37536 6 vssa1
port 627 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 37536 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 67628 2176 67948 37536 6 vdda2
port 629 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 37536 6 vdda2
port 630 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 37536 6 vdda2
port 631 nsew power bidirectional
rlabel metal4 s 82988 2176 83308 37536 6 vssa2
port 632 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 37536 6 vssa2
port 633 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 37536 6 vssa2
port 634 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
