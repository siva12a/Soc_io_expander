magic
tech sky130A
magscale 1 2
timestamp 1623239208
<< obsli1 >>
rect 1409 2261 98135 97291
<< obsm1 >>
rect 106 1368 99898 97640
<< metal2 >>
rect 386 99200 442 100000
rect 1214 99200 1270 100000
rect 2042 99200 2098 100000
rect 2962 99200 3018 100000
rect 3790 99200 3846 100000
rect 4710 99200 4766 100000
rect 5538 99200 5594 100000
rect 6458 99200 6514 100000
rect 7286 99200 7342 100000
rect 8206 99200 8262 100000
rect 9034 99200 9090 100000
rect 9862 99200 9918 100000
rect 10782 99200 10838 100000
rect 11610 99200 11666 100000
rect 12530 99200 12586 100000
rect 13358 99200 13414 100000
rect 14278 99200 14334 100000
rect 15106 99200 15162 100000
rect 16026 99200 16082 100000
rect 16854 99200 16910 100000
rect 17774 99200 17830 100000
rect 18602 99200 18658 100000
rect 19430 99200 19486 100000
rect 20350 99200 20406 100000
rect 21178 99200 21234 100000
rect 22098 99200 22154 100000
rect 22926 99200 22982 100000
rect 23846 99200 23902 100000
rect 24674 99200 24730 100000
rect 25594 99200 25650 100000
rect 26422 99200 26478 100000
rect 27342 99200 27398 100000
rect 28170 99200 28226 100000
rect 28998 99200 29054 100000
rect 29918 99200 29974 100000
rect 30746 99200 30802 100000
rect 31666 99200 31722 100000
rect 32494 99200 32550 100000
rect 33414 99200 33470 100000
rect 34242 99200 34298 100000
rect 35162 99200 35218 100000
rect 35990 99200 36046 100000
rect 36818 99200 36874 100000
rect 37738 99200 37794 100000
rect 38566 99200 38622 100000
rect 39486 99200 39542 100000
rect 40314 99200 40370 100000
rect 41234 99200 41290 100000
rect 42062 99200 42118 100000
rect 42982 99200 43038 100000
rect 43810 99200 43866 100000
rect 44730 99200 44786 100000
rect 45558 99200 45614 100000
rect 46386 99200 46442 100000
rect 47306 99200 47362 100000
rect 48134 99200 48190 100000
rect 49054 99200 49110 100000
rect 49882 99200 49938 100000
rect 50802 99200 50858 100000
rect 51630 99200 51686 100000
rect 52550 99200 52606 100000
rect 53378 99200 53434 100000
rect 54298 99200 54354 100000
rect 55126 99200 55182 100000
rect 55954 99200 56010 100000
rect 56874 99200 56930 100000
rect 57702 99200 57758 100000
rect 58622 99200 58678 100000
rect 59450 99200 59506 100000
rect 60370 99200 60426 100000
rect 61198 99200 61254 100000
rect 62118 99200 62174 100000
rect 62946 99200 63002 100000
rect 63866 99200 63922 100000
rect 64694 99200 64750 100000
rect 65522 99200 65578 100000
rect 66442 99200 66498 100000
rect 67270 99200 67326 100000
rect 68190 99200 68246 100000
rect 69018 99200 69074 100000
rect 69938 99200 69994 100000
rect 70766 99200 70822 100000
rect 71686 99200 71742 100000
rect 72514 99200 72570 100000
rect 73342 99200 73398 100000
rect 74262 99200 74318 100000
rect 75090 99200 75146 100000
rect 76010 99200 76066 100000
rect 76838 99200 76894 100000
rect 77758 99200 77814 100000
rect 78586 99200 78642 100000
rect 79506 99200 79562 100000
rect 80334 99200 80390 100000
rect 81254 99200 81310 100000
rect 82082 99200 82138 100000
rect 82910 99200 82966 100000
rect 83830 99200 83886 100000
rect 84658 99200 84714 100000
rect 85578 99200 85634 100000
rect 86406 99200 86462 100000
rect 87326 99200 87382 100000
rect 88154 99200 88210 100000
rect 89074 99200 89130 100000
rect 89902 99200 89958 100000
rect 90822 99200 90878 100000
rect 91650 99200 91706 100000
rect 92478 99200 92534 100000
rect 93398 99200 93454 100000
rect 94226 99200 94282 100000
rect 95146 99200 95202 100000
rect 95974 99200 96030 100000
rect 96894 99200 96950 100000
rect 97722 99200 97778 100000
rect 98642 99200 98698 100000
rect 99470 99200 99526 100000
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9678 0 9734 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10690 0 10746 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13726 0 13782 800
rect 13910 0 13966 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16762 0 16818 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18418 0 18474 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20442 0 20498 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22282 0 22338 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29826 0 29882 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30378 0 30434 800
rect 30654 0 30710 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31666 0 31722 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32218 0 32274 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 33046 0 33102 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34058 0 34114 800
rect 34242 0 34298 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39210 0 39266 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40590 0 40646 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 43074 0 43130 800
rect 43258 0 43314 800
rect 43442 0 43498 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44914 0 44970 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46938 0 46994 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53194 0 53250 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55218 0 55274 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56874 0 56930 800
rect 57058 0 57114 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58714 0 58770 800
rect 58898 0 58954 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60554 0 60610 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61566 0 61622 800
rect 61750 0 61806 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62394 0 62450 800
rect 62578 0 62634 800
rect 62762 0 62818 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 64050 0 64106 800
rect 64234 0 64290 800
rect 64418 0 64474 800
rect 64602 0 64658 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65246 0 65302 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65890 0 65946 800
rect 66074 0 66130 800
rect 66258 0 66314 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67086 0 67142 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67914 0 67970 800
rect 68098 0 68154 800
rect 68282 0 68338 800
rect 68466 0 68522 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69478 0 69534 800
rect 69754 0 69810 800
rect 69938 0 69994 800
rect 70122 0 70178 800
rect 70306 0 70362 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 71962 0 72018 800
rect 72146 0 72202 800
rect 72330 0 72386 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73618 0 73674 800
rect 73802 0 73858 800
rect 73986 0 74042 800
rect 74170 0 74226 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75826 0 75882 800
rect 76010 0 76066 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77022 0 77078 800
rect 77298 0 77354 800
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77850 0 77906 800
rect 78034 0 78090 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79046 0 79102 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79690 0 79746 800
rect 79874 0 79930 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80702 0 80758 800
rect 80886 0 80942 800
rect 81162 0 81218 800
rect 81346 0 81402 800
rect 81530 0 81586 800
rect 81714 0 81770 800
rect 81898 0 81954 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 83002 0 83058 800
rect 83186 0 83242 800
rect 83370 0 83426 800
rect 83554 0 83610 800
rect 83738 0 83794 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84566 0 84622 800
rect 84750 0 84806 800
rect 85026 0 85082 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85578 0 85634 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86590 0 86646 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87234 0 87290 800
rect 87418 0 87474 800
rect 87602 0 87658 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88430 0 88486 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89258 0 89314 800
rect 89442 0 89498 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90454 0 90510 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92294 0 92350 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 92938 0 92994 800
rect 93122 0 93178 800
rect 93306 0 93362 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95146 0 95202 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96158 0 96214 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< obsm2 >>
rect 112 99144 330 99200
rect 498 99144 1158 99200
rect 1326 99144 1986 99200
rect 2154 99144 2906 99200
rect 3074 99144 3734 99200
rect 3902 99144 4654 99200
rect 4822 99144 5482 99200
rect 5650 99144 6402 99200
rect 6570 99144 7230 99200
rect 7398 99144 8150 99200
rect 8318 99144 8978 99200
rect 9146 99144 9806 99200
rect 9974 99144 10726 99200
rect 10894 99144 11554 99200
rect 11722 99144 12474 99200
rect 12642 99144 13302 99200
rect 13470 99144 14222 99200
rect 14390 99144 15050 99200
rect 15218 99144 15970 99200
rect 16138 99144 16798 99200
rect 16966 99144 17718 99200
rect 17886 99144 18546 99200
rect 18714 99144 19374 99200
rect 19542 99144 20294 99200
rect 20462 99144 21122 99200
rect 21290 99144 22042 99200
rect 22210 99144 22870 99200
rect 23038 99144 23790 99200
rect 23958 99144 24618 99200
rect 24786 99144 25538 99200
rect 25706 99144 26366 99200
rect 26534 99144 27286 99200
rect 27454 99144 28114 99200
rect 28282 99144 28942 99200
rect 29110 99144 29862 99200
rect 30030 99144 30690 99200
rect 30858 99144 31610 99200
rect 31778 99144 32438 99200
rect 32606 99144 33358 99200
rect 33526 99144 34186 99200
rect 34354 99144 35106 99200
rect 35274 99144 35934 99200
rect 36102 99144 36762 99200
rect 36930 99144 37682 99200
rect 37850 99144 38510 99200
rect 38678 99144 39430 99200
rect 39598 99144 40258 99200
rect 40426 99144 41178 99200
rect 41346 99144 42006 99200
rect 42174 99144 42926 99200
rect 43094 99144 43754 99200
rect 43922 99144 44674 99200
rect 44842 99144 45502 99200
rect 45670 99144 46330 99200
rect 46498 99144 47250 99200
rect 47418 99144 48078 99200
rect 48246 99144 48998 99200
rect 49166 99144 49826 99200
rect 49994 99144 50746 99200
rect 50914 99144 51574 99200
rect 51742 99144 52494 99200
rect 52662 99144 53322 99200
rect 53490 99144 54242 99200
rect 54410 99144 55070 99200
rect 55238 99144 55898 99200
rect 56066 99144 56818 99200
rect 56986 99144 57646 99200
rect 57814 99144 58566 99200
rect 58734 99144 59394 99200
rect 59562 99144 60314 99200
rect 60482 99144 61142 99200
rect 61310 99144 62062 99200
rect 62230 99144 62890 99200
rect 63058 99144 63810 99200
rect 63978 99144 64638 99200
rect 64806 99144 65466 99200
rect 65634 99144 66386 99200
rect 66554 99144 67214 99200
rect 67382 99144 68134 99200
rect 68302 99144 68962 99200
rect 69130 99144 69882 99200
rect 70050 99144 70710 99200
rect 70878 99144 71630 99200
rect 71798 99144 72458 99200
rect 72626 99144 73286 99200
rect 73454 99144 74206 99200
rect 74374 99144 75034 99200
rect 75202 99144 75954 99200
rect 76122 99144 76782 99200
rect 76950 99144 77702 99200
rect 77870 99144 78530 99200
rect 78698 99144 79450 99200
rect 79618 99144 80278 99200
rect 80446 99144 81198 99200
rect 81366 99144 82026 99200
rect 82194 99144 82854 99200
rect 83022 99144 83774 99200
rect 83942 99144 84602 99200
rect 84770 99144 85522 99200
rect 85690 99144 86350 99200
rect 86518 99144 87270 99200
rect 87438 99144 88098 99200
rect 88266 99144 89018 99200
rect 89186 99144 89846 99200
rect 90014 99144 90766 99200
rect 90934 99144 91594 99200
rect 91762 99144 92422 99200
rect 92590 99144 93342 99200
rect 93510 99144 94170 99200
rect 94338 99144 95090 99200
rect 95258 99144 95918 99200
rect 96086 99144 96838 99200
rect 97006 99144 97666 99200
rect 97834 99144 98586 99200
rect 98754 99144 99414 99200
rect 99582 99144 99892 99200
rect 112 856 99892 99144
rect 222 800 238 856
rect 406 800 422 856
rect 590 800 606 856
rect 774 800 790 856
rect 958 800 1066 856
rect 1234 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1618 856
rect 1786 800 1802 856
rect 1970 800 2078 856
rect 2246 800 2262 856
rect 2430 800 2446 856
rect 2614 800 2630 856
rect 2798 800 2814 856
rect 2982 800 3090 856
rect 3258 800 3274 856
rect 3442 800 3458 856
rect 3626 800 3642 856
rect 3810 800 3918 856
rect 4086 800 4102 856
rect 4270 800 4286 856
rect 4454 800 4470 856
rect 4638 800 4654 856
rect 4822 800 4930 856
rect 5098 800 5114 856
rect 5282 800 5298 856
rect 5466 800 5482 856
rect 5650 800 5666 856
rect 5834 800 5942 856
rect 6110 800 6126 856
rect 6294 800 6310 856
rect 6478 800 6494 856
rect 6662 800 6770 856
rect 6938 800 6954 856
rect 7122 800 7138 856
rect 7306 800 7322 856
rect 7490 800 7506 856
rect 7674 800 7782 856
rect 7950 800 7966 856
rect 8134 800 8150 856
rect 8318 800 8334 856
rect 8502 800 8518 856
rect 8686 800 8794 856
rect 8962 800 8978 856
rect 9146 800 9162 856
rect 9330 800 9346 856
rect 9514 800 9622 856
rect 9790 800 9806 856
rect 9974 800 9990 856
rect 10158 800 10174 856
rect 10342 800 10358 856
rect 10526 800 10634 856
rect 10802 800 10818 856
rect 10986 800 11002 856
rect 11170 800 11186 856
rect 11354 800 11370 856
rect 11538 800 11646 856
rect 11814 800 11830 856
rect 11998 800 12014 856
rect 12182 800 12198 856
rect 12366 800 12474 856
rect 12642 800 12658 856
rect 12826 800 12842 856
rect 13010 800 13026 856
rect 13194 800 13210 856
rect 13378 800 13486 856
rect 13654 800 13670 856
rect 13838 800 13854 856
rect 14022 800 14038 856
rect 14206 800 14222 856
rect 14390 800 14498 856
rect 14666 800 14682 856
rect 14850 800 14866 856
rect 15034 800 15050 856
rect 15218 800 15326 856
rect 15494 800 15510 856
rect 15678 800 15694 856
rect 15862 800 15878 856
rect 16046 800 16062 856
rect 16230 800 16338 856
rect 16506 800 16522 856
rect 16690 800 16706 856
rect 16874 800 16890 856
rect 17058 800 17074 856
rect 17242 800 17350 856
rect 17518 800 17534 856
rect 17702 800 17718 856
rect 17886 800 17902 856
rect 18070 800 18178 856
rect 18346 800 18362 856
rect 18530 800 18546 856
rect 18714 800 18730 856
rect 18898 800 18914 856
rect 19082 800 19190 856
rect 19358 800 19374 856
rect 19542 800 19558 856
rect 19726 800 19742 856
rect 19910 800 19926 856
rect 20094 800 20202 856
rect 20370 800 20386 856
rect 20554 800 20570 856
rect 20738 800 20754 856
rect 20922 800 21030 856
rect 21198 800 21214 856
rect 21382 800 21398 856
rect 21566 800 21582 856
rect 21750 800 21766 856
rect 21934 800 22042 856
rect 22210 800 22226 856
rect 22394 800 22410 856
rect 22578 800 22594 856
rect 22762 800 22778 856
rect 22946 800 23054 856
rect 23222 800 23238 856
rect 23406 800 23422 856
rect 23590 800 23606 856
rect 23774 800 23882 856
rect 24050 800 24066 856
rect 24234 800 24250 856
rect 24418 800 24434 856
rect 24602 800 24618 856
rect 24786 800 24894 856
rect 25062 800 25078 856
rect 25246 800 25262 856
rect 25430 800 25446 856
rect 25614 800 25630 856
rect 25798 800 25906 856
rect 26074 800 26090 856
rect 26258 800 26274 856
rect 26442 800 26458 856
rect 26626 800 26734 856
rect 26902 800 26918 856
rect 27086 800 27102 856
rect 27270 800 27286 856
rect 27454 800 27470 856
rect 27638 800 27746 856
rect 27914 800 27930 856
rect 28098 800 28114 856
rect 28282 800 28298 856
rect 28466 800 28482 856
rect 28650 800 28758 856
rect 28926 800 28942 856
rect 29110 800 29126 856
rect 29294 800 29310 856
rect 29478 800 29586 856
rect 29754 800 29770 856
rect 29938 800 29954 856
rect 30122 800 30138 856
rect 30306 800 30322 856
rect 30490 800 30598 856
rect 30766 800 30782 856
rect 30950 800 30966 856
rect 31134 800 31150 856
rect 31318 800 31334 856
rect 31502 800 31610 856
rect 31778 800 31794 856
rect 31962 800 31978 856
rect 32146 800 32162 856
rect 32330 800 32438 856
rect 32606 800 32622 856
rect 32790 800 32806 856
rect 32974 800 32990 856
rect 33158 800 33174 856
rect 33342 800 33450 856
rect 33618 800 33634 856
rect 33802 800 33818 856
rect 33986 800 34002 856
rect 34170 800 34186 856
rect 34354 800 34462 856
rect 34630 800 34646 856
rect 34814 800 34830 856
rect 34998 800 35014 856
rect 35182 800 35198 856
rect 35366 800 35474 856
rect 35642 800 35658 856
rect 35826 800 35842 856
rect 36010 800 36026 856
rect 36194 800 36302 856
rect 36470 800 36486 856
rect 36654 800 36670 856
rect 36838 800 36854 856
rect 37022 800 37038 856
rect 37206 800 37314 856
rect 37482 800 37498 856
rect 37666 800 37682 856
rect 37850 800 37866 856
rect 38034 800 38050 856
rect 38218 800 38326 856
rect 38494 800 38510 856
rect 38678 800 38694 856
rect 38862 800 38878 856
rect 39046 800 39154 856
rect 39322 800 39338 856
rect 39506 800 39522 856
rect 39690 800 39706 856
rect 39874 800 39890 856
rect 40058 800 40166 856
rect 40334 800 40350 856
rect 40518 800 40534 856
rect 40702 800 40718 856
rect 40886 800 40902 856
rect 41070 800 41178 856
rect 41346 800 41362 856
rect 41530 800 41546 856
rect 41714 800 41730 856
rect 41898 800 42006 856
rect 42174 800 42190 856
rect 42358 800 42374 856
rect 42542 800 42558 856
rect 42726 800 42742 856
rect 42910 800 43018 856
rect 43186 800 43202 856
rect 43370 800 43386 856
rect 43554 800 43570 856
rect 43738 800 43754 856
rect 43922 800 44030 856
rect 44198 800 44214 856
rect 44382 800 44398 856
rect 44566 800 44582 856
rect 44750 800 44858 856
rect 45026 800 45042 856
rect 45210 800 45226 856
rect 45394 800 45410 856
rect 45578 800 45594 856
rect 45762 800 45870 856
rect 46038 800 46054 856
rect 46222 800 46238 856
rect 46406 800 46422 856
rect 46590 800 46606 856
rect 46774 800 46882 856
rect 47050 800 47066 856
rect 47234 800 47250 856
rect 47418 800 47434 856
rect 47602 800 47710 856
rect 47878 800 47894 856
rect 48062 800 48078 856
rect 48246 800 48262 856
rect 48430 800 48446 856
rect 48614 800 48722 856
rect 48890 800 48906 856
rect 49074 800 49090 856
rect 49258 800 49274 856
rect 49442 800 49458 856
rect 49626 800 49734 856
rect 49902 800 49918 856
rect 50086 800 50102 856
rect 50270 800 50286 856
rect 50454 800 50562 856
rect 50730 800 50746 856
rect 50914 800 50930 856
rect 51098 800 51114 856
rect 51282 800 51298 856
rect 51466 800 51574 856
rect 51742 800 51758 856
rect 51926 800 51942 856
rect 52110 800 52126 856
rect 52294 800 52310 856
rect 52478 800 52586 856
rect 52754 800 52770 856
rect 52938 800 52954 856
rect 53122 800 53138 856
rect 53306 800 53414 856
rect 53582 800 53598 856
rect 53766 800 53782 856
rect 53950 800 53966 856
rect 54134 800 54150 856
rect 54318 800 54426 856
rect 54594 800 54610 856
rect 54778 800 54794 856
rect 54962 800 54978 856
rect 55146 800 55162 856
rect 55330 800 55438 856
rect 55606 800 55622 856
rect 55790 800 55806 856
rect 55974 800 55990 856
rect 56158 800 56266 856
rect 56434 800 56450 856
rect 56618 800 56634 856
rect 56802 800 56818 856
rect 56986 800 57002 856
rect 57170 800 57278 856
rect 57446 800 57462 856
rect 57630 800 57646 856
rect 57814 800 57830 856
rect 57998 800 58014 856
rect 58182 800 58290 856
rect 58458 800 58474 856
rect 58642 800 58658 856
rect 58826 800 58842 856
rect 59010 800 59118 856
rect 59286 800 59302 856
rect 59470 800 59486 856
rect 59654 800 59670 856
rect 59838 800 59854 856
rect 60022 800 60130 856
rect 60298 800 60314 856
rect 60482 800 60498 856
rect 60666 800 60682 856
rect 60850 800 60866 856
rect 61034 800 61142 856
rect 61310 800 61326 856
rect 61494 800 61510 856
rect 61678 800 61694 856
rect 61862 800 61970 856
rect 62138 800 62154 856
rect 62322 800 62338 856
rect 62506 800 62522 856
rect 62690 800 62706 856
rect 62874 800 62982 856
rect 63150 800 63166 856
rect 63334 800 63350 856
rect 63518 800 63534 856
rect 63702 800 63718 856
rect 63886 800 63994 856
rect 64162 800 64178 856
rect 64346 800 64362 856
rect 64530 800 64546 856
rect 64714 800 64822 856
rect 64990 800 65006 856
rect 65174 800 65190 856
rect 65358 800 65374 856
rect 65542 800 65558 856
rect 65726 800 65834 856
rect 66002 800 66018 856
rect 66186 800 66202 856
rect 66370 800 66386 856
rect 66554 800 66570 856
rect 66738 800 66846 856
rect 67014 800 67030 856
rect 67198 800 67214 856
rect 67382 800 67398 856
rect 67566 800 67582 856
rect 67750 800 67858 856
rect 68026 800 68042 856
rect 68210 800 68226 856
rect 68394 800 68410 856
rect 68578 800 68686 856
rect 68854 800 68870 856
rect 69038 800 69054 856
rect 69222 800 69238 856
rect 69406 800 69422 856
rect 69590 800 69698 856
rect 69866 800 69882 856
rect 70050 800 70066 856
rect 70234 800 70250 856
rect 70418 800 70434 856
rect 70602 800 70710 856
rect 70878 800 70894 856
rect 71062 800 71078 856
rect 71246 800 71262 856
rect 71430 800 71538 856
rect 71706 800 71722 856
rect 71890 800 71906 856
rect 72074 800 72090 856
rect 72258 800 72274 856
rect 72442 800 72550 856
rect 72718 800 72734 856
rect 72902 800 72918 856
rect 73086 800 73102 856
rect 73270 800 73286 856
rect 73454 800 73562 856
rect 73730 800 73746 856
rect 73914 800 73930 856
rect 74098 800 74114 856
rect 74282 800 74390 856
rect 74558 800 74574 856
rect 74742 800 74758 856
rect 74926 800 74942 856
rect 75110 800 75126 856
rect 75294 800 75402 856
rect 75570 800 75586 856
rect 75754 800 75770 856
rect 75938 800 75954 856
rect 76122 800 76138 856
rect 76306 800 76414 856
rect 76582 800 76598 856
rect 76766 800 76782 856
rect 76950 800 76966 856
rect 77134 800 77242 856
rect 77410 800 77426 856
rect 77594 800 77610 856
rect 77778 800 77794 856
rect 77962 800 77978 856
rect 78146 800 78254 856
rect 78422 800 78438 856
rect 78606 800 78622 856
rect 78790 800 78806 856
rect 78974 800 78990 856
rect 79158 800 79266 856
rect 79434 800 79450 856
rect 79618 800 79634 856
rect 79802 800 79818 856
rect 79986 800 80094 856
rect 80262 800 80278 856
rect 80446 800 80462 856
rect 80630 800 80646 856
rect 80814 800 80830 856
rect 80998 800 81106 856
rect 81274 800 81290 856
rect 81458 800 81474 856
rect 81642 800 81658 856
rect 81826 800 81842 856
rect 82010 800 82118 856
rect 82286 800 82302 856
rect 82470 800 82486 856
rect 82654 800 82670 856
rect 82838 800 82946 856
rect 83114 800 83130 856
rect 83298 800 83314 856
rect 83482 800 83498 856
rect 83666 800 83682 856
rect 83850 800 83958 856
rect 84126 800 84142 856
rect 84310 800 84326 856
rect 84494 800 84510 856
rect 84678 800 84694 856
rect 84862 800 84970 856
rect 85138 800 85154 856
rect 85322 800 85338 856
rect 85506 800 85522 856
rect 85690 800 85798 856
rect 85966 800 85982 856
rect 86150 800 86166 856
rect 86334 800 86350 856
rect 86518 800 86534 856
rect 86702 800 86810 856
rect 86978 800 86994 856
rect 87162 800 87178 856
rect 87346 800 87362 856
rect 87530 800 87546 856
rect 87714 800 87822 856
rect 87990 800 88006 856
rect 88174 800 88190 856
rect 88358 800 88374 856
rect 88542 800 88650 856
rect 88818 800 88834 856
rect 89002 800 89018 856
rect 89186 800 89202 856
rect 89370 800 89386 856
rect 89554 800 89662 856
rect 89830 800 89846 856
rect 90014 800 90030 856
rect 90198 800 90214 856
rect 90382 800 90398 856
rect 90566 800 90674 856
rect 90842 800 90858 856
rect 91026 800 91042 856
rect 91210 800 91226 856
rect 91394 800 91502 856
rect 91670 800 91686 856
rect 91854 800 91870 856
rect 92038 800 92054 856
rect 92222 800 92238 856
rect 92406 800 92514 856
rect 92682 800 92698 856
rect 92866 800 92882 856
rect 93050 800 93066 856
rect 93234 800 93250 856
rect 93418 800 93526 856
rect 93694 800 93710 856
rect 93878 800 93894 856
rect 94062 800 94078 856
rect 94246 800 94354 856
rect 94522 800 94538 856
rect 94706 800 94722 856
rect 94890 800 94906 856
rect 95074 800 95090 856
rect 95258 800 95366 856
rect 95534 800 95550 856
rect 95718 800 95734 856
rect 95902 800 95918 856
rect 96086 800 96102 856
rect 96270 800 96378 856
rect 96546 800 96562 856
rect 96730 800 96746 856
rect 96914 800 96930 856
rect 97098 800 97206 856
rect 97374 800 97390 856
rect 97558 800 97574 856
rect 97742 800 97758 856
rect 97926 800 97942 856
rect 98110 800 98218 856
rect 98386 800 98402 856
rect 98570 800 98586 856
rect 98754 800 98770 856
rect 98938 800 98954 856
rect 99122 800 99230 856
rect 99398 800 99414 856
rect 99582 800 99598 856
rect 99766 800 99782 856
<< metal3 >>
rect 0 74808 800 74928
rect 0 24896 800 25016
<< obsm3 >>
rect 800 75008 96688 97409
rect 880 74728 96688 75008
rect 800 25096 96688 74728
rect 880 24816 96688 25096
rect 800 2143 96688 24816
<< metal4 >>
rect 4208 2128 4528 97424
rect 4868 2176 5188 97376
rect 5528 2176 5848 97376
rect 6188 2176 6508 97376
rect 19568 2128 19888 97424
rect 20228 2176 20548 97376
rect 20888 2176 21208 97376
rect 21548 2176 21868 97376
rect 34928 2128 35248 97424
rect 35588 2176 35908 97376
rect 36248 2176 36568 97376
rect 36908 2176 37228 97376
rect 50288 2128 50608 97424
rect 50948 2176 51268 97376
rect 51608 2176 51928 97376
rect 52268 2176 52588 97376
rect 65648 2128 65968 97424
rect 66308 2176 66628 97376
rect 66968 2176 67288 97376
rect 67628 2176 67948 97376
rect 81008 2128 81328 97424
rect 81668 2176 81988 97376
rect 82328 2176 82648 97376
rect 82988 2176 83308 97376
rect 96368 2128 96688 97424
rect 97028 2176 97348 97376
rect 97688 2176 98008 97376
<< labels >>
rlabel metal2 s 386 99200 442 100000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 26422 99200 26478 100000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 28998 99200 29054 100000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 31666 99200 31722 100000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 34242 99200 34298 100000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 36818 99200 36874 100000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 39486 99200 39542 100000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 42062 99200 42118 100000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 44730 99200 44786 100000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 47306 99200 47362 100000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 49882 99200 49938 100000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2962 99200 3018 100000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 52550 99200 52606 100000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 55126 99200 55182 100000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 57702 99200 57758 100000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 60370 99200 60426 100000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 62946 99200 63002 100000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 65522 99200 65578 100000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 68190 99200 68246 100000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 70766 99200 70822 100000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 73342 99200 73398 100000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 76010 99200 76066 100000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5538 99200 5594 100000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 78586 99200 78642 100000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 81254 99200 81310 100000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 83830 99200 83886 100000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 86406 99200 86462 100000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 89074 99200 89130 100000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 91650 99200 91706 100000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 94226 99200 94282 100000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 96894 99200 96950 100000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8206 99200 8262 100000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10782 99200 10838 100000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13358 99200 13414 100000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 16026 99200 16082 100000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 18602 99200 18658 100000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 21178 99200 21234 100000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 23846 99200 23902 100000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1214 99200 1270 100000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 27342 99200 27398 100000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 29918 99200 29974 100000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 32494 99200 32550 100000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 35162 99200 35218 100000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 37738 99200 37794 100000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 40314 99200 40370 100000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 42982 99200 43038 100000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 45558 99200 45614 100000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 48134 99200 48190 100000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 50802 99200 50858 100000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3790 99200 3846 100000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 53378 99200 53434 100000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 55954 99200 56010 100000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 58622 99200 58678 100000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 61198 99200 61254 100000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 63866 99200 63922 100000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 66442 99200 66498 100000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 69018 99200 69074 100000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 71686 99200 71742 100000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 74262 99200 74318 100000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 76838 99200 76894 100000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6458 99200 6514 100000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 79506 99200 79562 100000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 82082 99200 82138 100000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 84658 99200 84714 100000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 87326 99200 87382 100000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 89902 99200 89958 100000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 92478 99200 92534 100000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 95146 99200 95202 100000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 97722 99200 97778 100000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9034 99200 9090 100000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 11610 99200 11666 100000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 14278 99200 14334 100000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 16854 99200 16910 100000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 19430 99200 19486 100000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 22098 99200 22154 100000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 24674 99200 24730 100000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2042 99200 2098 100000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 28170 99200 28226 100000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 30746 99200 30802 100000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 33414 99200 33470 100000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 35990 99200 36046 100000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 38566 99200 38622 100000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 41234 99200 41290 100000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 43810 99200 43866 100000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 46386 99200 46442 100000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 49054 99200 49110 100000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 51630 99200 51686 100000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4710 99200 4766 100000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 54298 99200 54354 100000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 56874 99200 56930 100000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 59450 99200 59506 100000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 62118 99200 62174 100000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 64694 99200 64750 100000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 67270 99200 67326 100000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 69938 99200 69994 100000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 72514 99200 72570 100000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 75090 99200 75146 100000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 77758 99200 77814 100000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7286 99200 7342 100000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 80334 99200 80390 100000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 82910 99200 82966 100000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 85578 99200 85634 100000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 88154 99200 88210 100000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 90822 99200 90878 100000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 93398 99200 93454 100000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 95974 99200 96030 100000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 98642 99200 98698 100000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9862 99200 9918 100000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 12530 99200 12586 100000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 15106 99200 15162 100000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 17774 99200 17830 100000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 20350 99200 20406 100000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 22926 99200 22982 100000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 25594 99200 25650 100000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 99470 99200 99526 100000 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 user_clock2
port 502 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 503 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 504 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 505 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[0]
port 506 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[10]
port 507 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[11]
port 508 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[12]
port 509 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[13]
port 510 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_adr_i[14]
port 511 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[15]
port 512 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[16]
port 513 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[17]
port 514 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[18]
port 515 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_adr_i[19]
port 516 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[1]
port 517 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[20]
port 518 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[21]
port 519 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[22]
port 520 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[23]
port 521 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[24]
port 522 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[25]
port 523 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[26]
port 524 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[27]
port 525 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[28]
port 526 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[29]
port 527 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 528 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_adr_i[30]
port 529 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[31]
port 530 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[3]
port 531 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[4]
port 532 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[5]
port 533 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[6]
port 534 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[7]
port 535 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[8]
port 536 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[9]
port 537 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 538 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 539 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[10]
port 540 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[11]
port 541 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[12]
port 542 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[13]
port 543 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[14]
port 544 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[15]
port 545 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[16]
port 546 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_i[17]
port 547 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[18]
port 548 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[19]
port 549 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[1]
port 550 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_i[20]
port 551 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[21]
port 552 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[22]
port 553 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_i[23]
port 554 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[24]
port 555 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[25]
port 556 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[26]
port 557 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[27]
port 558 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[28]
port 559 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[29]
port 560 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[2]
port 561 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[30]
port 562 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_i[31]
port 563 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_i[3]
port 564 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[4]
port 565 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[5]
port 566 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[6]
port 567 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[7]
port 568 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[8]
port 569 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[9]
port 570 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 571 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[10]
port 572 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[11]
port 573 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[12]
port 574 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[13]
port 575 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[14]
port 576 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[15]
port 577 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[16]
port 578 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[17]
port 579 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[18]
port 580 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[19]
port 581 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[1]
port 582 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[20]
port 583 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_o[21]
port 584 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[22]
port 585 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[23]
port 586 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[24]
port 587 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[25]
port 588 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[26]
port 589 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[27]
port 590 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[28]
port 591 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_o[29]
port 592 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[2]
port 593 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[30]
port 594 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_o[31]
port 595 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[3]
port 596 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[4]
port 597 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[5]
port 598 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[6]
port 599 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_o[7]
port 600 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[8]
port 601 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[9]
port 602 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 603 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 604 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[2]
port 605 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_sel_i[3]
port 606 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 607 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 608 nsew signal input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 613 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 97028 2176 97348 97376 6 vccd2
port 616 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 97376 6 vccd2
port 617 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 97376 6 vccd2
port 618 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 97376 6 vccd2
port 619 nsew power bidirectional
rlabel metal4 s 81668 2176 81988 97376 6 vssd2
port 620 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 97376 6 vssd2
port 621 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 97376 6 vssd2
port 622 nsew ground bidirectional
rlabel metal4 s 97688 2176 98008 97376 6 vdda1
port 623 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 97376 6 vdda1
port 624 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 97376 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 97376 6 vdda1
port 626 nsew power bidirectional
rlabel metal4 s 82328 2176 82648 97376 6 vssa1
port 627 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 97376 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 97376 6 vssa1
port 629 nsew ground bidirectional
rlabel metal4 s 67628 2176 67948 97376 6 vdda2
port 630 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 97376 6 vdda2
port 631 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 97376 6 vdda2
port 632 nsew power bidirectional
rlabel metal4 s 82988 2176 83308 97376 6 vssa2
port 633 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 97376 6 vssa2
port 634 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 97376 6 vssa2
port 635 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 100000 100000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 2535208
string GDS_START 126
<< end >>

