magic
tech sky130A
magscale 1 2
timestamp 1623855674
<< locali >>
rect 74733 89879 74767 90049
rect 8309 88995 8343 89097
rect 14197 84983 14231 85221
rect 87613 83963 87647 84201
rect 96353 83963 96387 84201
rect 43269 76959 43303 77129
rect 25605 76279 25639 76449
rect 42993 59483 43027 59653
rect 41153 51255 41187 51425
rect 22293 49759 22327 49861
rect 86969 46495 87003 46665
rect 33149 39287 33183 39593
rect 25881 37655 25915 37893
rect 87337 37859 87371 37961
rect 27169 37655 27203 37757
rect 74365 31195 74399 31297
rect 27353 29699 27387 29801
rect 27445 29495 27479 29597
rect 48145 27863 48179 28101
rect 77125 27387 77159 27489
rect 59369 23035 59403 23205
rect 59311 23001 59403 23035
rect 61393 22967 61427 23069
rect 48237 19159 48271 19261
rect 96721 18615 96755 18717
rect 16681 14875 16715 14977
rect 71605 14807 71639 14909
rect 69213 12767 69247 12869
rect 79977 11611 80011 11713
rect 17141 10115 17175 10217
rect 16773 8347 16807 8517
rect 97273 2907 97307 3145
rect 84761 2499 84795 2601
<< viali >>
rect 2329 97257 2363 97291
rect 4445 97257 4479 97291
rect 7113 97257 7147 97291
rect 9781 97257 9815 97291
rect 12449 97257 12483 97291
rect 17785 97257 17819 97291
rect 20453 97257 20487 97291
rect 23121 97257 23155 97291
rect 28457 97257 28491 97291
rect 29929 97257 29963 97291
rect 31125 97257 31159 97291
rect 32597 97257 32631 97291
rect 34437 97257 34471 97291
rect 35265 97257 35299 97291
rect 37933 97257 37967 97291
rect 40601 97257 40635 97291
rect 43177 97257 43211 97291
rect 90465 97257 90499 97291
rect 95709 97257 95743 97291
rect 2973 97189 3007 97223
rect 4353 97189 4387 97223
rect 10885 97189 10919 97223
rect 15209 97189 15243 97223
rect 16129 97189 16163 97223
rect 18705 97189 18739 97223
rect 23581 97189 23615 97223
rect 23857 97189 23891 97223
rect 24685 97189 24719 97223
rect 26525 97189 26559 97223
rect 29101 97189 29135 97223
rect 31769 97189 31803 97223
rect 36921 97189 36955 97223
rect 39589 97189 39623 97223
rect 42165 97189 42199 97223
rect 44833 97189 44867 97223
rect 47409 97189 47443 97223
rect 48513 97189 48547 97223
rect 51089 97189 51123 97223
rect 53665 97189 53699 97223
rect 56333 97189 56367 97223
rect 57805 97189 57839 97223
rect 58909 97189 58943 97223
rect 60473 97189 60507 97223
rect 61577 97189 61611 97223
rect 64153 97189 64187 97223
rect 65717 97189 65751 97223
rect 66729 97189 66763 97223
rect 68569 97189 68603 97223
rect 69489 97189 69523 97223
rect 72709 97189 72743 97223
rect 74641 97189 74675 97223
rect 76389 97189 76423 97223
rect 77493 97189 77527 97223
rect 80161 97189 80195 97223
rect 82369 97189 82403 97223
rect 84669 97189 84703 97223
rect 87337 97189 87371 97223
rect 89913 97189 89947 97223
rect 90833 97189 90867 97223
rect 92489 97189 92523 97223
rect 95157 97189 95191 97223
rect 96077 97189 96111 97223
rect 97733 97189 97767 97223
rect 1409 97121 1443 97155
rect 2237 97121 2271 97155
rect 5549 97121 5583 97155
rect 7021 97121 7055 97155
rect 8217 97121 8251 97155
rect 9689 97121 9723 97155
rect 12357 97121 12391 97155
rect 13369 97121 13403 97155
rect 15025 97121 15059 97155
rect 17693 97121 17727 97155
rect 20361 97121 20395 97155
rect 21189 97121 21223 97155
rect 23029 97121 23063 97155
rect 24501 97121 24535 97155
rect 25789 97121 25823 97155
rect 28365 97121 28399 97155
rect 29837 97121 29871 97155
rect 31033 97121 31067 97155
rect 32505 97121 32539 97155
rect 34253 97121 34287 97155
rect 35173 97121 35207 97155
rect 37841 97121 37875 97155
rect 40509 97121 40543 97155
rect 43085 97121 43119 97155
rect 45661 97121 45695 97155
rect 48329 97121 48363 97155
rect 49893 97121 49927 97155
rect 50905 97121 50939 97155
rect 52561 97121 52595 97155
rect 53481 97121 53515 97155
rect 55137 97121 55171 97155
rect 56149 97121 56183 97155
rect 58725 97121 58759 97155
rect 61393 97121 61427 97155
rect 62957 97121 62991 97155
rect 63969 97121 64003 97155
rect 66545 97121 66579 97155
rect 68293 97121 68327 97155
rect 69305 97121 69339 97155
rect 71053 97121 71087 97155
rect 71789 97121 71823 97155
rect 72525 97121 72559 97155
rect 73629 97121 73663 97155
rect 74457 97121 74491 97155
rect 75193 97121 75227 97155
rect 77309 97121 77343 97155
rect 78965 97121 78999 97155
rect 79977 97121 80011 97155
rect 82185 97121 82219 97155
rect 82921 97121 82955 97155
rect 84577 97121 84611 97155
rect 84853 97121 84887 97155
rect 85497 97121 85531 97155
rect 87521 97121 87555 97155
rect 88165 97121 88199 97155
rect 90097 97121 90131 97155
rect 92673 97121 92707 97155
rect 93133 97121 93167 97155
rect 93409 97121 93443 97155
rect 95341 97121 95375 97155
rect 97917 97121 97951 97155
rect 5733 97053 5767 97087
rect 8493 97053 8527 97087
rect 13645 97053 13679 97087
rect 21373 97053 21407 97087
rect 25973 97053 26007 97087
rect 50077 97053 50111 97087
rect 55321 97053 55355 97087
rect 79149 97053 79183 97087
rect 85681 97053 85715 97087
rect 47593 96985 47627 97019
rect 57989 96985 58023 97019
rect 65901 96985 65935 97019
rect 73813 96985 73847 97019
rect 88349 96985 88383 97019
rect 90649 96985 90683 97019
rect 93225 96985 93259 97019
rect 95893 96985 95927 97019
rect 1593 96917 1627 96951
rect 3065 96917 3099 96951
rect 11161 96917 11195 96951
rect 16221 96917 16255 96951
rect 18797 96917 18831 96951
rect 23765 96917 23799 96951
rect 24317 96917 24351 96951
rect 26617 96917 26651 96951
rect 29193 96917 29227 96951
rect 31861 96917 31895 96951
rect 37197 96917 37231 96951
rect 39681 96917 39715 96951
rect 42257 96917 42291 96951
rect 44925 96917 44959 96951
rect 45753 96917 45787 96951
rect 52745 96917 52779 96951
rect 60749 96917 60783 96951
rect 63141 96917 63175 96951
rect 71145 96917 71179 96951
rect 71881 96917 71915 96951
rect 75285 96917 75319 96951
rect 76481 96917 76515 96951
rect 83013 96917 83047 96951
rect 85037 96917 85071 96951
rect 87245 96917 87279 96951
rect 87705 96917 87739 96951
rect 89729 96917 89763 96951
rect 92305 96917 92339 96951
rect 92857 96917 92891 96951
rect 94973 96917 95007 96951
rect 95525 96917 95559 96951
rect 97549 96917 97583 96951
rect 98101 96917 98135 96951
rect 16037 96713 16071 96747
rect 16313 96713 16347 96747
rect 2329 96577 2363 96611
rect 4997 96577 5031 96611
rect 7297 96577 7331 96611
rect 10149 96577 10183 96611
rect 12817 96577 12851 96611
rect 15393 96577 15427 96611
rect 18061 96577 18095 96611
rect 23213 96577 23247 96611
rect 25881 96577 25915 96611
rect 33701 96577 33735 96611
rect 36277 96577 36311 96611
rect 38853 96577 38887 96611
rect 41521 96577 41555 96611
rect 44097 96577 44131 96611
rect 49341 96577 49375 96611
rect 51917 96577 51951 96611
rect 54585 96577 54619 96611
rect 57161 96577 57195 96611
rect 59737 96577 59771 96611
rect 62405 96577 62439 96611
rect 64981 96577 65015 96611
rect 75377 96577 75411 96611
rect 93409 96577 93443 96611
rect 96261 96577 96295 96611
rect 98101 96577 98135 96611
rect 23857 96509 23891 96543
rect 43913 96509 43947 96543
rect 46305 96509 46339 96543
rect 46627 96509 46661 96543
rect 46765 96509 46799 96543
rect 47041 96509 47075 96543
rect 47225 96509 47259 96543
rect 70777 96509 70811 96543
rect 81265 96509 81299 96543
rect 83841 96509 83875 96543
rect 86417 96509 86451 96543
rect 89085 96509 89119 96543
rect 91661 96509 91695 96543
rect 94237 96509 94271 96543
rect 97365 96509 97399 96543
rect 2145 96441 2179 96475
rect 4813 96441 4847 96475
rect 7481 96441 7515 96475
rect 9965 96441 9999 96475
rect 12633 96441 12667 96475
rect 15209 96441 15243 96475
rect 17877 96441 17911 96475
rect 23029 96441 23063 96475
rect 25697 96441 25731 96475
rect 33517 96441 33551 96475
rect 36093 96441 36127 96475
rect 38669 96441 38703 96475
rect 41337 96441 41371 96475
rect 49157 96441 49191 96475
rect 51733 96441 51767 96475
rect 54401 96441 54435 96475
rect 56977 96441 57011 96475
rect 59553 96441 59587 96475
rect 62221 96441 62255 96475
rect 64797 96441 64831 96475
rect 75193 96441 75227 96475
rect 93593 96441 93627 96475
rect 96077 96441 96111 96475
rect 97181 96441 97215 96475
rect 97733 96441 97767 96475
rect 97917 96441 97951 96475
rect 98193 96441 98227 96475
rect 7113 96373 7147 96407
rect 24041 96373 24075 96407
rect 47501 96373 47535 96407
rect 70961 96373 70995 96407
rect 81449 96373 81483 96407
rect 93225 96373 93259 96407
rect 93777 96373 93811 96407
rect 96905 96373 96939 96407
rect 97457 96373 97491 96407
rect 46581 96169 46615 96203
rect 26525 96033 26559 96067
rect 46489 96033 46523 96067
rect 57437 96033 57471 96067
rect 57805 96033 57839 96067
rect 58173 96033 58207 96067
rect 83381 96033 83415 96067
rect 83749 96033 83783 96067
rect 96905 96033 96939 96067
rect 26801 95965 26835 95999
rect 28181 95965 28215 95999
rect 57621 95965 57655 95999
rect 58081 95965 58115 95999
rect 82921 95965 82955 95999
rect 83841 95965 83875 95999
rect 58541 95897 58575 95931
rect 53849 95557 53883 95591
rect 54217 95557 54251 95591
rect 35081 95489 35115 95523
rect 10149 95421 10183 95455
rect 34989 95421 35023 95455
rect 35357 95421 35391 95455
rect 35541 95421 35575 95455
rect 10885 95353 10919 95387
rect 34621 95285 34655 95319
rect 15117 95013 15151 95047
rect 2237 94945 2271 94979
rect 2421 94945 2455 94979
rect 2513 94945 2547 94979
rect 5089 94945 5123 94979
rect 14933 94945 14967 94979
rect 15209 94945 15243 94979
rect 15353 94945 15387 94979
rect 54125 94945 54159 94979
rect 54493 94945 54527 94979
rect 54585 94877 54619 94911
rect 1869 94809 1903 94843
rect 53941 94809 53975 94843
rect 2053 94741 2087 94775
rect 5181 94741 5215 94775
rect 15485 94741 15519 94775
rect 62773 94537 62807 94571
rect 25513 94333 25547 94367
rect 25789 94333 25823 94367
rect 41613 94333 41647 94367
rect 41889 94333 41923 94367
rect 54585 94333 54619 94367
rect 62957 94333 62991 94367
rect 63233 94333 63267 94367
rect 54401 94265 54435 94299
rect 63417 94265 63451 94299
rect 63049 94197 63083 94231
rect 95713 93925 95747 93959
rect 95525 93857 95559 93891
rect 95801 93857 95835 93891
rect 95985 93857 96019 93891
rect 96169 93653 96203 93687
rect 92581 92293 92615 92327
rect 93777 92293 93811 92327
rect 92673 92225 92707 92259
rect 93869 92225 93903 92259
rect 36369 92157 36403 92191
rect 92452 92157 92486 92191
rect 93648 92157 93682 92191
rect 23489 92089 23523 92123
rect 23673 92089 23707 92123
rect 36277 92089 36311 92123
rect 92305 92089 92339 92123
rect 93501 92089 93535 92123
rect 92949 92021 92983 92055
rect 94145 92021 94179 92055
rect 47317 91681 47351 91715
rect 47500 91681 47534 91715
rect 47590 91681 47624 91715
rect 47685 91681 47719 91715
rect 47869 91681 47903 91715
rect 73629 91681 73663 91715
rect 73812 91681 73846 91715
rect 73905 91681 73939 91715
rect 74181 91681 74215 91715
rect 73997 91613 74031 91647
rect 74365 91545 74399 91579
rect 47961 91477 47995 91511
rect 73445 91477 73479 91511
rect 44097 91069 44131 91103
rect 97733 91069 97767 91103
rect 97917 91069 97951 91103
rect 44281 90933 44315 90967
rect 9505 90593 9539 90627
rect 69857 90593 69891 90627
rect 70317 90525 70351 90559
rect 9689 90389 9723 90423
rect 52285 90389 52319 90423
rect 52469 90389 52503 90423
rect 45293 90117 45327 90151
rect 75101 90117 75135 90151
rect 29561 90049 29595 90083
rect 29653 90049 29687 90083
rect 74733 90049 74767 90083
rect 74917 90049 74951 90083
rect 29285 89981 29319 90015
rect 29468 89981 29502 90015
rect 29837 89981 29871 90015
rect 30481 89981 30515 90015
rect 30757 89981 30791 90015
rect 43913 89981 43947 90015
rect 44180 89913 44214 89947
rect 75280 89981 75314 90015
rect 75469 89981 75503 90015
rect 75653 89981 75687 90015
rect 75377 89913 75411 89947
rect 76205 89913 76239 89947
rect 29929 89845 29963 89879
rect 32045 89845 32079 89879
rect 74733 89845 74767 89879
rect 75745 89845 75779 89879
rect 76297 89845 76331 89879
rect 73813 89505 73847 89539
rect 74181 89505 74215 89539
rect 74549 89505 74583 89539
rect 88809 89505 88843 89539
rect 89177 89505 89211 89539
rect 73997 89437 74031 89471
rect 74641 89437 74675 89471
rect 88257 89437 88291 89471
rect 88625 89437 88659 89471
rect 89085 89437 89119 89471
rect 74917 89369 74951 89403
rect 8309 89097 8343 89131
rect 3893 89029 3927 89063
rect 6745 88961 6779 88995
rect 8309 88961 8343 88995
rect 2513 88893 2547 88927
rect 2780 88893 2814 88927
rect 7297 88893 7331 88927
rect 7573 88893 7607 88927
rect 7665 88893 7699 88927
rect 7941 88893 7975 88927
rect 8217 88893 8251 88927
rect 17693 88893 17727 88927
rect 17969 88893 18003 88927
rect 55045 88893 55079 88927
rect 55873 88825 55907 88859
rect 6929 88757 6963 88791
rect 19073 88757 19107 88791
rect 16037 88553 16071 88587
rect 15853 88417 15887 88451
rect 67281 88349 67315 88383
rect 67557 88349 67591 88383
rect 77585 87941 77619 87975
rect 8309 87805 8343 87839
rect 8585 87805 8619 87839
rect 15669 87805 15703 87839
rect 77677 87805 77711 87839
rect 77953 87805 77987 87839
rect 15945 87737 15979 87771
rect 79057 87669 79091 87703
rect 2053 87329 2087 87363
rect 2422 87329 2456 87363
rect 2605 87329 2639 87363
rect 27905 87329 27939 87363
rect 73169 87329 73203 87363
rect 73537 87329 73571 87363
rect 73905 87329 73939 87363
rect 74089 87329 74123 87363
rect 89913 87329 89947 87363
rect 90281 87329 90315 87363
rect 90649 87329 90683 87363
rect 2237 87261 2271 87295
rect 2329 87261 2363 87295
rect 28457 87261 28491 87295
rect 73629 87261 73663 87295
rect 90097 87261 90131 87295
rect 90557 87261 90591 87295
rect 1777 87193 1811 87227
rect 74273 87193 74307 87227
rect 89821 87193 89855 87227
rect 91017 87193 91051 87227
rect 1961 87125 1995 87159
rect 12357 86785 12391 86819
rect 12909 86785 12943 86819
rect 12081 86717 12115 86751
rect 12449 86717 12483 86751
rect 12817 86717 12851 86751
rect 29469 86717 29503 86751
rect 29745 86717 29779 86751
rect 55873 86717 55907 86751
rect 56149 86717 56183 86751
rect 31125 86649 31159 86683
rect 13277 86581 13311 86615
rect 43545 86241 43579 86275
rect 44189 86173 44223 86207
rect 82829 86173 82863 86207
rect 84301 86173 84335 86207
rect 84577 86173 84611 86207
rect 83013 86037 83047 86071
rect 89821 86037 89855 86071
rect 89913 86037 89947 86071
rect 97457 86037 97491 86071
rect 97733 86037 97767 86071
rect 80989 85629 81023 85663
rect 81265 85629 81299 85663
rect 87245 85629 87279 85663
rect 23673 85561 23707 85595
rect 24409 85561 24443 85595
rect 87061 85561 87095 85595
rect 14197 85221 14231 85255
rect 4721 85153 4755 85187
rect 5089 85153 5123 85187
rect 10149 85153 10183 85187
rect 10517 85153 10551 85187
rect 5181 85085 5215 85119
rect 9597 85085 9631 85119
rect 10241 85085 10275 85119
rect 10425 85085 10459 85119
rect 4537 85017 4571 85051
rect 31861 85153 31895 85187
rect 46305 85153 46339 85187
rect 46488 85153 46522 85187
rect 46673 85153 46707 85187
rect 46857 85153 46891 85187
rect 72525 85153 72559 85187
rect 32505 85085 32539 85119
rect 46581 85085 46615 85119
rect 47041 85085 47075 85119
rect 73077 85085 73111 85119
rect 14197 84949 14231 84983
rect 61761 84949 61795 84983
rect 61945 84949 61979 84983
rect 38485 84745 38519 84779
rect 62037 84541 62071 84575
rect 62313 84541 62347 84575
rect 85773 84541 85807 84575
rect 85957 84405 85991 84439
rect 87613 84201 87647 84235
rect 85865 84065 85899 84099
rect 86233 84065 86267 84099
rect 85313 83997 85347 84031
rect 85681 83997 85715 84031
rect 86141 83997 86175 84031
rect 87613 83929 87647 83963
rect 96353 84201 96387 84235
rect 97181 84065 97215 84099
rect 97549 84065 97583 84099
rect 96997 83997 97031 84031
rect 97457 83997 97491 84031
rect 96353 83929 96387 83963
rect 34529 83861 34563 83895
rect 34805 83861 34839 83895
rect 96813 83861 96847 83895
rect 19349 83453 19383 83487
rect 19625 83453 19659 83487
rect 97917 83385 97951 83419
rect 98009 83317 98043 83351
rect 76205 82977 76239 83011
rect 76573 82977 76607 83011
rect 75653 82909 75687 82943
rect 76021 82909 76055 82943
rect 76481 82909 76515 82943
rect 65349 82365 65383 82399
rect 65625 82365 65659 82399
rect 93685 82025 93719 82059
rect 74089 81889 74123 81923
rect 83013 81889 83047 81923
rect 94145 81889 94179 81923
rect 74457 81821 74491 81855
rect 83289 81821 83323 81855
rect 93869 81821 93903 81855
rect 41245 81685 41279 81719
rect 95249 81685 95283 81719
rect 27813 81277 27847 81311
rect 29837 81209 29871 81243
rect 82461 81209 82495 81243
rect 82737 81209 82771 81243
rect 83105 81209 83139 81243
rect 27629 81141 27663 81175
rect 29929 81141 29963 81175
rect 74089 80869 74123 80903
rect 84301 80869 84335 80903
rect 73905 80801 73939 80835
rect 84669 80733 84703 80767
rect 84577 80665 84611 80699
rect 73629 80597 73663 80631
rect 84466 80597 84500 80631
rect 84761 80597 84795 80631
rect 50261 80257 50295 80291
rect 29101 80189 29135 80223
rect 29377 80189 29411 80223
rect 49617 80189 49651 80223
rect 49801 80189 49835 80223
rect 49985 80189 50019 80223
rect 50353 80189 50387 80223
rect 30665 80053 30699 80087
rect 50813 80053 50847 80087
rect 42901 79781 42935 79815
rect 42625 79713 42659 79747
rect 42809 79713 42843 79747
rect 42998 79713 43032 79747
rect 43194 79713 43228 79747
rect 89085 79713 89119 79747
rect 89233 79713 89267 79747
rect 89453 79713 89487 79747
rect 89637 79713 89671 79747
rect 89361 79645 89395 79679
rect 89821 79577 89855 79611
rect 42533 79509 42567 79543
rect 43453 79509 43487 79543
rect 88993 79509 89027 79543
rect 89913 79509 89947 79543
rect 3249 79169 3283 79203
rect 4077 79169 4111 79203
rect 4445 79169 4479 79203
rect 97365 79169 97399 79203
rect 3985 79101 4019 79135
rect 4353 79101 4387 79135
rect 4721 79101 4755 79135
rect 28181 79101 28215 79135
rect 28457 79101 28491 79135
rect 96721 79101 96755 79135
rect 96905 79101 96939 79135
rect 97089 79101 97123 79135
rect 97457 79101 97491 79135
rect 3433 79033 3467 79067
rect 97917 78965 97951 78999
rect 30757 78693 30791 78727
rect 11069 78625 11103 78659
rect 11529 78625 11563 78659
rect 17325 78625 17359 78659
rect 17509 78625 17543 78659
rect 17729 78625 17763 78659
rect 17877 78625 17911 78659
rect 30481 78625 30515 78659
rect 30665 78625 30699 78659
rect 30854 78625 30888 78659
rect 83105 78625 83139 78659
rect 11253 78557 11287 78591
rect 17601 78557 17635 78591
rect 30389 78557 30423 78591
rect 83289 78557 83323 78591
rect 18061 78489 18095 78523
rect 17049 78421 17083 78455
rect 17233 78421 17267 78455
rect 31033 78421 31067 78455
rect 84301 78421 84335 78455
rect 84577 78421 84611 78455
rect 23397 78013 23431 78047
rect 23673 78013 23707 78047
rect 78413 78013 78447 78047
rect 78689 78013 78723 78047
rect 82737 78013 82771 78047
rect 82921 78013 82955 78047
rect 83105 78013 83139 78047
rect 77033 77945 77067 77979
rect 82277 77945 82311 77979
rect 76849 77877 76883 77911
rect 20729 77605 20763 77639
rect 25973 77537 26007 77571
rect 26156 77537 26190 77571
rect 26341 77537 26375 77571
rect 26525 77537 26559 77571
rect 21557 77469 21591 77503
rect 26249 77469 26283 77503
rect 25881 77333 25915 77367
rect 26617 77333 26651 77367
rect 28273 77129 28307 77163
rect 43269 77129 43303 77163
rect 43361 77129 43395 77163
rect 20729 77061 20763 77095
rect 28457 76925 28491 76959
rect 28641 76925 28675 76959
rect 28825 76925 28859 76959
rect 29193 76925 29227 76959
rect 29377 76925 29411 76959
rect 43269 76925 43303 76959
rect 43545 76925 43579 76959
rect 43821 76925 43855 76959
rect 54217 76925 54251 76959
rect 54493 76925 54527 76959
rect 93133 76925 93167 76959
rect 20545 76857 20579 76891
rect 29653 76789 29687 76823
rect 92949 76789 92983 76823
rect 58081 76585 58115 76619
rect 25605 76449 25639 76483
rect 26157 76449 26191 76483
rect 30573 76449 30607 76483
rect 56977 76449 57011 76483
rect 94053 76449 94087 76483
rect 25881 76381 25915 76415
rect 31125 76381 31159 76415
rect 56701 76381 56735 76415
rect 93777 76381 93811 76415
rect 25605 76245 25639 76279
rect 25697 76245 25731 76279
rect 27261 76245 27295 76279
rect 37473 76245 37507 76279
rect 37565 76245 37599 76279
rect 93593 76245 93627 76279
rect 95157 76245 95191 76279
rect 4905 75973 4939 76007
rect 44557 75905 44591 75939
rect 5089 75837 5123 75871
rect 5273 75837 5307 75871
rect 5457 75837 5491 75871
rect 30021 75837 30055 75871
rect 44097 75837 44131 75871
rect 30297 75769 30331 75803
rect 94973 75157 95007 75191
rect 95157 75157 95191 75191
rect 2605 74817 2639 74851
rect 2881 74749 2915 74783
rect 72617 74749 72651 74783
rect 72765 74749 72799 74783
rect 72893 74749 72927 74783
rect 72985 74749 73019 74783
rect 73169 74749 73203 74783
rect 77953 74681 77987 74715
rect 4169 74613 4203 74647
rect 73261 74613 73295 74647
rect 78045 74613 78079 74647
rect 76573 74341 76607 74375
rect 51457 74273 51491 74307
rect 51640 74273 51674 74307
rect 51733 74273 51767 74307
rect 52009 74273 52043 74307
rect 56701 74273 56735 74307
rect 78321 74273 78355 74307
rect 51825 74205 51859 74239
rect 56977 74205 57011 74239
rect 78505 74205 78539 74239
rect 52101 74069 52135 74103
rect 58081 74069 58115 74103
rect 76849 73593 76883 73627
rect 76941 73525 76975 73559
rect 46213 73185 46247 73219
rect 47041 73185 47075 73219
rect 13277 72641 13311 72675
rect 82921 72641 82955 72675
rect 13553 72573 13587 72607
rect 83197 72573 83231 72607
rect 14657 72437 14691 72471
rect 84301 72437 84335 72471
rect 30849 72233 30883 72267
rect 60197 72165 60231 72199
rect 9597 72097 9631 72131
rect 31309 72097 31343 72131
rect 55045 72097 55079 72131
rect 55229 72097 55263 72131
rect 55321 72097 55355 72131
rect 59829 72097 59863 72131
rect 59922 72097 59956 72131
rect 60105 72097 60139 72131
rect 60294 72097 60328 72131
rect 79149 72097 79183 72131
rect 31033 72029 31067 72063
rect 78873 72029 78907 72063
rect 9689 71893 9723 71927
rect 25145 71893 25179 71927
rect 25421 71893 25455 71927
rect 32413 71893 32447 71927
rect 54861 71893 54895 71927
rect 60473 71893 60507 71927
rect 78689 71893 78723 71927
rect 80253 71893 80287 71927
rect 89269 71893 89303 71927
rect 89453 71893 89487 71927
rect 71237 71621 71271 71655
rect 65901 71553 65935 71587
rect 22477 71485 22511 71519
rect 22753 71485 22787 71519
rect 54309 71485 54343 71519
rect 65349 71485 65383 71519
rect 66545 71485 66579 71519
rect 70685 71485 70719 71519
rect 70869 71485 70903 71519
rect 71105 71485 71139 71519
rect 54033 71417 54067 71451
rect 70961 71417 70995 71451
rect 66637 71349 66671 71383
rect 26801 71077 26835 71111
rect 26525 71009 26559 71043
rect 26709 71009 26743 71043
rect 26898 71009 26932 71043
rect 2513 70873 2547 70907
rect 2789 70873 2823 70907
rect 27077 70873 27111 70907
rect 25421 70805 25455 70839
rect 25697 70805 25731 70839
rect 83565 70805 83599 70839
rect 83749 70805 83783 70839
rect 52745 70465 52779 70499
rect 53021 70465 53055 70499
rect 87153 70465 87187 70499
rect 85313 70397 85347 70431
rect 86877 70397 86911 70431
rect 85589 70261 85623 70295
rect 15761 69921 15795 69955
rect 15945 69785 15979 69819
rect 2421 69445 2455 69479
rect 61301 69377 61335 69411
rect 61485 69377 61519 69411
rect 52561 69309 52595 69343
rect 88717 69309 88751 69343
rect 2053 69241 2087 69275
rect 2237 69241 2271 69275
rect 52469 69173 52503 69207
rect 88625 69173 88659 69207
rect 77493 68969 77527 69003
rect 85957 68969 85991 69003
rect 15945 68833 15979 68867
rect 77677 68833 77711 68867
rect 78045 68833 78079 68867
rect 78137 68833 78171 68867
rect 78413 68833 78447 68867
rect 90373 68833 90407 68867
rect 92029 68833 92063 68867
rect 16497 68765 16531 68799
rect 61945 68765 61979 68799
rect 62221 68765 62255 68799
rect 78321 68765 78355 68799
rect 84577 68765 84611 68799
rect 84853 68765 84887 68799
rect 91753 68765 91787 68799
rect 78781 68697 78815 68731
rect 63509 68629 63543 68663
rect 90189 68629 90223 68663
rect 92581 68425 92615 68459
rect 10057 68289 10091 68323
rect 46489 68289 46523 68323
rect 46581 68289 46615 68323
rect 6745 68221 6779 68255
rect 7021 68221 7055 68255
rect 9781 68221 9815 68255
rect 10149 68221 10183 68255
rect 10517 68221 10551 68255
rect 10701 68221 10735 68255
rect 46121 68221 46155 68255
rect 46305 68221 46339 68255
rect 46674 68221 46708 68255
rect 46857 68221 46891 68255
rect 92029 68221 92063 68255
rect 92213 68221 92247 68255
rect 92397 68221 92431 68255
rect 92305 68153 92339 68187
rect 10977 68085 11011 68119
rect 45937 68085 45971 68119
rect 16129 67745 16163 67779
rect 44005 67745 44039 67779
rect 16957 67677 16991 67711
rect 44833 67677 44867 67711
rect 90649 67609 90683 67643
rect 90925 67609 90959 67643
rect 3617 67337 3651 67371
rect 33793 67269 33827 67303
rect 52193 67269 52227 67303
rect 4160 67201 4194 67235
rect 19717 67201 19751 67235
rect 20637 67201 20671 67235
rect 3893 67133 3927 67167
rect 4077 67133 4111 67167
rect 4261 67133 4295 67167
rect 4441 67133 4475 67167
rect 4629 67133 4663 67167
rect 19533 67133 19567 67167
rect 19901 67133 19935 67167
rect 20269 67133 20303 67167
rect 20453 67133 20487 67167
rect 33977 67133 34011 67167
rect 52377 67133 52411 67167
rect 63141 67133 63175 67167
rect 63417 67133 63451 67167
rect 72709 67133 72743 67167
rect 86141 67133 86175 67167
rect 90741 67133 90775 67167
rect 3709 67065 3743 67099
rect 52653 67065 52687 67099
rect 73261 67065 73295 67099
rect 86417 67065 86451 67099
rect 91017 67065 91051 67099
rect 52561 66997 52595 67031
rect 34161 66793 34195 66827
rect 20453 66657 20487 66691
rect 77953 66657 77987 66691
rect 4261 66589 4295 66623
rect 4537 66589 4571 66623
rect 32781 66589 32815 66623
rect 33057 66589 33091 66623
rect 5825 66521 5859 66555
rect 20269 66453 20303 66487
rect 64889 66453 64923 66487
rect 65073 66453 65107 66487
rect 77953 66453 77987 66487
rect 80161 66113 80195 66147
rect 80253 66045 80287 66079
rect 80529 66045 80563 66079
rect 82369 66045 82403 66079
rect 82553 66045 82587 66079
rect 82737 66045 82771 66079
rect 83105 66045 83139 66079
rect 83289 66045 83323 66079
rect 81633 65909 81667 65943
rect 83565 65909 83599 65943
rect 6653 65569 6687 65603
rect 7389 65569 7423 65603
rect 81725 65569 81759 65603
rect 7113 65501 7147 65535
rect 81541 65433 81575 65467
rect 90557 65161 90591 65195
rect 80161 65093 80195 65127
rect 80437 65093 80471 65127
rect 60381 65025 60415 65059
rect 92397 65025 92431 65059
rect 27813 64957 27847 64991
rect 59277 64957 59311 64991
rect 59461 64957 59495 64991
rect 59645 64957 59679 64991
rect 60013 64957 60047 64991
rect 60197 64957 60231 64991
rect 90741 64957 90775 64991
rect 92121 64957 92155 64991
rect 28641 64889 28675 64923
rect 27353 64617 27387 64651
rect 50537 64617 50571 64651
rect 27169 64481 27203 64515
rect 49433 64481 49467 64515
rect 49715 64481 49749 64515
rect 49892 64481 49926 64515
rect 49985 64481 50019 64515
rect 50261 64481 50295 64515
rect 91569 64481 91603 64515
rect 91753 64481 91787 64515
rect 91845 64481 91879 64515
rect 92029 64481 92063 64515
rect 95065 64481 95099 64515
rect 95433 64481 95467 64515
rect 95801 64481 95835 64515
rect 50077 64413 50111 64447
rect 92213 64413 92247 64447
rect 95249 64413 95283 64447
rect 95709 64413 95743 64447
rect 26157 64277 26191 64311
rect 26433 64277 26467 64311
rect 49617 64277 49651 64311
rect 50353 64277 50387 64311
rect 67189 64277 67223 64311
rect 67373 64277 67407 64311
rect 96261 64277 96295 64311
rect 8953 64073 8987 64107
rect 66361 64073 66395 64107
rect 68477 64073 68511 64107
rect 82461 64005 82495 64039
rect 67097 63937 67131 63971
rect 8309 63869 8343 63903
rect 8492 63869 8526 63903
rect 8585 63869 8619 63903
rect 8677 63869 8711 63903
rect 8861 63869 8895 63903
rect 66545 63869 66579 63903
rect 67373 63869 67407 63903
rect 81909 63869 81943 63903
rect 82185 63869 82219 63903
rect 82282 63869 82316 63903
rect 93133 63869 93167 63903
rect 82093 63801 82127 63835
rect 66913 63733 66947 63767
rect 92949 63733 92983 63767
rect 18613 63393 18647 63427
rect 27445 63393 27479 63427
rect 27261 63257 27295 63291
rect 9413 63189 9447 63223
rect 9689 63189 9723 63223
rect 18797 63189 18831 63223
rect 44649 63189 44683 63223
rect 44925 63189 44959 63223
rect 79701 63189 79735 63223
rect 79885 63189 79919 63223
rect 13553 62917 13587 62951
rect 14197 62849 14231 62883
rect 13737 62781 13771 62815
rect 14105 62781 14139 62815
rect 33793 62781 33827 62815
rect 33976 62781 34010 62815
rect 34069 62781 34103 62815
rect 34161 62781 34195 62815
rect 34345 62781 34379 62815
rect 33701 62645 33735 62679
rect 34437 62645 34471 62679
rect 13001 62305 13035 62339
rect 13185 62305 13219 62339
rect 13277 62305 13311 62339
rect 73997 62305 74031 62339
rect 74365 62305 74399 62339
rect 74733 62305 74767 62339
rect 74917 62305 74951 62339
rect 83473 62305 83507 62339
rect 74273 62237 74307 62271
rect 83749 62237 83783 62271
rect 75101 62169 75135 62203
rect 12817 62101 12851 62135
rect 75009 61897 75043 61931
rect 30665 61761 30699 61795
rect 50721 61761 50755 61795
rect 30481 61693 30515 61727
rect 30849 61693 30883 61727
rect 31217 61693 31251 61727
rect 31401 61693 31435 61727
rect 48789 61693 48823 61727
rect 50997 61693 51031 61727
rect 75193 61693 75227 61727
rect 83289 61693 83323 61727
rect 93225 61693 93259 61727
rect 49617 61625 49651 61659
rect 83657 61625 83691 61659
rect 31677 61557 31711 61591
rect 52101 61557 52135 61591
rect 93409 61557 93443 61591
rect 9505 61217 9539 61251
rect 9781 61217 9815 61251
rect 41153 61217 41187 61251
rect 41429 61217 41463 61251
rect 41705 61217 41739 61251
rect 41797 61217 41831 61251
rect 57621 61217 57655 61251
rect 92029 61217 92063 61251
rect 41981 61149 42015 61183
rect 57897 61149 57931 61183
rect 92213 61149 92247 61183
rect 4169 61013 4203 61047
rect 4445 61013 4479 61047
rect 11069 61013 11103 61047
rect 59001 61013 59035 61047
rect 75009 61013 75043 61047
rect 75285 61013 75319 61047
rect 96997 61013 97031 61047
rect 97181 61013 97215 61047
rect 68109 60809 68143 60843
rect 75377 60673 75411 60707
rect 4997 60605 5031 60639
rect 5273 60605 5307 60639
rect 67557 60605 67591 60639
rect 67741 60605 67775 60639
rect 67833 60605 67867 60639
rect 67971 60605 68005 60639
rect 75101 60605 75135 60639
rect 83013 60605 83047 60639
rect 83197 60605 83231 60639
rect 83381 60605 83415 60639
rect 83657 60605 83691 60639
rect 83749 60605 83783 60639
rect 91753 60605 91787 60639
rect 92029 60605 92063 60639
rect 84209 60469 84243 60503
rect 5181 60129 5215 60163
rect 36553 60129 36587 60163
rect 74825 60129 74859 60163
rect 89821 60129 89855 60163
rect 6009 60061 6043 60095
rect 36277 60061 36311 60095
rect 75009 60061 75043 60095
rect 90005 60061 90039 60095
rect 37841 59925 37875 59959
rect 67189 59925 67223 59959
rect 67373 59925 67407 59959
rect 38117 59721 38151 59755
rect 42993 59653 43027 59687
rect 38577 59585 38611 59619
rect 18061 59517 18095 59551
rect 38301 59517 38335 59551
rect 38484 59517 38518 59551
rect 38669 59517 38703 59551
rect 38853 59517 38887 59551
rect 60749 59517 60783 59551
rect 61025 59517 61059 59551
rect 39037 59449 39071 59483
rect 42993 59449 43027 59483
rect 18245 59381 18279 59415
rect 60565 59381 60599 59415
rect 60933 59381 60967 59415
rect 37657 59177 37691 59211
rect 38025 59177 38059 59211
rect 93225 59177 93259 59211
rect 21281 59041 21315 59075
rect 37841 59041 37875 59075
rect 38117 59041 38151 59075
rect 21833 58973 21867 59007
rect 93409 58973 93443 59007
rect 93685 58973 93719 59007
rect 94789 58973 94823 59007
rect 37565 58837 37599 58871
rect 57621 58497 57655 58531
rect 57345 58429 57379 58463
rect 81173 58429 81207 58463
rect 81081 58293 81115 58327
rect 53941 57749 53975 57783
rect 54217 57749 54251 57783
rect 10333 57545 10367 57579
rect 10425 57409 10459 57443
rect 84209 57409 84243 57443
rect 10204 57341 10238 57375
rect 13737 57341 13771 57375
rect 14013 57341 14047 57375
rect 20729 57341 20763 57375
rect 21005 57341 21039 57375
rect 83933 57341 83967 57375
rect 85405 57341 85439 57375
rect 85681 57341 85715 57375
rect 10057 57273 10091 57307
rect 82553 57273 82587 57307
rect 10701 57205 10735 57239
rect 82369 57205 82403 57239
rect 64797 57001 64831 57035
rect 64061 56933 64095 56967
rect 64521 56933 64555 56967
rect 37473 56865 37507 56899
rect 64245 56865 64279 56899
rect 64429 56865 64463 56899
rect 64613 56865 64647 56899
rect 68753 56865 68787 56899
rect 96721 56865 96755 56899
rect 97181 56865 97215 56899
rect 97365 56865 97399 56899
rect 97549 56865 97583 56899
rect 38025 56797 38059 56831
rect 68937 56797 68971 56831
rect 59277 56661 59311 56695
rect 59553 56661 59587 56695
rect 3249 56253 3283 56287
rect 10885 56253 10919 56287
rect 33977 56253 34011 56287
rect 34253 56253 34287 56287
rect 42257 56253 42291 56287
rect 50445 56253 50479 56287
rect 50721 56253 50755 56287
rect 54217 56253 54251 56287
rect 54493 56253 54527 56287
rect 3801 56185 3835 56219
rect 41889 56185 41923 56219
rect 11069 56117 11103 56151
rect 35357 56117 35391 56151
rect 55781 56117 55815 56151
rect 49065 55777 49099 55811
rect 49213 55777 49247 55811
rect 49479 55777 49513 55811
rect 49617 55777 49651 55811
rect 49801 55777 49835 55811
rect 68569 55777 68603 55811
rect 49341 55709 49375 55743
rect 68845 55709 68879 55743
rect 44281 55233 44315 55267
rect 43637 55165 43671 55199
rect 44189 55165 44223 55199
rect 44465 55165 44499 55199
rect 61025 55165 61059 55199
rect 91937 55165 91971 55199
rect 61301 55097 61335 55131
rect 92765 55097 92799 55131
rect 84117 54757 84151 54791
rect 36553 54689 36587 54723
rect 83657 54689 83691 54723
rect 36277 54621 36311 54655
rect 86141 54621 86175 54655
rect 86417 54621 86451 54655
rect 37841 54485 37875 54519
rect 47777 54485 47811 54519
rect 48053 54485 48087 54519
rect 84577 54485 84611 54519
rect 84853 54485 84887 54519
rect 25421 54145 25455 54179
rect 24317 54077 24351 54111
rect 25605 54077 25639 54111
rect 25789 54009 25823 54043
rect 24041 53941 24075 53975
rect 53389 53669 53423 53703
rect 53757 53669 53791 53703
rect 53849 53669 53883 53703
rect 14749 53601 14783 53635
rect 21005 53601 21039 53635
rect 21188 53601 21222 53635
rect 21557 53601 21591 53635
rect 53573 53601 53607 53635
rect 53993 53601 54027 53635
rect 63141 53601 63175 53635
rect 75469 53601 75503 53635
rect 84945 53601 84979 53635
rect 15025 53533 15059 53567
rect 21281 53533 21315 53567
rect 21373 53533 21407 53567
rect 63509 53533 63543 53567
rect 75745 53533 75779 53567
rect 85221 53533 85255 53567
rect 16313 53465 16347 53499
rect 54309 53465 54343 53499
rect 21649 53397 21683 53431
rect 54125 53397 54159 53431
rect 58173 53125 58207 53159
rect 60473 53125 60507 53159
rect 61209 53125 61243 53159
rect 61485 53125 61519 53159
rect 67005 53125 67039 53159
rect 73629 53057 73663 53091
rect 81081 53057 81115 53091
rect 18797 52989 18831 53023
rect 57437 52989 57471 53023
rect 57585 52989 57619 53023
rect 57713 52989 57747 53023
rect 57805 52989 57839 53023
rect 57989 52989 58023 53023
rect 60657 52989 60691 53023
rect 60933 52989 60967 53023
rect 61077 52989 61111 53023
rect 66913 52989 66947 53023
rect 67189 52989 67223 53023
rect 73353 52989 73387 53023
rect 80805 52989 80839 53023
rect 19625 52921 19659 52955
rect 60841 52921 60875 52955
rect 71973 52921 72007 52955
rect 67373 52853 67407 52887
rect 71789 52853 71823 52887
rect 3985 52649 4019 52683
rect 4261 52649 4295 52683
rect 5181 52649 5215 52683
rect 7389 52649 7423 52683
rect 8033 52649 8067 52683
rect 7665 52581 7699 52615
rect 7757 52581 7791 52615
rect 42717 52581 42751 52615
rect 4445 52513 4479 52547
rect 4809 52513 4843 52547
rect 4997 52513 5031 52547
rect 7481 52513 7515 52547
rect 7849 52513 7883 52547
rect 36277 52513 36311 52547
rect 36645 52513 36679 52547
rect 37013 52513 37047 52547
rect 37197 52513 37231 52547
rect 42165 52513 42199 52547
rect 80161 52513 80195 52547
rect 80345 52513 80379 52547
rect 80529 52513 80563 52547
rect 80897 52513 80931 52547
rect 89637 52513 89671 52547
rect 4169 52445 4203 52479
rect 4629 52445 4663 52479
rect 4721 52445 4755 52479
rect 8125 52445 8159 52479
rect 36461 52445 36495 52479
rect 37381 52445 37415 52479
rect 80805 52445 80839 52479
rect 81265 52445 81299 52479
rect 89545 52445 89579 52479
rect 13553 52309 13587 52343
rect 13829 52309 13863 52343
rect 82829 52309 82863 52343
rect 82921 52309 82955 52343
rect 59461 52105 59495 52139
rect 9781 51901 9815 51935
rect 41797 51901 41831 51935
rect 54585 51901 54619 51935
rect 59277 51901 59311 51935
rect 10425 51833 10459 51867
rect 42073 51833 42107 51867
rect 55137 51833 55171 51867
rect 41153 51425 41187 51459
rect 41429 51425 41463 51459
rect 41613 51425 41647 51459
rect 42073 51357 42107 51391
rect 41153 51221 41187 51255
rect 41245 51221 41279 51255
rect 41705 51221 41739 51255
rect 77493 51221 77527 51255
rect 77677 51221 77711 51255
rect 47593 50813 47627 50847
rect 47501 50677 47535 50711
rect 21741 50473 21775 50507
rect 21925 50473 21959 50507
rect 48053 50405 48087 50439
rect 90649 50405 90683 50439
rect 21833 50337 21867 50371
rect 22109 50337 22143 50371
rect 37841 50337 37875 50371
rect 49617 50337 49651 50371
rect 58633 50337 58667 50371
rect 72617 50337 72651 50371
rect 90465 50337 90499 50371
rect 22477 50269 22511 50303
rect 31953 50269 31987 50303
rect 32229 50269 32263 50303
rect 73077 50269 73111 50303
rect 37657 50201 37691 50235
rect 58449 50201 58483 50235
rect 22293 50133 22327 50167
rect 33517 50133 33551 50167
rect 36185 50133 36219 50167
rect 36461 50133 36495 50167
rect 13461 49929 13495 49963
rect 22293 49861 22327 49895
rect 24041 49861 24075 49895
rect 70133 49861 70167 49895
rect 12725 49793 12759 49827
rect 1409 49725 1443 49759
rect 12265 49725 12299 49759
rect 12633 49725 12667 49759
rect 13001 49725 13035 49759
rect 13185 49725 13219 49759
rect 22293 49725 22327 49759
rect 22569 49725 22603 49759
rect 22753 49725 22787 49759
rect 22937 49725 22971 49759
rect 23213 49725 23247 49759
rect 23305 49725 23339 49759
rect 23857 49725 23891 49759
rect 30297 49725 30331 49759
rect 30573 49725 30607 49759
rect 31953 49725 31987 49759
rect 48789 49725 48823 49759
rect 49617 49725 49651 49759
rect 55965 49725 55999 49759
rect 71421 49725 71455 49759
rect 71697 49725 71731 49759
rect 56701 49657 56735 49691
rect 22385 49589 22419 49623
rect 69857 49589 69891 49623
rect 42349 49181 42383 49215
rect 42625 49181 42659 49215
rect 84209 49181 84243 49215
rect 85681 49181 85715 49215
rect 85957 49181 85991 49215
rect 84393 49113 84427 49147
rect 1501 49045 1535 49079
rect 1777 49045 1811 49079
rect 22385 49045 22419 49079
rect 22661 49045 22695 49079
rect 24041 49045 24075 49079
rect 24317 49045 24351 49079
rect 43729 49045 43763 49079
rect 18889 48705 18923 48739
rect 68017 48705 68051 48739
rect 18981 48637 19015 48671
rect 19257 48637 19291 48671
rect 19349 48637 19383 48671
rect 34253 48637 34287 48671
rect 67741 48637 67775 48671
rect 19165 48569 19199 48603
rect 35081 48569 35115 48603
rect 19533 48501 19567 48535
rect 4905 48161 4939 48195
rect 5273 48161 5307 48195
rect 5457 48161 5491 48195
rect 41797 48161 41831 48195
rect 57753 48161 57787 48195
rect 57897 48161 57931 48195
rect 57989 48161 58023 48195
rect 58173 48161 58207 48195
rect 4997 48093 5031 48127
rect 42073 48093 42107 48127
rect 43453 48093 43487 48127
rect 4537 47957 4571 47991
rect 37565 47957 37599 47991
rect 37841 47957 37875 47991
rect 46029 47957 46063 47991
rect 46213 47957 46247 47991
rect 57345 47957 57379 47991
rect 57621 47957 57655 47991
rect 58265 47957 58299 47991
rect 28457 47753 28491 47787
rect 92949 47753 92983 47787
rect 28181 47617 28215 47651
rect 92121 47617 92155 47651
rect 92489 47617 92523 47651
rect 92581 47617 92615 47651
rect 27813 47549 27847 47583
rect 27996 47549 28030 47583
rect 28089 47549 28123 47583
rect 28365 47549 28399 47583
rect 86969 47549 87003 47583
rect 87153 47549 87187 47583
rect 87337 47549 87371 47583
rect 87705 47549 87739 47583
rect 87889 47549 87923 47583
rect 92305 47549 92339 47583
rect 92674 47549 92708 47583
rect 92857 47549 92891 47583
rect 91937 47481 91971 47515
rect 27629 47413 27663 47447
rect 86785 47413 86819 47447
rect 88165 47413 88199 47447
rect 17693 47209 17727 47243
rect 64981 47141 65015 47175
rect 16313 47073 16347 47107
rect 64521 47073 64555 47107
rect 64705 47073 64739 47107
rect 64889 47073 64923 47107
rect 65078 47073 65112 47107
rect 75837 47073 75871 47107
rect 16589 47005 16623 47039
rect 76113 47005 76147 47039
rect 65257 46937 65291 46971
rect 86969 46665 87003 46699
rect 13369 46529 13403 46563
rect 14657 46529 14691 46563
rect 19257 46529 19291 46563
rect 87337 46529 87371 46563
rect 88257 46529 88291 46563
rect 14105 46461 14139 46495
rect 14197 46461 14231 46495
rect 14473 46461 14507 46495
rect 14841 46461 14875 46495
rect 18705 46461 18739 46495
rect 86969 46461 87003 46495
rect 87153 46461 87187 46495
rect 87521 46461 87555 46495
rect 87797 46461 87831 46495
rect 87889 46461 87923 46495
rect 13645 46325 13679 46359
rect 7481 45441 7515 45475
rect 76297 45441 76331 45475
rect 6929 45373 6963 45407
rect 76573 45373 76607 45407
rect 77677 45237 77711 45271
rect 18061 44965 18095 44999
rect 74273 44965 74307 44999
rect 6469 44897 6503 44931
rect 6837 44897 6871 44931
rect 17872 44897 17906 44931
rect 17969 44897 18003 44931
rect 18245 44897 18279 44931
rect 74089 44897 74123 44931
rect 74365 44897 74399 44931
rect 74462 44897 74496 44931
rect 17693 44761 17727 44795
rect 1685 44693 1719 44727
rect 1961 44693 1995 44727
rect 6653 44693 6687 44727
rect 17509 44693 17543 44727
rect 21741 44693 21775 44727
rect 22017 44693 22051 44727
rect 74641 44693 74675 44727
rect 23305 44285 23339 44319
rect 23581 44285 23615 44319
rect 58081 44285 58115 44319
rect 58357 44285 58391 44319
rect 69765 44285 69799 44319
rect 24869 44149 24903 44183
rect 69581 44149 69615 44183
rect 25237 43809 25271 43843
rect 25605 43741 25639 43775
rect 37289 43741 37323 43775
rect 37565 43741 37599 43775
rect 38853 43673 38887 43707
rect 23213 43605 23247 43639
rect 23489 43605 23523 43639
rect 40049 43333 40083 43367
rect 45109 43265 45143 43299
rect 59369 43265 59403 43299
rect 40233 43197 40267 43231
rect 40417 43197 40451 43231
rect 44741 43197 44775 43231
rect 59553 43197 59587 43231
rect 88717 43197 88751 43231
rect 40509 43129 40543 43163
rect 59829 43129 59863 43163
rect 59737 43061 59771 43095
rect 88533 43061 88567 43095
rect 73169 42721 73203 42755
rect 73537 42721 73571 42755
rect 73721 42721 73755 42755
rect 80529 42721 80563 42755
rect 91661 42721 91695 42755
rect 72525 42653 72559 42687
rect 73077 42653 73111 42687
rect 80713 42585 80747 42619
rect 91845 42585 91879 42619
rect 92857 42177 92891 42211
rect 44741 42109 44775 42143
rect 92581 42109 92615 42143
rect 44373 41973 44407 42007
rect 30481 41633 30515 41667
rect 48789 41633 48823 41667
rect 96353 41633 96387 41667
rect 96721 41633 96755 41667
rect 97089 41633 97123 41667
rect 97273 41633 97307 41667
rect 31309 41565 31343 41599
rect 49433 41565 49467 41599
rect 96169 41565 96203 41599
rect 96537 41565 96571 41599
rect 97457 41497 97491 41531
rect 90557 40681 90591 40715
rect 95525 40681 95559 40715
rect 92121 40545 92155 40579
rect 95433 40545 95467 40579
rect 92397 40477 92431 40511
rect 90833 40409 90867 40443
rect 77677 40341 77711 40375
rect 77861 40341 77895 40375
rect 32965 40069 32999 40103
rect 33241 40069 33275 40103
rect 41068 40001 41102 40035
rect 41521 40001 41555 40035
rect 50077 40001 50111 40035
rect 50261 40001 50295 40035
rect 59277 40001 59311 40035
rect 60933 40001 60967 40035
rect 71789 40001 71823 40035
rect 2789 39933 2823 39967
rect 28365 39933 28399 39967
rect 28641 39933 28675 39967
rect 34437 39933 34471 39967
rect 34621 39933 34655 39967
rect 34857 39933 34891 39967
rect 40785 39933 40819 39967
rect 40968 39933 41002 39967
rect 41153 39933 41187 39967
rect 41337 39933 41371 39967
rect 41613 39933 41647 39967
rect 50537 39933 50571 39967
rect 59093 39933 59127 39967
rect 59553 39933 59587 39967
rect 67741 39933 67775 39967
rect 68017 39933 68051 39967
rect 72065 39933 72099 39967
rect 3341 39865 3375 39899
rect 34713 39865 34747 39899
rect 29745 39797 29779 39831
rect 34997 39797 35031 39831
rect 40601 39797 40635 39831
rect 51641 39797 51675 39831
rect 73169 39797 73203 39831
rect 6193 39593 6227 39627
rect 33149 39593 33183 39627
rect 33333 39593 33367 39627
rect 34161 39593 34195 39627
rect 31677 39525 31711 39559
rect 5089 39457 5123 39491
rect 31125 39457 31159 39491
rect 32137 39457 32171 39491
rect 32689 39457 32723 39491
rect 32965 39457 32999 39491
rect 4813 39389 4847 39423
rect 32505 39389 32539 39423
rect 32873 39321 32907 39355
rect 33425 39457 33459 39491
rect 33609 39457 33643 39491
rect 33977 39457 34011 39491
rect 69029 39457 69063 39491
rect 33701 39389 33735 39423
rect 33793 39389 33827 39423
rect 33149 39253 33183 39287
rect 68937 39253 68971 39287
rect 33057 38777 33091 38811
rect 33885 38777 33919 38811
rect 33333 38505 33367 38539
rect 43177 38505 43211 38539
rect 32689 38437 32723 38471
rect 73261 38437 73295 38471
rect 10413 38369 10447 38403
rect 10701 38369 10735 38403
rect 10793 38369 10827 38403
rect 11069 38369 11103 38403
rect 11253 38369 11287 38403
rect 33241 38369 33275 38403
rect 42533 38369 42567 38403
rect 42716 38369 42750 38403
rect 42901 38369 42935 38403
rect 43085 38369 43119 38403
rect 46397 38369 46431 38403
rect 48145 38369 48179 38403
rect 31033 38301 31067 38335
rect 31309 38301 31343 38335
rect 42816 38301 42850 38335
rect 46673 38301 46707 38335
rect 73353 38301 73387 38335
rect 73629 38301 73663 38335
rect 74733 38301 74767 38335
rect 10057 38233 10091 38267
rect 48329 38233 48363 38267
rect 7297 38165 7331 38199
rect 7573 38165 7607 38199
rect 33793 38165 33827 38199
rect 34069 38165 34103 38199
rect 78413 37961 78447 37995
rect 87337 37961 87371 37995
rect 25881 37893 25915 37927
rect 47041 37893 47075 37927
rect 9137 37825 9171 37859
rect 9413 37757 9447 37791
rect 19625 37757 19659 37791
rect 19901 37757 19935 37791
rect 10793 37689 10827 37723
rect 46673 37825 46707 37859
rect 78965 37825 78999 37859
rect 81173 37825 81207 37859
rect 81449 37825 81483 37859
rect 87337 37825 87371 37859
rect 87705 37825 87739 37859
rect 87889 37825 87923 37859
rect 88441 37825 88475 37859
rect 26065 37757 26099 37791
rect 26341 37757 26375 37791
rect 27169 37757 27203 37791
rect 46121 37757 46155 37791
rect 46305 37757 46339 37791
rect 46488 37757 46522 37791
rect 46581 37757 46615 37791
rect 46857 37757 46891 37791
rect 50629 37757 50663 37791
rect 50905 37757 50939 37791
rect 73721 37757 73755 37791
rect 78597 37757 78631 37791
rect 78780 37757 78814 37791
rect 78873 37757 78907 37791
rect 79122 37757 79156 37791
rect 25881 37621 25915 37655
rect 87521 37689 87555 37723
rect 87981 37689 88015 37723
rect 27169 37621 27203 37655
rect 50445 37621 50479 37655
rect 50813 37621 50847 37655
rect 73537 37621 73571 37655
rect 79241 37621 79275 37655
rect 82553 37621 82587 37655
rect 88349 37621 88383 37655
rect 17601 37417 17635 37451
rect 12909 37349 12943 37383
rect 73537 37349 73571 37383
rect 78689 37349 78723 37383
rect 11253 37281 11287 37315
rect 11529 37281 11563 37315
rect 17785 37281 17819 37315
rect 18153 37281 18187 37315
rect 18337 37281 18371 37315
rect 18613 37281 18647 37315
rect 18705 37281 18739 37315
rect 19073 37281 19107 37315
rect 73997 37281 74031 37315
rect 74181 37281 74215 37315
rect 74549 37281 74583 37315
rect 77953 37281 77987 37315
rect 93869 37281 93903 37315
rect 94237 37281 94271 37315
rect 74457 37213 74491 37247
rect 94329 37213 94363 37247
rect 93685 37145 93719 37179
rect 84761 37077 84795 37111
rect 84853 37077 84887 37111
rect 3341 36873 3375 36907
rect 76205 36873 76239 36907
rect 3157 36737 3191 36771
rect 3525 36669 3559 36703
rect 3709 36669 3743 36703
rect 75009 36669 75043 36703
rect 75193 36669 75227 36703
rect 75377 36669 75411 36703
rect 75745 36669 75779 36703
rect 75929 36669 75963 36703
rect 87613 36669 87647 36703
rect 88441 36669 88475 36703
rect 90833 36669 90867 36703
rect 3801 36601 3835 36635
rect 91201 36601 91235 36635
rect 3985 36533 4019 36567
rect 88441 36533 88475 36567
rect 51273 36329 51307 36363
rect 78965 36261 78999 36295
rect 35817 36193 35851 36227
rect 51457 36193 51491 36227
rect 51640 36193 51674 36227
rect 51825 36193 51859 36227
rect 52009 36193 52043 36227
rect 52193 36193 52227 36227
rect 63049 36193 63083 36227
rect 63232 36193 63266 36227
rect 63601 36193 63635 36227
rect 77677 36193 77711 36227
rect 78045 36193 78079 36227
rect 78321 36193 78355 36227
rect 78413 36193 78447 36227
rect 36553 36125 36587 36159
rect 51733 36125 51767 36159
rect 63325 36125 63359 36159
rect 63417 36125 63451 36159
rect 77953 36125 77987 36159
rect 63693 35989 63727 36023
rect 75009 35581 75043 35615
rect 74825 35445 74859 35479
rect 27721 35105 27755 35139
rect 72433 35105 72467 35139
rect 27445 35037 27479 35071
rect 72249 35037 72283 35071
rect 72801 35037 72835 35071
rect 72709 34969 72743 35003
rect 29009 34901 29043 34935
rect 72571 34901 72605 34935
rect 73077 34901 73111 34935
rect 65901 34697 65935 34731
rect 66913 34629 66947 34663
rect 66545 34561 66579 34595
rect 66085 34493 66119 34527
rect 66269 34493 66303 34527
rect 66453 34493 66487 34527
rect 66638 34493 66672 34527
rect 66824 34493 66858 34527
rect 67833 34493 67867 34527
rect 68661 34493 68695 34527
rect 56609 34153 56643 34187
rect 21649 34085 21683 34119
rect 19993 34017 20027 34051
rect 36001 34017 36035 34051
rect 56701 34017 56735 34051
rect 56885 34017 56919 34051
rect 57069 34017 57103 34051
rect 57253 34017 57287 34051
rect 20269 33949 20303 33983
rect 56977 33949 57011 33983
rect 57529 33949 57563 33983
rect 36185 33881 36219 33915
rect 35817 33813 35851 33847
rect 57437 33813 57471 33847
rect 60013 33813 60047 33847
rect 60289 33813 60323 33847
rect 33057 33405 33091 33439
rect 33333 33405 33367 33439
rect 40509 33405 40543 33439
rect 40785 33405 40819 33439
rect 34713 33337 34747 33371
rect 58909 32997 58943 33031
rect 58081 32929 58115 32963
rect 30389 32725 30423 32759
rect 30665 32725 30699 32759
rect 10793 32521 10827 32555
rect 91937 32453 91971 32487
rect 92259 32453 92293 32487
rect 92397 32453 92431 32487
rect 2789 32385 2823 32419
rect 92489 32385 92523 32419
rect 3065 32317 3099 32351
rect 9229 32317 9263 32351
rect 9505 32317 9539 32351
rect 92121 32249 92155 32283
rect 4353 32181 4387 32215
rect 92765 32181 92799 32215
rect 95065 31977 95099 32011
rect 32045 31841 32079 31875
rect 32321 31841 32355 31875
rect 93869 31841 93903 31875
rect 94237 31841 94271 31875
rect 94605 31841 94639 31875
rect 41797 31773 41831 31807
rect 41981 31773 42015 31807
rect 43085 31773 43119 31807
rect 43361 31773 43395 31807
rect 44741 31773 44775 31807
rect 94053 31773 94087 31807
rect 94513 31773 94547 31807
rect 64613 31433 64647 31467
rect 70593 31297 70627 31331
rect 72801 31297 72835 31331
rect 74365 31297 74399 31331
rect 70317 31229 70351 31263
rect 71605 31229 71639 31263
rect 72525 31229 72559 31263
rect 74365 31161 74399 31195
rect 64429 31093 64463 31127
rect 71421 31093 71455 31127
rect 69489 30821 69523 30855
rect 9965 30753 9999 30787
rect 10333 30753 10367 30787
rect 10425 30753 10459 30787
rect 21097 30753 21131 30787
rect 67649 30753 67683 30787
rect 67833 30753 67867 30787
rect 68201 30753 68235 30787
rect 68569 30753 68603 30787
rect 69673 30753 69707 30787
rect 70041 30753 70075 30787
rect 70317 30753 70351 30787
rect 70409 30753 70443 30787
rect 21465 30685 21499 30719
rect 68385 30685 68419 30719
rect 69857 30685 69891 30719
rect 9781 30617 9815 30651
rect 67373 30617 67407 30651
rect 67097 30549 67131 30583
rect 70869 30549 70903 30583
rect 78505 30209 78539 30243
rect 41245 30141 41279 30175
rect 58081 30141 58115 30175
rect 77861 30141 77895 30175
rect 41613 30073 41647 30107
rect 58265 30005 58299 30039
rect 27353 29801 27387 29835
rect 21281 29733 21315 29767
rect 26617 29733 26651 29767
rect 26985 29733 27019 29767
rect 27261 29733 27295 29767
rect 20729 29665 20763 29699
rect 21925 29665 21959 29699
rect 26433 29665 26467 29699
rect 26801 29665 26835 29699
rect 27077 29665 27111 29699
rect 27353 29665 27387 29699
rect 27721 29665 27755 29699
rect 88809 29665 88843 29699
rect 88993 29665 89027 29699
rect 89158 29665 89192 29699
rect 89545 29665 89579 29699
rect 26249 29597 26283 29631
rect 27445 29597 27479 29631
rect 89269 29597 89303 29631
rect 89361 29597 89395 29631
rect 22201 29461 22235 29495
rect 27445 29461 27479 29495
rect 27537 29461 27571 29495
rect 89637 29461 89671 29495
rect 17325 29257 17359 29291
rect 25513 29257 25547 29291
rect 45293 29257 45327 29291
rect 75101 29189 75135 29223
rect 44925 29121 44959 29155
rect 46397 29121 46431 29155
rect 14473 29053 14507 29087
rect 17509 29053 17543 29087
rect 25237 29053 25271 29087
rect 25973 29053 26007 29087
rect 26065 29053 26099 29087
rect 26341 29053 26375 29087
rect 26525 29053 26559 29087
rect 26709 29053 26743 29087
rect 46673 29053 46707 29087
rect 75101 29053 75135 29087
rect 14841 28985 14875 29019
rect 15577 28645 15611 28679
rect 63509 28645 63543 28679
rect 63969 28645 64003 28679
rect 15393 28577 15427 28611
rect 15669 28577 15703 28611
rect 60381 28577 60415 28611
rect 63693 28577 63727 28611
rect 63877 28577 63911 28611
rect 77677 28577 77711 28611
rect 60657 28509 60691 28543
rect 77953 28509 77987 28543
rect 15209 28373 15243 28407
rect 43821 28101 43855 28135
rect 48145 28101 48179 28135
rect 44281 28033 44315 28067
rect 43545 27965 43579 27999
rect 44005 27965 44039 27999
rect 44189 27965 44223 27999
rect 44391 27965 44425 27999
rect 44557 27965 44591 27999
rect 44649 27897 44683 27931
rect 55965 28033 55999 28067
rect 55597 27965 55631 27999
rect 55780 27965 55814 27999
rect 55873 27965 55907 27999
rect 56149 27965 56183 27999
rect 82093 27965 82127 27999
rect 82369 27965 82403 27999
rect 43729 27829 43763 27863
rect 48145 27829 48179 27863
rect 56241 27829 56275 27863
rect 12817 27489 12851 27523
rect 13645 27489 13679 27523
rect 42441 27489 42475 27523
rect 42809 27489 42843 27523
rect 43085 27489 43119 27523
rect 43177 27489 43211 27523
rect 73445 27489 73479 27523
rect 74273 27489 74307 27523
rect 77125 27489 77159 27523
rect 77861 27489 77895 27523
rect 85405 27489 85439 27523
rect 14933 27421 14967 27455
rect 15209 27421 15243 27455
rect 25421 27421 25455 27455
rect 42717 27421 42751 27455
rect 43545 27421 43579 27455
rect 85589 27421 85623 27455
rect 77125 27353 77159 27387
rect 77677 27353 77711 27387
rect 16497 27285 16531 27319
rect 56609 27285 56643 27319
rect 56701 27285 56735 27319
rect 7021 27081 7055 27115
rect 87870 27013 87904 27047
rect 87981 27013 88015 27047
rect 88717 27013 88751 27047
rect 7573 26945 7607 26979
rect 20361 26945 20395 26979
rect 87429 26945 87463 26979
rect 88533 26945 88567 26979
rect 7481 26877 7515 26911
rect 7849 26877 7883 26911
rect 8033 26877 8067 26911
rect 8217 26877 8251 26911
rect 20177 26877 20211 26911
rect 20545 26877 20579 26911
rect 20913 26877 20947 26911
rect 21097 26877 21131 26911
rect 65349 26877 65383 26911
rect 87521 26877 87555 26911
rect 87705 26877 87739 26911
rect 88044 26877 88078 26911
rect 6745 26809 6779 26843
rect 21465 26809 21499 26843
rect 65165 26741 65199 26775
rect 88349 26741 88383 26775
rect 21833 26537 21867 26571
rect 20729 26401 20763 26435
rect 34713 26401 34747 26435
rect 20453 26333 20487 26367
rect 84761 26265 84795 26299
rect 96629 26265 96663 26299
rect 96721 26265 96755 26299
rect 34529 26197 34563 26231
rect 2881 25789 2915 25823
rect 49157 25789 49191 25823
rect 49801 25789 49835 25823
rect 75009 25789 75043 25823
rect 75837 25721 75871 25755
rect 80161 25381 80195 25415
rect 47777 25313 47811 25347
rect 80345 25313 80379 25347
rect 80528 25313 80562 25347
rect 80897 25313 80931 25347
rect 47961 25245 47995 25279
rect 78229 25245 78263 25279
rect 78505 25245 78539 25279
rect 80621 25245 80655 25279
rect 80713 25245 80747 25279
rect 37841 25109 37875 25143
rect 72617 25109 72651 25143
rect 79609 25109 79643 25143
rect 80989 25109 81023 25143
rect 9873 24905 9907 24939
rect 9965 24837 9999 24871
rect 9413 24769 9447 24803
rect 10057 24769 10091 24803
rect 10425 24769 10459 24803
rect 19625 24769 19659 24803
rect 9505 24701 9539 24735
rect 19717 24701 19751 24735
rect 19993 24701 20027 24735
rect 37105 24701 37139 24735
rect 59461 24701 59495 24735
rect 85497 24701 85531 24735
rect 85681 24701 85715 24735
rect 85865 24701 85899 24735
rect 86233 24701 86267 24735
rect 86417 24701 86451 24735
rect 36838 24633 36872 24667
rect 9137 24565 9171 24599
rect 10609 24565 10643 24599
rect 21281 24565 21315 24599
rect 35449 24565 35483 24599
rect 35725 24565 35759 24599
rect 85313 24565 85347 24599
rect 86693 24565 86727 24599
rect 6837 23681 6871 23715
rect 40785 23681 40819 23715
rect 7113 23613 7147 23647
rect 40049 23613 40083 23647
rect 77401 23613 77435 23647
rect 77585 23613 77619 23647
rect 77677 23613 77711 23647
rect 8493 23545 8527 23579
rect 77217 23545 77251 23579
rect 76941 23477 76975 23511
rect 59369 23205 59403 23239
rect 59553 23205 59587 23239
rect 59829 23137 59863 23171
rect 60013 23137 60047 23171
rect 60197 23137 60231 23171
rect 60381 23137 60415 23171
rect 60749 23137 60783 23171
rect 77677 23137 77711 23171
rect 60105 23069 60139 23103
rect 61393 23069 61427 23103
rect 77953 23069 77987 23103
rect 59277 23001 59311 23035
rect 60565 23001 60599 23035
rect 20085 22933 20119 22967
rect 20361 22933 20395 22967
rect 59737 22933 59771 22967
rect 61393 22933 61427 22967
rect 79241 22933 79275 22967
rect 84945 22933 84979 22967
rect 19165 22525 19199 22559
rect 19441 22525 19475 22559
rect 38485 22525 38519 22559
rect 45477 22525 45511 22559
rect 20821 22457 20855 22491
rect 36185 22117 36219 22151
rect 83013 22117 83047 22151
rect 36921 22049 36955 22083
rect 47501 22049 47535 22083
rect 47593 21981 47627 22015
rect 47869 21981 47903 22015
rect 48973 21845 49007 21879
rect 83105 21845 83139 21879
rect 36020 21641 36054 21675
rect 35909 21573 35943 21607
rect 35817 21505 35851 21539
rect 80621 21437 80655 21471
rect 80805 21437 80839 21471
rect 80989 21437 81023 21471
rect 81265 21437 81299 21471
rect 81357 21437 81391 21471
rect 35449 21369 35483 21403
rect 36185 21369 36219 21403
rect 35357 21301 35391 21335
rect 81817 21301 81851 21335
rect 77953 21029 77987 21063
rect 77677 20961 77711 20995
rect 94329 20961 94363 20995
rect 94605 20893 94639 20927
rect 94145 20757 94179 20791
rect 95709 20757 95743 20791
rect 24317 20417 24351 20451
rect 51273 20417 51307 20451
rect 3617 20349 3651 20383
rect 19533 20349 19567 20383
rect 23949 20349 23983 20383
rect 24132 20349 24166 20383
rect 24225 20349 24259 20383
rect 24501 20349 24535 20383
rect 50997 20349 51031 20383
rect 78137 20349 78171 20383
rect 19809 20281 19843 20315
rect 3801 20213 3835 20247
rect 23857 20213 23891 20247
rect 24593 20213 24627 20247
rect 52377 20213 52411 20247
rect 65165 20009 65199 20043
rect 88809 19941 88843 19975
rect 64981 19873 65015 19907
rect 72433 19873 72467 19907
rect 72893 19873 72927 19907
rect 73077 19873 73111 19907
rect 73261 19873 73295 19907
rect 90373 19873 90407 19907
rect 91109 19873 91143 19907
rect 90649 19805 90683 19839
rect 89085 19737 89119 19771
rect 91293 19669 91327 19703
rect 44925 19329 44959 19363
rect 4997 19261 5031 19295
rect 44649 19261 44683 19295
rect 44832 19261 44866 19295
rect 45017 19261 45051 19295
rect 45201 19261 45235 19295
rect 48237 19261 48271 19295
rect 50077 19261 50111 19295
rect 50629 19261 50663 19295
rect 5549 19193 5583 19227
rect 45293 19125 45327 19159
rect 48237 19125 48271 19159
rect 65165 18921 65199 18955
rect 49065 18853 49099 18887
rect 63601 18853 63635 18887
rect 64797 18853 64831 18887
rect 65257 18853 65291 18887
rect 47225 18785 47259 18819
rect 47685 18785 47719 18819
rect 62221 18785 62255 18819
rect 64981 18785 65015 18819
rect 96997 18785 97031 18819
rect 97181 18785 97215 18819
rect 97273 18785 97307 18819
rect 97549 18785 97583 18819
rect 47409 18717 47443 18751
rect 61945 18717 61979 18751
rect 96721 18717 96755 18751
rect 97365 18717 97399 18751
rect 97733 18649 97767 18683
rect 96721 18581 96755 18615
rect 96813 18581 96847 18615
rect 56609 18377 56643 18411
rect 73353 18377 73387 18411
rect 71329 18309 71363 18343
rect 19533 18241 19567 18275
rect 29929 18241 29963 18275
rect 70869 18241 70903 18275
rect 70961 18241 70995 18275
rect 19349 18173 19383 18207
rect 30205 18173 30239 18207
rect 31585 18173 31619 18207
rect 55045 18173 55079 18207
rect 55321 18173 55355 18207
rect 70409 18173 70443 18207
rect 70593 18173 70627 18207
rect 70765 18173 70799 18207
rect 71145 18173 71179 18207
rect 73169 18173 73203 18207
rect 17141 17493 17175 17527
rect 20453 17493 20487 17527
rect 32597 17493 32631 17527
rect 62129 17493 62163 17527
rect 87061 17153 87095 17187
rect 87153 17153 87187 17187
rect 14933 17085 14967 17119
rect 44557 17085 44591 17119
rect 86693 17085 86727 17119
rect 86877 17085 86911 17119
rect 87246 17085 87280 17119
rect 87429 17085 87463 17119
rect 97181 17085 97215 17119
rect 86509 16949 86543 16983
rect 44741 16745 44775 16779
rect 47685 16745 47719 16779
rect 8033 16677 8067 16711
rect 8493 16677 8527 16711
rect 44649 16677 44683 16711
rect 7849 16609 7883 16643
rect 8217 16609 8251 16643
rect 8401 16609 8435 16643
rect 48041 16609 48075 16643
rect 48329 16609 48363 16643
rect 48467 16609 48501 16643
rect 48697 16609 48731 16643
rect 48973 16609 49007 16643
rect 58081 15657 58115 15691
rect 57989 15589 58023 15623
rect 21925 15317 21959 15351
rect 22201 15317 22235 15351
rect 16681 14977 16715 15011
rect 71789 14977 71823 15011
rect 72065 14977 72099 15011
rect 13369 14909 13403 14943
rect 13645 14909 13679 14943
rect 13737 14909 13771 14943
rect 14013 14909 14047 14943
rect 14289 14909 14323 14943
rect 54769 14909 54803 14943
rect 71605 14909 71639 14943
rect 16681 14841 16715 14875
rect 54033 14841 54067 14875
rect 13001 14773 13035 14807
rect 71605 14773 71639 14807
rect 44373 14433 44407 14467
rect 44556 14433 44590 14467
rect 44741 14433 44775 14467
rect 44879 14433 44913 14467
rect 82921 14433 82955 14467
rect 44649 14365 44683 14399
rect 45293 14365 45327 14399
rect 44189 14297 44223 14331
rect 37749 14229 37783 14263
rect 45017 14229 45051 14263
rect 83105 14229 83139 14263
rect 8677 13957 8711 13991
rect 8861 13957 8895 13991
rect 9137 13957 9171 13991
rect 9321 13957 9355 13991
rect 20177 13821 20211 13855
rect 39773 13821 39807 13855
rect 39957 13685 39991 13719
rect 11529 13345 11563 13379
rect 11897 13345 11931 13379
rect 12173 13345 12207 13379
rect 12265 13345 12299 13379
rect 67373 13345 67407 13379
rect 11713 13277 11747 13311
rect 12725 13209 12759 13243
rect 16957 13141 16991 13175
rect 27721 13141 27755 13175
rect 52193 13141 52227 13175
rect 40601 12869 40635 12903
rect 40923 12869 40957 12903
rect 41061 12869 41095 12903
rect 69213 12869 69247 12903
rect 97825 12869 97859 12903
rect 41153 12801 41187 12835
rect 96629 12801 96663 12835
rect 96905 12801 96939 12835
rect 18429 12733 18463 12767
rect 19073 12733 19107 12767
rect 41705 12733 41739 12767
rect 66269 12733 66303 12767
rect 66637 12733 66671 12767
rect 66729 12733 66763 12767
rect 67005 12733 67039 12767
rect 67189 12733 67223 12767
rect 67557 12733 67591 12767
rect 69213 12733 69247 12767
rect 96721 12733 96755 12767
rect 97089 12733 97123 12767
rect 97365 12733 97399 12767
rect 97457 12733 97491 12767
rect 40785 12665 40819 12699
rect 41521 12665 41555 12699
rect 38117 12257 38151 12291
rect 38393 12257 38427 12291
rect 85773 12257 85807 12291
rect 85957 12257 85991 12291
rect 86141 12257 86175 12291
rect 86509 12257 86543 12291
rect 96353 12257 96387 12291
rect 96721 12257 96755 12291
rect 97089 12257 97123 12291
rect 86417 12189 86451 12223
rect 96813 12189 96847 12223
rect 96997 12189 97031 12223
rect 86877 12121 86911 12155
rect 39681 12053 39715 12087
rect 97549 12053 97583 12087
rect 3433 11849 3467 11883
rect 19533 11781 19567 11815
rect 80391 11781 80425 11815
rect 80529 11781 80563 11815
rect 3709 11713 3743 11747
rect 3801 11713 3835 11747
rect 79977 11713 80011 11747
rect 80069 11713 80103 11747
rect 80621 11713 80655 11747
rect 3525 11645 3559 11679
rect 3929 11645 3963 11679
rect 4077 11645 4111 11679
rect 3249 11577 3283 11611
rect 79977 11577 80011 11611
rect 80253 11577 80287 11611
rect 80897 11509 80931 11543
rect 26985 11305 27019 11339
rect 27169 11169 27203 11203
rect 27353 11169 27387 11203
rect 27721 11169 27755 11203
rect 27905 11169 27939 11203
rect 42901 11169 42935 11203
rect 53389 11169 53423 11203
rect 53573 11169 53607 11203
rect 53849 11169 53883 11203
rect 53942 11169 53976 11203
rect 54125 11169 54159 11203
rect 5733 11101 5767 11135
rect 6009 11101 6043 11135
rect 43177 11101 43211 11135
rect 53757 11101 53791 11135
rect 7297 11033 7331 11067
rect 44465 11033 44499 11067
rect 53205 11033 53239 11067
rect 36921 10693 36955 10727
rect 1685 10625 1719 10659
rect 3893 10625 3927 10659
rect 4537 10625 4571 10659
rect 12909 10625 12943 10659
rect 39865 10625 39899 10659
rect 40141 10625 40175 10659
rect 1961 10557 1995 10591
rect 4445 10557 4479 10591
rect 4813 10557 4847 10591
rect 4997 10557 5031 10591
rect 12081 10557 12115 10591
rect 24041 10557 24075 10591
rect 24685 10557 24719 10591
rect 36369 10557 36403 10591
rect 36645 10557 36679 10591
rect 36742 10557 36776 10591
rect 54677 10557 54711 10591
rect 54861 10557 54895 10591
rect 55045 10557 55079 10591
rect 55413 10557 55447 10591
rect 55597 10557 55631 10591
rect 36553 10489 36587 10523
rect 54493 10489 54527 10523
rect 3249 10421 3283 10455
rect 55873 10421 55907 10455
rect 17141 10217 17175 10251
rect 61761 10217 61795 10251
rect 62221 10217 62255 10251
rect 17141 10081 17175 10115
rect 17233 10081 17267 10115
rect 23581 10081 23615 10115
rect 63331 10081 63365 10115
rect 63594 10081 63628 10115
rect 91477 10081 91511 10115
rect 91753 10081 91787 10115
rect 17572 10013 17606 10047
rect 17398 9945 17432 9979
rect 17509 9877 17543 9911
rect 17877 9877 17911 9911
rect 23765 9877 23799 9911
rect 94237 9605 94271 9639
rect 45109 9469 45143 9503
rect 45293 9469 45327 9503
rect 45477 9469 45511 9503
rect 46489 9469 46523 9503
rect 61117 9469 61151 9503
rect 44649 9401 44683 9435
rect 94053 9401 94087 9435
rect 4813 8585 4847 8619
rect 13921 8517 13955 8551
rect 16773 8517 16807 8551
rect 4905 8381 4939 8415
rect 5089 8381 5123 8415
rect 4445 8313 4479 8347
rect 16773 8313 16807 8347
rect 64429 7973 64463 8007
rect 93869 7905 93903 7939
rect 94145 7905 94179 7939
rect 94238 7905 94272 7939
rect 94421 7905 94455 7939
rect 62773 7837 62807 7871
rect 63049 7837 63083 7871
rect 94053 7837 94087 7871
rect 93685 7769 93719 7803
rect 93501 7701 93535 7735
rect 94513 7701 94547 7735
rect 43729 7429 43763 7463
rect 13093 7293 13127 7327
rect 45017 7293 45051 7327
rect 45293 7293 45327 7327
rect 57345 7293 57379 7327
rect 57437 7293 57471 7327
rect 90925 7293 90959 7327
rect 43453 7157 43487 7191
rect 57805 7157 57839 7191
rect 50537 6817 50571 6851
rect 59921 6817 59955 6851
rect 97549 6817 97583 6851
rect 50261 6749 50295 6783
rect 60289 6749 60323 6783
rect 48973 6681 49007 6715
rect 60059 6681 60093 6715
rect 60197 6681 60231 6715
rect 48697 6613 48731 6647
rect 56977 6613 57011 6647
rect 59737 6613 59771 6647
rect 60565 6613 60599 6647
rect 81633 6613 81667 6647
rect 96905 6613 96939 6647
rect 92121 6409 92155 6443
rect 93685 6273 93719 6307
rect 14657 6205 14691 6239
rect 93961 6205 93995 6239
rect 96997 6205 97031 6239
rect 97641 6205 97675 6239
rect 92305 6137 92339 6171
rect 50353 5865 50387 5899
rect 85221 5865 85255 5899
rect 50261 5797 50295 5831
rect 91201 5797 91235 5831
rect 2697 5729 2731 5763
rect 84117 5729 84151 5763
rect 91661 5729 91695 5763
rect 91845 5729 91879 5763
rect 92029 5729 92063 5763
rect 96261 5729 96295 5763
rect 96905 5729 96939 5763
rect 97549 5729 97583 5763
rect 83841 5661 83875 5695
rect 2513 5117 2547 5151
rect 4077 5117 4111 5151
rect 4721 5117 4755 5151
rect 7021 5117 7055 5151
rect 10609 5117 10643 5151
rect 12081 5117 12115 5151
rect 13093 5117 13127 5151
rect 14289 5117 14323 5151
rect 15485 5117 15519 5151
rect 17325 5117 17359 5151
rect 18613 5117 18647 5151
rect 24409 5117 24443 5151
rect 80529 5117 80563 5151
rect 96445 5117 96479 5151
rect 97181 5117 97215 5151
rect 97825 5117 97859 5151
rect 1685 5049 1719 5083
rect 1961 5049 1995 5083
rect 3341 5049 3375 5083
rect 3525 5049 3559 5083
rect 1869 4981 1903 5015
rect 3249 4981 3283 5015
rect 24593 4981 24627 5015
rect 15209 4777 15243 4811
rect 1685 4709 1719 4743
rect 4169 4709 4203 4743
rect 4445 4709 4479 4743
rect 4905 4709 4939 4743
rect 5181 4709 5215 4743
rect 5641 4709 5675 4743
rect 5917 4709 5951 4743
rect 6377 4709 6411 4743
rect 6653 4709 6687 4743
rect 7481 4709 7515 4743
rect 11161 4709 11195 4743
rect 11345 4709 11379 4743
rect 11897 4709 11931 4743
rect 1409 4641 1443 4675
rect 2329 4641 2363 4675
rect 8125 4641 8159 4675
rect 10057 4641 10091 4675
rect 12541 4641 12575 4675
rect 13185 4641 13219 4675
rect 14933 4641 14967 4675
rect 15117 4641 15151 4675
rect 15761 4641 15795 4675
rect 16405 4641 16439 4675
rect 17233 4641 17267 4675
rect 17877 4641 17911 4675
rect 18521 4641 18555 4675
rect 19993 4641 20027 4675
rect 20637 4641 20671 4675
rect 21281 4641 21315 4675
rect 25237 4641 25271 4675
rect 25881 4641 25915 4675
rect 26525 4641 26559 4675
rect 27169 4641 27203 4675
rect 37289 4641 37323 4675
rect 39129 4641 39163 4675
rect 39773 4641 39807 4675
rect 41705 4641 41739 4675
rect 44557 4641 44591 4675
rect 46213 4641 46247 4675
rect 47041 4641 47075 4675
rect 47685 4641 47719 4675
rect 48329 4641 48363 4675
rect 52561 4641 52595 4675
rect 53205 4641 53239 4675
rect 62865 4641 62899 4675
rect 73813 4641 73847 4675
rect 78781 4641 78815 4675
rect 79425 4641 79459 4675
rect 80069 4641 80103 4675
rect 80805 4641 80839 4675
rect 81449 4641 81483 4675
rect 82921 4641 82955 4675
rect 90189 4641 90223 4675
rect 93409 4641 93443 4675
rect 94053 4641 94087 4675
rect 94697 4641 94731 4675
rect 95341 4641 95375 4675
rect 95985 4641 96019 4675
rect 96629 4641 96663 4675
rect 97273 4641 97307 4675
rect 2605 4573 2639 4607
rect 5733 4573 5767 4607
rect 6469 4573 6503 4607
rect 41981 4573 42015 4607
rect 43269 4505 43303 4539
rect 4353 4437 4387 4471
rect 5089 4437 5123 4471
rect 7573 4437 7607 4471
rect 11989 4437 12023 4471
rect 17325 4437 17359 4471
rect 65165 4437 65199 4471
rect 89729 4437 89763 4471
rect 1685 4097 1719 4131
rect 2605 4097 2639 4131
rect 11989 4097 12023 4131
rect 13553 4097 13587 4131
rect 81633 4097 81667 4131
rect 96813 4097 96847 4131
rect 96905 4097 96939 4131
rect 97457 4097 97491 4131
rect 1409 4029 1443 4063
rect 2329 4029 2363 4063
rect 4261 4029 4295 4063
rect 5181 4029 5215 4063
rect 6837 4029 6871 4063
rect 7665 4029 7699 4063
rect 8401 4029 8435 4063
rect 9045 4029 9079 4063
rect 9689 4029 9723 4063
rect 10517 4029 10551 4063
rect 12265 4029 12299 4063
rect 12909 4029 12943 4063
rect 13461 4029 13495 4063
rect 13737 4029 13771 4063
rect 14381 4029 14415 4063
rect 15025 4029 15059 4063
rect 16037 4029 16071 4063
rect 17417 4029 17451 4063
rect 18153 4029 18187 4063
rect 18889 4029 18923 4063
rect 19625 4029 19659 4063
rect 21005 4029 21039 4063
rect 22569 4029 22603 4063
rect 23213 4029 23247 4063
rect 23857 4029 23891 4063
rect 24501 4029 24535 4063
rect 25145 4029 25179 4063
rect 25881 4029 25915 4063
rect 26525 4029 26559 4063
rect 27813 4029 27847 4063
rect 28733 4029 28767 4063
rect 29377 4029 29411 4063
rect 30573 4029 30607 4063
rect 31217 4029 31251 4063
rect 31861 4029 31895 4063
rect 33609 4029 33643 4063
rect 34253 4029 34287 4063
rect 34897 4029 34931 4063
rect 35541 4029 35575 4063
rect 36185 4029 36219 4063
rect 36829 4029 36863 4063
rect 38301 4029 38335 4063
rect 38945 4029 38979 4063
rect 39957 4029 39991 4063
rect 40601 4029 40635 4063
rect 41245 4029 41279 4063
rect 41889 4029 41923 4063
rect 43545 4029 43579 4063
rect 44189 4029 44223 4063
rect 44833 4029 44867 4063
rect 46029 4029 46063 4063
rect 46673 4029 46707 4063
rect 47317 4029 47351 4063
rect 48789 4029 48823 4063
rect 49433 4029 49467 4063
rect 50077 4029 50111 4063
rect 50721 4029 50755 4063
rect 51365 4029 51399 4063
rect 52009 4029 52043 4063
rect 52653 4029 52687 4063
rect 54033 4029 54067 4063
rect 54677 4029 54711 4063
rect 55321 4029 55355 4063
rect 55965 4029 55999 4063
rect 56609 4029 56643 4063
rect 57253 4029 57287 4063
rect 57897 4029 57931 4063
rect 59277 4029 59311 4063
rect 59921 4029 59955 4063
rect 60565 4029 60599 4063
rect 61209 4029 61243 4063
rect 61853 4029 61887 4063
rect 62497 4029 62531 4063
rect 63141 4029 63175 4063
rect 64521 4029 64555 4063
rect 65165 4029 65199 4063
rect 65901 4029 65935 4063
rect 66545 4029 66579 4063
rect 67189 4029 67223 4063
rect 67833 4029 67867 4063
rect 68477 4029 68511 4063
rect 69765 4029 69799 4063
rect 70409 4029 70443 4063
rect 71053 4029 71087 4063
rect 71697 4029 71731 4063
rect 72341 4029 72375 4063
rect 72985 4029 73019 4063
rect 73629 4029 73663 4063
rect 75009 4029 75043 4063
rect 75653 4029 75687 4063
rect 76297 4029 76331 4063
rect 76941 4029 76975 4063
rect 77585 4029 77619 4063
rect 78229 4029 78263 4063
rect 78873 4029 78907 4063
rect 80253 4029 80287 4063
rect 80529 4029 80563 4063
rect 82369 4029 82403 4063
rect 83013 4029 83047 4063
rect 83657 4029 83691 4063
rect 84301 4029 84335 4063
rect 85497 4029 85531 4063
rect 86141 4029 86175 4063
rect 86785 4029 86819 4063
rect 87429 4029 87463 4063
rect 88533 4029 88567 4063
rect 89177 4029 89211 4063
rect 90741 4029 90775 4063
rect 91385 4029 91419 4063
rect 92029 4029 92063 4063
rect 92673 4029 92707 4063
rect 93317 4029 93351 4063
rect 94145 4029 94179 4063
rect 94789 4029 94823 4063
rect 95985 4029 96019 4063
rect 97181 4029 97215 4063
rect 97365 4029 97399 4063
rect 3341 3961 3375 3995
rect 4077 3961 4111 3995
rect 7849 3961 7883 3995
rect 12081 3961 12115 3995
rect 20361 3961 20395 3995
rect 97641 3961 97675 3995
rect 97917 3961 97951 3995
rect 3433 3893 3467 3927
rect 5365 3893 5399 3927
rect 7021 3893 7055 3927
rect 8493 3893 8527 3927
rect 10609 3893 10643 3927
rect 13001 3893 13035 3927
rect 14473 3893 14507 3927
rect 16129 3893 16163 3927
rect 17509 3893 17543 3927
rect 18245 3893 18279 3927
rect 18981 3893 19015 3927
rect 19717 3893 19751 3927
rect 20453 3893 20487 3927
rect 98009 3893 98043 3927
rect 2973 3689 3007 3723
rect 12081 3689 12115 3723
rect 85037 3689 85071 3723
rect 94881 3689 94915 3723
rect 2053 3621 2087 3655
rect 5365 3621 5399 3655
rect 6469 3621 6503 3655
rect 7481 3621 7515 3655
rect 8401 3621 8435 3655
rect 9781 3621 9815 3655
rect 10701 3621 10735 3655
rect 13277 3621 13311 3655
rect 15393 3621 15427 3655
rect 16497 3621 16531 3655
rect 18613 3621 18647 3655
rect 20269 3621 20303 3655
rect 21005 3621 21039 3655
rect 21741 3621 21775 3655
rect 26617 3621 26651 3655
rect 26893 3621 26927 3655
rect 31677 3621 31711 3655
rect 46765 3621 46799 3655
rect 81449 3621 81483 3655
rect 81725 3621 81759 3655
rect 95157 3621 95191 3655
rect 97365 3621 97399 3655
rect 97641 3621 97675 3655
rect 1501 3553 1535 3587
rect 2697 3553 2731 3587
rect 4813 3553 4847 3587
rect 6009 3553 6043 3587
rect 7205 3553 7239 3587
rect 8125 3553 8159 3587
rect 9505 3553 9539 3587
rect 10425 3553 10459 3587
rect 11805 3553 11839 3587
rect 12725 3553 12759 3587
rect 14841 3553 14875 3587
rect 16037 3553 16071 3587
rect 17233 3553 17267 3587
rect 18337 3553 18371 3587
rect 19993 3553 20027 3587
rect 23029 3553 23063 3587
rect 23673 3553 23707 3587
rect 25237 3553 25271 3587
rect 25881 3553 25915 3587
rect 27445 3553 27479 3587
rect 28089 3553 28123 3587
rect 28917 3553 28951 3587
rect 30481 3553 30515 3587
rect 31309 3553 31343 3587
rect 32413 3553 32447 3587
rect 33057 3553 33091 3587
rect 33701 3553 33735 3587
rect 34437 3553 34471 3587
rect 35725 3553 35759 3587
rect 36829 3553 36863 3587
rect 37473 3553 37507 3587
rect 38117 3553 38151 3587
rect 39313 3553 39347 3587
rect 40969 3553 41003 3587
rect 41705 3553 41739 3587
rect 42349 3553 42383 3587
rect 42993 3553 43027 3587
rect 43637 3553 43671 3587
rect 44833 3553 44867 3587
rect 46305 3553 46339 3587
rect 47409 3553 47443 3587
rect 48053 3553 48087 3587
rect 48697 3553 48731 3587
rect 49341 3553 49375 3587
rect 49985 3553 50019 3587
rect 51457 3553 51491 3587
rect 52101 3553 52135 3587
rect 52745 3553 52779 3587
rect 53389 3553 53423 3587
rect 54033 3553 54067 3587
rect 54677 3553 54711 3587
rect 55321 3553 55355 3587
rect 56701 3553 56735 3587
rect 57345 3553 57379 3587
rect 58173 3553 58207 3587
rect 58817 3553 58851 3587
rect 59461 3553 59495 3587
rect 60657 3553 60691 3587
rect 61945 3553 61979 3587
rect 62589 3553 62623 3587
rect 63233 3553 63267 3587
rect 63877 3553 63911 3587
rect 64521 3553 64555 3587
rect 65165 3553 65199 3587
rect 65809 3553 65843 3587
rect 67189 3553 67223 3587
rect 67925 3553 67959 3587
rect 68569 3553 68603 3587
rect 69213 3553 69247 3587
rect 69857 3553 69891 3587
rect 70501 3553 70535 3587
rect 71145 3553 71179 3587
rect 72433 3553 72467 3587
rect 73077 3553 73111 3587
rect 74089 3553 74123 3587
rect 74733 3553 74767 3587
rect 75929 3553 75963 3587
rect 76573 3553 76607 3587
rect 77677 3553 77711 3587
rect 78321 3553 78355 3587
rect 78965 3553 78999 3587
rect 79609 3553 79643 3587
rect 80253 3553 80287 3587
rect 80897 3553 80931 3587
rect 82921 3553 82955 3587
rect 83565 3553 83599 3587
rect 84393 3553 84427 3587
rect 84541 3553 84575 3587
rect 84669 3553 84703 3587
rect 84761 3553 84795 3587
rect 84945 3553 84979 3587
rect 85589 3553 85623 3587
rect 86233 3553 86267 3587
rect 86877 3553 86911 3587
rect 88165 3553 88199 3587
rect 89269 3553 89303 3587
rect 89913 3553 89947 3587
rect 90557 3553 90591 3587
rect 91201 3553 91235 3587
rect 92305 3553 92339 3587
rect 93409 3553 93443 3587
rect 94053 3553 94087 3587
rect 95709 3553 95743 3587
rect 96813 3553 96847 3587
rect 97089 3553 97123 3587
rect 17785 3485 17819 3519
rect 96629 3485 96663 3519
rect 96997 3485 97031 3519
rect 21925 3417 21959 3451
rect 26709 3417 26743 3451
rect 94973 3417 95007 3451
rect 97457 3417 97491 3451
rect 21097 3349 21131 3383
rect 22569 3349 22603 3383
rect 81633 3349 81667 3383
rect 84301 3349 84335 3383
rect 7205 3145 7239 3179
rect 25329 3145 25363 3179
rect 27721 3145 27755 3179
rect 38209 3145 38243 3179
rect 47317 3145 47351 3179
rect 55229 3145 55263 3179
rect 62497 3145 62531 3179
rect 66729 3145 66763 3179
rect 72249 3145 72283 3179
rect 80161 3145 80195 3179
rect 81909 3145 81943 3179
rect 90649 3145 90683 3179
rect 91293 3145 91327 3179
rect 93685 3145 93719 3179
rect 96629 3145 96663 3179
rect 97089 3145 97123 3179
rect 97273 3145 97307 3179
rect 15853 3077 15887 3111
rect 2421 3009 2455 3043
rect 5273 3009 5307 3043
rect 10977 3009 11011 3043
rect 12817 3009 12851 3043
rect 13737 3009 13771 3043
rect 13829 3009 13863 3043
rect 14197 3009 14231 3043
rect 15117 3009 15151 3043
rect 17693 3009 17727 3043
rect 19257 3009 19291 3043
rect 20361 3009 20395 3043
rect 21465 3009 21499 3043
rect 50629 3009 50663 3043
rect 70409 3009 70443 3043
rect 94513 3009 94547 3043
rect 2053 2941 2087 2975
rect 3157 2941 3191 2975
rect 4721 2941 4755 2975
rect 7757 2941 7791 2975
rect 8493 2941 8527 2975
rect 8861 2941 8895 2975
rect 9689 2941 9723 2975
rect 10517 2941 10551 2975
rect 13461 2941 13495 2975
rect 13644 2941 13678 2975
rect 14013 2941 14047 2975
rect 14749 2941 14783 2975
rect 17417 2941 17451 2975
rect 18889 2941 18923 2975
rect 20085 2941 20119 2975
rect 21189 2941 21223 2975
rect 22661 2941 22695 2975
rect 23305 2941 23339 2975
rect 23949 2941 23983 2975
rect 24593 2941 24627 2975
rect 25697 2941 25731 2975
rect 26341 2941 26375 2975
rect 27997 2941 28031 2975
rect 28549 2941 28583 2975
rect 29193 2941 29227 2975
rect 29837 2941 29871 2975
rect 30481 2941 30515 2975
rect 31125 2941 31159 2975
rect 31769 2941 31803 2975
rect 33057 2941 33091 2975
rect 33701 2941 33735 2975
rect 34345 2941 34379 2975
rect 35173 2941 35207 2975
rect 35449 2941 35483 2975
rect 36001 2941 36035 2975
rect 36645 2941 36679 2975
rect 38485 2941 38519 2975
rect 39037 2941 39071 2975
rect 40233 2941 40267 2975
rect 41245 2941 41279 2975
rect 41521 2941 41555 2975
rect 42073 2941 42107 2975
rect 43453 2941 43487 2975
rect 43729 2941 43763 2975
rect 44281 2941 44315 2975
rect 44925 2941 44959 2975
rect 45477 2941 45511 2975
rect 45753 2941 45787 2975
rect 46305 2941 46339 2975
rect 47593 2941 47627 2975
rect 49157 2941 49191 2975
rect 49433 2941 49467 2975
rect 50997 2941 51031 2975
rect 51273 2941 51307 2975
rect 51825 2941 51859 2975
rect 52469 2941 52503 2975
rect 54125 2941 54159 2975
rect 55505 2941 55539 2975
rect 56517 2941 56551 2975
rect 56793 2941 56827 2975
rect 57345 2941 57379 2975
rect 57989 2941 58023 2975
rect 59185 2941 59219 2975
rect 60013 2941 60047 2975
rect 60657 2941 60691 2975
rect 61393 2941 61427 2975
rect 61669 2941 61703 2975
rect 62865 2941 62899 2975
rect 63417 2941 63451 2975
rect 64429 2941 64463 2975
rect 64705 2941 64739 2975
rect 65257 2941 65291 2975
rect 65901 2941 65935 2975
rect 67097 2941 67131 2975
rect 67649 2941 67683 2975
rect 68293 2941 68327 2975
rect 69673 2941 69707 2975
rect 69949 2941 69983 2975
rect 70777 2941 70811 2975
rect 71329 2941 71363 2975
rect 72617 2941 72651 2975
rect 73169 2941 73203 2975
rect 73813 2941 73847 2975
rect 74825 2941 74859 2975
rect 75193 2941 75227 2975
rect 75745 2941 75779 2975
rect 76573 2941 76607 2975
rect 76849 2941 76883 2975
rect 77861 2941 77895 2975
rect 78137 2941 78171 2975
rect 79149 2941 79183 2975
rect 80897 2941 80931 2975
rect 81173 2941 81207 2975
rect 81817 2941 81851 2975
rect 83197 2941 83231 2975
rect 83841 2941 83875 2975
rect 85497 2941 85531 2975
rect 86141 2941 86175 2975
rect 86785 2941 86819 2975
rect 87429 2941 87463 2975
rect 88073 2941 88107 2975
rect 88717 2941 88751 2975
rect 89361 2941 89395 2975
rect 90925 2941 90959 2975
rect 91477 2941 91511 2975
rect 91661 2941 91695 2975
rect 92213 2941 92247 2975
rect 94053 2941 94087 2975
rect 94605 2941 94639 2975
rect 94789 2941 94823 2975
rect 96077 2941 96111 2975
rect 97733 2941 97767 2975
rect 3985 2873 4019 2907
rect 6929 2873 6963 2907
rect 12081 2873 12115 2907
rect 15669 2873 15703 2907
rect 16037 2873 16071 2907
rect 25513 2873 25547 2907
rect 35265 2873 35299 2907
rect 38301 2873 38335 2907
rect 41337 2873 41371 2907
rect 43545 2873 43579 2907
rect 45569 2873 45603 2907
rect 47409 2873 47443 2907
rect 49249 2873 49283 2907
rect 51089 2873 51123 2907
rect 55321 2873 55355 2907
rect 56609 2873 56643 2907
rect 59277 2873 59311 2907
rect 59461 2873 59495 2907
rect 61485 2873 61519 2907
rect 62681 2873 62715 2907
rect 64521 2873 64555 2907
rect 66913 2873 66947 2907
rect 69765 2873 69799 2907
rect 70593 2873 70627 2907
rect 72433 2873 72467 2907
rect 75009 2873 75043 2907
rect 76665 2873 76699 2907
rect 77953 2873 77987 2907
rect 80253 2873 80287 2907
rect 80437 2873 80471 2907
rect 82553 2873 82587 2907
rect 90741 2873 90775 2907
rect 93133 2873 93167 2907
rect 93317 2873 93351 2907
rect 93869 2873 93903 2907
rect 96721 2873 96755 2907
rect 96905 2873 96939 2907
rect 97273 2873 97307 2907
rect 97549 2873 97583 2907
rect 9781 2805 9815 2839
rect 22753 2805 22787 2839
rect 26433 2805 26467 2839
rect 27905 2805 27939 2839
rect 40325 2805 40359 2839
rect 54217 2805 54251 2839
rect 79241 2805 79275 2839
rect 81081 2805 81115 2839
rect 82645 2805 82679 2839
rect 92949 2805 92983 2839
rect 96169 2805 96203 2839
rect 8493 2601 8527 2635
rect 13461 2601 13495 2635
rect 22753 2601 22787 2635
rect 26893 2601 26927 2635
rect 28181 2601 28215 2635
rect 28641 2601 28675 2635
rect 28825 2601 28859 2635
rect 29653 2601 29687 2635
rect 30757 2601 30791 2635
rect 31493 2601 31527 2635
rect 32045 2601 32079 2635
rect 34161 2601 34195 2635
rect 36185 2601 36219 2635
rect 36645 2601 36679 2635
rect 36921 2601 36955 2635
rect 38853 2601 38887 2635
rect 39405 2601 39439 2635
rect 40233 2601 40267 2635
rect 41429 2601 41463 2635
rect 48605 2601 48639 2635
rect 49433 2601 49467 2635
rect 50905 2601 50939 2635
rect 54769 2601 54803 2635
rect 58173 2601 58207 2635
rect 60197 2601 60231 2635
rect 61669 2601 61703 2635
rect 65717 2601 65751 2635
rect 66269 2601 66303 2635
rect 68845 2601 68879 2635
rect 69581 2601 69615 2635
rect 70133 2601 70167 2635
rect 70777 2601 70811 2635
rect 71513 2601 71547 2635
rect 74181 2601 74215 2635
rect 74917 2601 74951 2635
rect 77585 2601 77619 2635
rect 78873 2601 78907 2635
rect 79517 2601 79551 2635
rect 81541 2601 81575 2635
rect 82093 2601 82127 2635
rect 84761 2601 84795 2635
rect 84853 2601 84887 2635
rect 88349 2601 88383 2635
rect 89453 2601 89487 2635
rect 90005 2601 90039 2635
rect 90741 2601 90775 2635
rect 92121 2601 92155 2635
rect 92857 2601 92891 2635
rect 94789 2601 94823 2635
rect 95525 2601 95559 2635
rect 96261 2601 96295 2635
rect 2237 2533 2271 2567
rect 3157 2533 3191 2567
rect 4997 2533 5031 2567
rect 7665 2533 7699 2567
rect 10425 2533 10459 2567
rect 11161 2533 11195 2567
rect 12265 2533 12299 2567
rect 13093 2533 13127 2567
rect 13829 2533 13863 2567
rect 15577 2533 15611 2567
rect 16681 2533 16715 2567
rect 18429 2533 18463 2567
rect 18981 2533 19015 2567
rect 19257 2533 19291 2567
rect 20361 2533 20395 2567
rect 21833 2533 21867 2567
rect 23121 2533 23155 2567
rect 23581 2533 23615 2567
rect 23857 2533 23891 2567
rect 24501 2533 24535 2567
rect 25513 2533 25547 2567
rect 25789 2533 25823 2567
rect 27261 2533 27295 2567
rect 28457 2533 28491 2567
rect 29193 2533 29227 2567
rect 29929 2533 29963 2567
rect 31125 2533 31159 2567
rect 31861 2533 31895 2567
rect 32321 2533 32355 2567
rect 32597 2533 32631 2567
rect 33701 2533 33735 2567
rect 34529 2533 34563 2567
rect 35173 2533 35207 2567
rect 36461 2533 36495 2567
rect 37197 2533 37231 2567
rect 37657 2533 37691 2567
rect 37933 2533 37967 2567
rect 38945 2533 38979 2567
rect 39129 2533 39163 2567
rect 39589 2533 39623 2567
rect 39865 2533 39899 2567
rect 40601 2533 40635 2567
rect 42441 2533 42475 2567
rect 42993 2533 43027 2567
rect 43269 2533 43303 2567
rect 44189 2533 44223 2567
rect 44465 2533 44499 2567
rect 45109 2533 45143 2567
rect 45661 2533 45695 2567
rect 45937 2533 45971 2567
rect 46121 2533 46155 2567
rect 47041 2533 47075 2567
rect 48513 2533 48547 2567
rect 49801 2533 49835 2567
rect 50261 2533 50295 2567
rect 50537 2533 50571 2567
rect 51273 2533 51307 2567
rect 52377 2533 52411 2567
rect 52929 2533 52963 2567
rect 53205 2533 53239 2567
rect 53849 2533 53883 2567
rect 55137 2533 55171 2567
rect 55781 2533 55815 2567
rect 56333 2533 56367 2567
rect 56609 2533 56643 2567
rect 57529 2533 57563 2567
rect 57805 2533 57839 2567
rect 58357 2533 58391 2567
rect 58541 2533 58575 2567
rect 59001 2533 59035 2567
rect 59277 2533 59311 2567
rect 60473 2533 60507 2567
rect 60933 2533 60967 2567
rect 61209 2533 61243 2567
rect 61761 2533 61795 2567
rect 61945 2533 61979 2567
rect 62865 2533 62899 2567
rect 63141 2533 63175 2567
rect 63325 2533 63359 2567
rect 63601 2533 63635 2567
rect 63877 2533 63911 2567
rect 65533 2533 65567 2567
rect 65809 2533 65843 2567
rect 66545 2533 66579 2567
rect 67189 2533 67223 2567
rect 68385 2533 68419 2567
rect 69213 2533 69247 2567
rect 69949 2533 69983 2567
rect 71145 2533 71179 2567
rect 71881 2533 71915 2567
rect 72341 2533 72375 2567
rect 72617 2533 72651 2567
rect 72801 2533 72835 2567
rect 74365 2533 74399 2567
rect 74549 2533 74583 2567
rect 75285 2533 75319 2567
rect 76205 2533 76239 2567
rect 76481 2533 76515 2567
rect 76941 2533 76975 2567
rect 77217 2533 77251 2567
rect 77953 2533 77987 2567
rect 79149 2533 79183 2567
rect 79885 2533 79919 2567
rect 80529 2533 80563 2567
rect 81817 2533 81851 2567
rect 82921 2533 82955 2567
rect 84393 2533 84427 2567
rect 85681 2533 85715 2567
rect 85957 2533 85991 2567
rect 87061 2533 87095 2567
rect 87613 2533 87647 2567
rect 87889 2533 87923 2567
rect 88625 2533 88659 2567
rect 89637 2533 89671 2567
rect 89821 2533 89855 2567
rect 90281 2533 90315 2567
rect 90557 2533 90591 2567
rect 91201 2533 91235 2567
rect 92489 2533 92523 2567
rect 93225 2533 93259 2567
rect 93685 2533 93719 2567
rect 93961 2533 93995 2567
rect 95157 2533 95191 2567
rect 95893 2533 95927 2567
rect 96537 2533 96571 2567
rect 96721 2533 96755 2567
rect 1409 2465 1443 2499
rect 2881 2465 2915 2499
rect 4261 2465 4295 2499
rect 5641 2465 5675 2499
rect 6929 2465 6963 2499
rect 8309 2465 8343 2499
rect 9689 2465 9723 2499
rect 15025 2465 15059 2499
rect 16313 2465 16347 2499
rect 17601 2465 17635 2499
rect 21189 2465 21223 2499
rect 26249 2465 26283 2499
rect 26525 2465 26559 2499
rect 36277 2465 36311 2499
rect 40417 2465 40451 2499
rect 41797 2465 41831 2499
rect 44281 2465 44315 2499
rect 47777 2465 47811 2499
rect 53021 2465 53055 2499
rect 57621 2465 57655 2499
rect 60289 2465 60323 2499
rect 64521 2465 64555 2499
rect 69765 2465 69799 2499
rect 73721 2465 73755 2499
rect 77769 2465 77803 2499
rect 79701 2465 79735 2499
rect 84761 2465 84795 2499
rect 85221 2465 85255 2499
rect 97641 2465 97675 2499
rect 97917 2465 97951 2499
rect 19073 2397 19107 2431
rect 25605 2397 25639 2431
rect 26341 2397 26375 2431
rect 31677 2397 31711 2431
rect 34345 2397 34379 2431
rect 37749 2397 37783 2431
rect 41613 2397 41647 2431
rect 43085 2397 43119 2431
rect 47225 2397 47259 2431
rect 51089 2397 51123 2431
rect 54953 2397 54987 2431
rect 55965 2397 55999 2431
rect 62957 2397 62991 2431
rect 63693 2397 63727 2431
rect 67373 2397 67407 2431
rect 70961 2397 70995 2431
rect 72433 2397 72467 2431
rect 76297 2397 76331 2431
rect 80713 2397 80747 2431
rect 85773 2397 85807 2431
rect 88441 2397 88475 2431
rect 90373 2397 90407 2431
rect 91385 2397 91419 2431
rect 94973 2397 95007 2431
rect 5825 2329 5859 2363
rect 13645 2329 13679 2363
rect 20545 2329 20579 2363
rect 22937 2329 22971 2363
rect 24685 2329 24719 2363
rect 27077 2329 27111 2363
rect 28273 2329 28307 2363
rect 29009 2329 29043 2363
rect 29745 2329 29779 2363
rect 30941 2329 30975 2363
rect 32413 2329 32447 2363
rect 37013 2329 37047 2363
rect 42625 2329 42659 2363
rect 45753 2329 45787 2363
rect 49617 2329 49651 2363
rect 56425 2329 56459 2363
rect 61025 2329 61059 2363
rect 66361 2329 66395 2363
rect 69029 2329 69063 2363
rect 71697 2329 71731 2363
rect 75101 2329 75135 2363
rect 81633 2329 81667 2363
rect 85037 2329 85071 2363
rect 87705 2329 87739 2363
rect 92305 2329 92339 2363
rect 93041 2329 93075 2363
rect 93777 2329 93811 2363
rect 95709 2329 95743 2363
rect 98101 2329 98135 2363
rect 11253 2261 11287 2295
rect 23765 2261 23799 2295
rect 33793 2261 33827 2295
rect 35265 2261 35299 2295
rect 39773 2261 39807 2295
rect 45201 2261 45235 2295
rect 47869 2261 47903 2295
rect 50445 2261 50479 2295
rect 52469 2261 52503 2295
rect 53941 2261 53975 2295
rect 59185 2261 59219 2295
rect 64613 2261 64647 2295
rect 68477 2261 68511 2295
rect 73813 2261 73847 2295
rect 77125 2261 77159 2295
rect 79057 2261 79091 2295
rect 83013 2261 83047 2295
rect 84485 2261 84519 2295
rect 87153 2261 87187 2295
<< metal1 >>
rect 16298 97588 16304 97640
rect 16356 97628 16362 97640
rect 90450 97628 90456 97640
rect 16356 97600 90456 97628
rect 16356 97588 16362 97600
rect 90450 97588 90456 97600
rect 90508 97588 90514 97640
rect 23934 97520 23940 97572
rect 23992 97560 23998 97572
rect 56502 97560 56508 97572
rect 23992 97532 56508 97560
rect 23992 97520 23998 97532
rect 56502 97520 56508 97532
rect 56560 97520 56566 97572
rect 7650 97452 7656 97504
rect 7708 97492 7714 97504
rect 68554 97492 68560 97504
rect 7708 97464 68560 97492
rect 7708 97452 7714 97464
rect 68554 97452 68560 97464
rect 68612 97452 68618 97504
rect 1104 97402 98808 97424
rect 1104 97350 19606 97402
rect 19658 97350 19670 97402
rect 19722 97350 19734 97402
rect 19786 97350 19798 97402
rect 19850 97350 50326 97402
rect 50378 97350 50390 97402
rect 50442 97350 50454 97402
rect 50506 97350 50518 97402
rect 50570 97350 81046 97402
rect 81098 97350 81110 97402
rect 81162 97350 81174 97402
rect 81226 97350 81238 97402
rect 81290 97350 98808 97402
rect 1104 97328 98808 97350
rect 1210 97248 1216 97300
rect 1268 97288 1274 97300
rect 2317 97291 2375 97297
rect 2317 97288 2329 97291
rect 1268 97260 2329 97288
rect 1268 97248 1274 97260
rect 2317 97257 2329 97260
rect 2363 97257 2375 97291
rect 2317 97251 2375 97257
rect 3786 97248 3792 97300
rect 3844 97288 3850 97300
rect 4433 97291 4491 97297
rect 4433 97288 4445 97291
rect 3844 97260 4445 97288
rect 3844 97248 3850 97260
rect 4433 97257 4445 97260
rect 4479 97257 4491 97291
rect 4433 97251 4491 97257
rect 6454 97248 6460 97300
rect 6512 97288 6518 97300
rect 7101 97291 7159 97297
rect 7101 97288 7113 97291
rect 6512 97260 7113 97288
rect 6512 97248 6518 97260
rect 7101 97257 7113 97260
rect 7147 97257 7159 97291
rect 7101 97251 7159 97257
rect 9030 97248 9036 97300
rect 9088 97288 9094 97300
rect 9769 97291 9827 97297
rect 9769 97288 9781 97291
rect 9088 97260 9781 97288
rect 9088 97248 9094 97260
rect 9769 97257 9781 97260
rect 9815 97257 9827 97291
rect 9769 97251 9827 97257
rect 11606 97248 11612 97300
rect 11664 97288 11670 97300
rect 12437 97291 12495 97297
rect 12437 97288 12449 97291
rect 11664 97260 12449 97288
rect 11664 97248 11670 97260
rect 12437 97257 12449 97260
rect 12483 97257 12495 97291
rect 12437 97251 12495 97257
rect 14200 97260 16574 97288
rect 2958 97220 2964 97232
rect 2919 97192 2964 97220
rect 2958 97180 2964 97192
rect 3016 97180 3022 97232
rect 4341 97223 4399 97229
rect 4341 97189 4353 97223
rect 4387 97220 4399 97223
rect 6178 97220 6184 97232
rect 4387 97192 6184 97220
rect 4387 97189 4399 97192
rect 4341 97183 4399 97189
rect 6178 97180 6184 97192
rect 6236 97180 6242 97232
rect 10778 97180 10784 97232
rect 10836 97220 10842 97232
rect 10873 97223 10931 97229
rect 10873 97220 10885 97223
rect 10836 97192 10885 97220
rect 10836 97180 10842 97192
rect 10873 97189 10885 97192
rect 10919 97189 10931 97223
rect 14200 97220 14228 97260
rect 10873 97183 10931 97189
rect 12176 97192 14228 97220
rect 382 97112 388 97164
rect 440 97152 446 97164
rect 1397 97155 1455 97161
rect 1397 97152 1409 97155
rect 440 97124 1409 97152
rect 440 97112 446 97124
rect 1397 97121 1409 97124
rect 1443 97121 1455 97155
rect 1397 97115 1455 97121
rect 2225 97155 2283 97161
rect 2225 97121 2237 97155
rect 2271 97152 2283 97155
rect 2498 97152 2504 97164
rect 2271 97124 2504 97152
rect 2271 97121 2283 97124
rect 2225 97115 2283 97121
rect 2498 97112 2504 97124
rect 2556 97112 2562 97164
rect 5534 97152 5540 97164
rect 5495 97124 5540 97152
rect 5534 97112 5540 97124
rect 5592 97112 5598 97164
rect 7006 97152 7012 97164
rect 6967 97124 7012 97152
rect 7006 97112 7012 97124
rect 7064 97112 7070 97164
rect 8202 97152 8208 97164
rect 8163 97124 8208 97152
rect 8202 97112 8208 97124
rect 8260 97112 8266 97164
rect 9677 97155 9735 97161
rect 9677 97121 9689 97155
rect 9723 97152 9735 97155
rect 12176 97152 12204 97192
rect 14274 97180 14280 97232
rect 14332 97220 14338 97232
rect 15197 97223 15255 97229
rect 15197 97220 15209 97223
rect 14332 97192 15209 97220
rect 14332 97180 14338 97192
rect 15197 97189 15209 97192
rect 15243 97189 15255 97223
rect 15197 97183 15255 97189
rect 16022 97180 16028 97232
rect 16080 97220 16086 97232
rect 16117 97223 16175 97229
rect 16117 97220 16129 97223
rect 16080 97192 16129 97220
rect 16080 97180 16086 97192
rect 16117 97189 16129 97192
rect 16163 97189 16175 97223
rect 16546 97220 16574 97260
rect 16850 97248 16856 97300
rect 16908 97288 16914 97300
rect 17773 97291 17831 97297
rect 17773 97288 17785 97291
rect 16908 97260 17785 97288
rect 16908 97248 16914 97260
rect 17773 97257 17785 97260
rect 17819 97257 17831 97291
rect 17773 97251 17831 97257
rect 19426 97248 19432 97300
rect 19484 97288 19490 97300
rect 20441 97291 20499 97297
rect 20441 97288 20453 97291
rect 19484 97260 20453 97288
rect 19484 97248 19490 97260
rect 20441 97257 20453 97260
rect 20487 97257 20499 97291
rect 20441 97251 20499 97257
rect 22094 97248 22100 97300
rect 22152 97288 22158 97300
rect 23109 97291 23167 97297
rect 23109 97288 23121 97291
rect 22152 97260 23121 97288
rect 22152 97248 22158 97260
rect 23109 97257 23121 97260
rect 23155 97257 23167 97291
rect 23109 97251 23167 97257
rect 23216 97260 26648 97288
rect 16546 97192 17816 97220
rect 16117 97183 16175 97189
rect 12342 97152 12348 97164
rect 9723 97124 12204 97152
rect 12303 97124 12348 97152
rect 9723 97121 9735 97124
rect 9677 97115 9735 97121
rect 12342 97112 12348 97124
rect 12400 97112 12406 97164
rect 13354 97152 13360 97164
rect 13315 97124 13360 97152
rect 13354 97112 13360 97124
rect 13412 97112 13418 97164
rect 15010 97152 15016 97164
rect 14971 97124 15016 97152
rect 15010 97112 15016 97124
rect 15068 97112 15074 97164
rect 17678 97152 17684 97164
rect 17639 97124 17684 97152
rect 17678 97112 17684 97124
rect 17736 97112 17742 97164
rect 17788 97152 17816 97192
rect 18598 97180 18604 97232
rect 18656 97220 18662 97232
rect 18693 97223 18751 97229
rect 18693 97220 18705 97223
rect 18656 97192 18705 97220
rect 18656 97180 18662 97192
rect 18693 97189 18705 97192
rect 18739 97189 18751 97223
rect 21450 97220 21456 97232
rect 18693 97183 18751 97189
rect 18800 97192 21456 97220
rect 18800 97152 18828 97192
rect 21450 97180 21456 97192
rect 21508 97180 21514 97232
rect 22830 97180 22836 97232
rect 22888 97220 22894 97232
rect 23216 97220 23244 97260
rect 22888 97192 23244 97220
rect 23569 97223 23627 97229
rect 22888 97180 22894 97192
rect 23569 97189 23581 97223
rect 23615 97220 23627 97223
rect 23845 97223 23903 97229
rect 23845 97220 23857 97223
rect 23615 97192 23857 97220
rect 23615 97189 23627 97192
rect 23569 97183 23627 97189
rect 23845 97189 23857 97192
rect 23891 97220 23903 97223
rect 23934 97220 23940 97232
rect 23891 97192 23940 97220
rect 23891 97189 23903 97192
rect 23845 97183 23903 97189
rect 23934 97180 23940 97192
rect 23992 97180 23998 97232
rect 24670 97220 24676 97232
rect 24631 97192 24676 97220
rect 24670 97180 24676 97192
rect 24728 97180 24734 97232
rect 26418 97180 26424 97232
rect 26476 97220 26482 97232
rect 26513 97223 26571 97229
rect 26513 97220 26525 97223
rect 26476 97192 26525 97220
rect 26476 97180 26482 97192
rect 26513 97189 26525 97192
rect 26559 97189 26571 97223
rect 26620 97220 26648 97260
rect 27338 97248 27344 97300
rect 27396 97288 27402 97300
rect 28445 97291 28503 97297
rect 28445 97288 28457 97291
rect 27396 97260 28457 97288
rect 27396 97248 27402 97260
rect 28445 97257 28457 97260
rect 28491 97257 28503 97291
rect 29914 97288 29920 97300
rect 29875 97260 29920 97288
rect 28445 97251 28503 97257
rect 29914 97248 29920 97260
rect 29972 97248 29978 97300
rect 30742 97248 30748 97300
rect 30800 97288 30806 97300
rect 31113 97291 31171 97297
rect 31113 97288 31125 97291
rect 30800 97260 31125 97288
rect 30800 97248 30806 97260
rect 31113 97257 31125 97260
rect 31159 97257 31171 97291
rect 31113 97251 31171 97257
rect 32490 97248 32496 97300
rect 32548 97288 32554 97300
rect 32585 97291 32643 97297
rect 32585 97288 32597 97291
rect 32548 97260 32597 97288
rect 32548 97248 32554 97260
rect 32585 97257 32597 97260
rect 32631 97257 32643 97291
rect 32585 97251 32643 97257
rect 34425 97291 34483 97297
rect 34425 97257 34437 97291
rect 34471 97257 34483 97291
rect 34425 97251 34483 97257
rect 26620 97192 28488 97220
rect 26513 97183 26571 97189
rect 20346 97152 20352 97164
rect 17788 97124 18828 97152
rect 20307 97124 20352 97152
rect 20346 97112 20352 97124
rect 20404 97112 20410 97164
rect 21174 97152 21180 97164
rect 21135 97124 21180 97152
rect 21174 97112 21180 97124
rect 21232 97112 21238 97164
rect 23017 97155 23075 97161
rect 23017 97121 23029 97155
rect 23063 97152 23075 97155
rect 23106 97152 23112 97164
rect 23063 97124 23112 97152
rect 23063 97121 23075 97124
rect 23017 97115 23075 97121
rect 23106 97112 23112 97124
rect 23164 97112 23170 97164
rect 24486 97152 24492 97164
rect 24447 97124 24492 97152
rect 24486 97112 24492 97124
rect 24544 97112 24550 97164
rect 25777 97155 25835 97161
rect 25777 97121 25789 97155
rect 25823 97152 25835 97155
rect 26050 97152 26056 97164
rect 25823 97124 26056 97152
rect 25823 97121 25835 97124
rect 25777 97115 25835 97121
rect 26050 97112 26056 97124
rect 26108 97112 26114 97164
rect 28258 97112 28264 97164
rect 28316 97152 28322 97164
rect 28353 97155 28411 97161
rect 28353 97152 28365 97155
rect 28316 97124 28365 97152
rect 28316 97112 28322 97124
rect 28353 97121 28365 97124
rect 28399 97121 28411 97155
rect 28353 97115 28411 97121
rect 5718 97084 5724 97096
rect 5679 97056 5724 97084
rect 5718 97044 5724 97056
rect 5776 97044 5782 97096
rect 8481 97087 8539 97093
rect 8481 97053 8493 97087
rect 8527 97084 8539 97087
rect 8754 97084 8760 97096
rect 8527 97056 8760 97084
rect 8527 97053 8539 97056
rect 8481 97047 8539 97053
rect 8754 97044 8760 97056
rect 8812 97044 8818 97096
rect 13633 97087 13691 97093
rect 13633 97053 13645 97087
rect 13679 97084 13691 97087
rect 14826 97084 14832 97096
rect 13679 97056 14832 97084
rect 13679 97053 13691 97056
rect 13633 97047 13691 97053
rect 14826 97044 14832 97056
rect 14884 97044 14890 97096
rect 21358 97084 21364 97096
rect 21319 97056 21364 97084
rect 21358 97044 21364 97056
rect 21416 97044 21422 97096
rect 25961 97087 26019 97093
rect 25961 97053 25973 97087
rect 26007 97084 26019 97087
rect 28166 97084 28172 97096
rect 26007 97056 28172 97084
rect 26007 97053 26019 97056
rect 25961 97047 26019 97053
rect 28166 97044 28172 97056
rect 28224 97044 28230 97096
rect 28460 97084 28488 97192
rect 28994 97180 29000 97232
rect 29052 97220 29058 97232
rect 29089 97223 29147 97229
rect 29089 97220 29101 97223
rect 29052 97192 29101 97220
rect 29052 97180 29058 97192
rect 29089 97189 29101 97192
rect 29135 97189 29147 97223
rect 31754 97220 31760 97232
rect 31715 97192 31760 97220
rect 29089 97183 29147 97189
rect 31754 97180 31760 97192
rect 31812 97180 31818 97232
rect 29822 97152 29828 97164
rect 29783 97124 29828 97152
rect 29822 97112 29828 97124
rect 29880 97112 29886 97164
rect 31018 97152 31024 97164
rect 30979 97124 31024 97152
rect 31018 97112 31024 97124
rect 31076 97112 31082 97164
rect 32490 97152 32496 97164
rect 32451 97124 32496 97152
rect 32490 97112 32496 97124
rect 32548 97112 32554 97164
rect 34238 97152 34244 97164
rect 34199 97124 34244 97152
rect 34238 97112 34244 97124
rect 34296 97112 34302 97164
rect 34440 97084 34468 97251
rect 35158 97248 35164 97300
rect 35216 97288 35222 97300
rect 35253 97291 35311 97297
rect 35253 97288 35265 97291
rect 35216 97260 35265 97288
rect 35216 97248 35222 97260
rect 35253 97257 35265 97260
rect 35299 97257 35311 97291
rect 35253 97251 35311 97257
rect 37734 97248 37740 97300
rect 37792 97288 37798 97300
rect 37921 97291 37979 97297
rect 37921 97288 37933 97291
rect 37792 97260 37933 97288
rect 37792 97248 37798 97260
rect 37921 97257 37933 97260
rect 37967 97257 37979 97291
rect 37921 97251 37979 97257
rect 40310 97248 40316 97300
rect 40368 97288 40374 97300
rect 40589 97291 40647 97297
rect 40589 97288 40601 97291
rect 40368 97260 40601 97288
rect 40368 97248 40374 97260
rect 40589 97257 40601 97260
rect 40635 97257 40647 97291
rect 40589 97251 40647 97257
rect 42978 97248 42984 97300
rect 43036 97288 43042 97300
rect 43165 97291 43223 97297
rect 43165 97288 43177 97291
rect 43036 97260 43177 97288
rect 43036 97248 43042 97260
rect 43165 97257 43177 97260
rect 43211 97257 43223 97291
rect 90450 97288 90456 97300
rect 43165 97251 43223 97257
rect 43548 97260 44956 97288
rect 36814 97180 36820 97232
rect 36872 97220 36878 97232
rect 36909 97223 36967 97229
rect 36909 97220 36921 97223
rect 36872 97192 36921 97220
rect 36872 97180 36878 97192
rect 36909 97189 36921 97192
rect 36955 97189 36967 97223
rect 36909 97183 36967 97189
rect 39482 97180 39488 97232
rect 39540 97220 39546 97232
rect 39577 97223 39635 97229
rect 39577 97220 39589 97223
rect 39540 97192 39589 97220
rect 39540 97180 39546 97192
rect 39577 97189 39589 97192
rect 39623 97189 39635 97223
rect 39577 97183 39635 97189
rect 42058 97180 42064 97232
rect 42116 97220 42122 97232
rect 42153 97223 42211 97229
rect 42153 97220 42165 97223
rect 42116 97192 42165 97220
rect 42116 97180 42122 97192
rect 42153 97189 42165 97192
rect 42199 97189 42211 97223
rect 42153 97183 42211 97189
rect 34790 97112 34796 97164
rect 34848 97152 34854 97164
rect 35161 97155 35219 97161
rect 35161 97152 35173 97155
rect 34848 97124 35173 97152
rect 34848 97112 34854 97124
rect 35161 97121 35173 97124
rect 35207 97121 35219 97155
rect 37826 97152 37832 97164
rect 37787 97124 37832 97152
rect 35161 97115 35219 97121
rect 37826 97112 37832 97124
rect 37884 97112 37890 97164
rect 40494 97152 40500 97164
rect 40455 97124 40500 97152
rect 40494 97112 40500 97124
rect 40552 97112 40558 97164
rect 43070 97152 43076 97164
rect 43031 97124 43076 97152
rect 43070 97112 43076 97124
rect 43128 97112 43134 97164
rect 43548 97152 43576 97260
rect 44726 97180 44732 97232
rect 44784 97220 44790 97232
rect 44821 97223 44879 97229
rect 44821 97220 44833 97223
rect 44784 97192 44833 97220
rect 44784 97180 44790 97192
rect 44821 97189 44833 97192
rect 44867 97189 44879 97223
rect 44928 97220 44956 97260
rect 45526 97260 90312 97288
rect 90411 97260 90456 97288
rect 45526 97220 45554 97260
rect 44928 97192 45554 97220
rect 44821 97183 44879 97189
rect 47302 97180 47308 97232
rect 47360 97220 47366 97232
rect 47397 97223 47455 97229
rect 47397 97220 47409 97223
rect 47360 97192 47409 97220
rect 47360 97180 47366 97192
rect 47397 97189 47409 97192
rect 47443 97189 47455 97223
rect 47397 97183 47455 97189
rect 48130 97180 48136 97232
rect 48188 97220 48194 97232
rect 48501 97223 48559 97229
rect 48501 97220 48513 97223
rect 48188 97192 48513 97220
rect 48188 97180 48194 97192
rect 48501 97189 48513 97192
rect 48547 97189 48559 97223
rect 48501 97183 48559 97189
rect 50798 97180 50804 97232
rect 50856 97220 50862 97232
rect 51077 97223 51135 97229
rect 51077 97220 51089 97223
rect 50856 97192 51089 97220
rect 50856 97180 50862 97192
rect 51077 97189 51089 97192
rect 51123 97189 51135 97223
rect 51077 97183 51135 97189
rect 53374 97180 53380 97232
rect 53432 97220 53438 97232
rect 53653 97223 53711 97229
rect 53653 97220 53665 97223
rect 53432 97192 53665 97220
rect 53432 97180 53438 97192
rect 53653 97189 53665 97192
rect 53699 97189 53711 97223
rect 53653 97183 53711 97189
rect 55950 97180 55956 97232
rect 56008 97220 56014 97232
rect 56321 97223 56379 97229
rect 56321 97220 56333 97223
rect 56008 97192 56333 97220
rect 56008 97180 56014 97192
rect 56321 97189 56333 97192
rect 56367 97189 56379 97223
rect 56321 97183 56379 97189
rect 57698 97180 57704 97232
rect 57756 97220 57762 97232
rect 57793 97223 57851 97229
rect 57793 97220 57805 97223
rect 57756 97192 57805 97220
rect 57756 97180 57762 97192
rect 57793 97189 57805 97192
rect 57839 97189 57851 97223
rect 57793 97183 57851 97189
rect 58618 97180 58624 97232
rect 58676 97220 58682 97232
rect 58897 97223 58955 97229
rect 58897 97220 58909 97223
rect 58676 97192 58909 97220
rect 58676 97180 58682 97192
rect 58897 97189 58909 97192
rect 58943 97189 58955 97223
rect 58897 97183 58955 97189
rect 60366 97180 60372 97232
rect 60424 97220 60430 97232
rect 60461 97223 60519 97229
rect 60461 97220 60473 97223
rect 60424 97192 60473 97220
rect 60424 97180 60430 97192
rect 60461 97189 60473 97192
rect 60507 97189 60519 97223
rect 60461 97183 60519 97189
rect 61194 97180 61200 97232
rect 61252 97220 61258 97232
rect 61565 97223 61623 97229
rect 61565 97220 61577 97223
rect 61252 97192 61577 97220
rect 61252 97180 61258 97192
rect 61565 97189 61577 97192
rect 61611 97189 61623 97223
rect 61565 97183 61623 97189
rect 63862 97180 63868 97232
rect 63920 97220 63926 97232
rect 64141 97223 64199 97229
rect 64141 97220 64153 97223
rect 63920 97192 64153 97220
rect 63920 97180 63926 97192
rect 64141 97189 64153 97192
rect 64187 97189 64199 97223
rect 64141 97183 64199 97189
rect 65518 97180 65524 97232
rect 65576 97220 65582 97232
rect 65705 97223 65763 97229
rect 65705 97220 65717 97223
rect 65576 97192 65717 97220
rect 65576 97180 65582 97192
rect 65705 97189 65717 97192
rect 65751 97189 65763 97223
rect 65705 97183 65763 97189
rect 66438 97180 66444 97232
rect 66496 97220 66502 97232
rect 66717 97223 66775 97229
rect 66717 97220 66729 97223
rect 66496 97192 66729 97220
rect 66496 97180 66502 97192
rect 66717 97189 66729 97192
rect 66763 97189 66775 97223
rect 68554 97220 68560 97232
rect 68515 97192 68560 97220
rect 66717 97183 66775 97189
rect 68554 97180 68560 97192
rect 68612 97180 68618 97232
rect 69014 97180 69020 97232
rect 69072 97220 69078 97232
rect 69477 97223 69535 97229
rect 69477 97220 69489 97223
rect 69072 97192 69489 97220
rect 69072 97180 69078 97192
rect 69477 97189 69489 97192
rect 69523 97189 69535 97223
rect 69477 97183 69535 97189
rect 69934 97180 69940 97232
rect 69992 97220 69998 97232
rect 72697 97223 72755 97229
rect 72697 97220 72709 97223
rect 69992 97192 72709 97220
rect 69992 97180 69998 97192
rect 72697 97189 72709 97192
rect 72743 97189 72755 97223
rect 72697 97183 72755 97189
rect 74258 97180 74264 97232
rect 74316 97220 74322 97232
rect 74629 97223 74687 97229
rect 74629 97220 74641 97223
rect 74316 97192 74641 97220
rect 74316 97180 74322 97192
rect 74629 97189 74641 97192
rect 74675 97189 74687 97223
rect 74629 97183 74687 97189
rect 76006 97180 76012 97232
rect 76064 97220 76070 97232
rect 76377 97223 76435 97229
rect 76377 97220 76389 97223
rect 76064 97192 76389 97220
rect 76064 97180 76070 97192
rect 76377 97189 76389 97192
rect 76423 97189 76435 97223
rect 76377 97183 76435 97189
rect 76834 97180 76840 97232
rect 76892 97220 76898 97232
rect 77481 97223 77539 97229
rect 77481 97220 77493 97223
rect 76892 97192 77493 97220
rect 76892 97180 76898 97192
rect 77481 97189 77493 97192
rect 77527 97189 77539 97223
rect 77481 97183 77539 97189
rect 79502 97180 79508 97232
rect 79560 97220 79566 97232
rect 80149 97223 80207 97229
rect 80149 97220 80161 97223
rect 79560 97192 80161 97220
rect 79560 97180 79566 97192
rect 80149 97189 80161 97192
rect 80195 97189 80207 97223
rect 80149 97183 80207 97189
rect 82078 97180 82084 97232
rect 82136 97220 82142 97232
rect 82357 97223 82415 97229
rect 82357 97220 82369 97223
rect 82136 97192 82369 97220
rect 82136 97180 82142 97192
rect 82357 97189 82369 97192
rect 82403 97189 82415 97223
rect 84654 97220 84660 97232
rect 84615 97192 84660 97220
rect 82357 97183 82415 97189
rect 84654 97180 84660 97192
rect 84712 97180 84718 97232
rect 87322 97220 87328 97232
rect 87283 97192 87328 97220
rect 87322 97180 87328 97192
rect 87380 97180 87386 97232
rect 89898 97220 89904 97232
rect 89859 97192 89904 97220
rect 89898 97180 89904 97192
rect 89956 97180 89962 97232
rect 43364 97124 43576 97152
rect 28460 97056 34468 97084
rect 42058 97044 42064 97096
rect 42116 97084 42122 97096
rect 43364 97084 43392 97124
rect 45462 97112 45468 97164
rect 45520 97152 45526 97164
rect 45649 97155 45707 97161
rect 45649 97152 45661 97155
rect 45520 97124 45661 97152
rect 45520 97112 45526 97124
rect 45649 97121 45661 97124
rect 45695 97121 45707 97155
rect 48314 97152 48320 97164
rect 48275 97124 48320 97152
rect 45649 97115 45707 97121
rect 48314 97112 48320 97124
rect 48372 97112 48378 97164
rect 49878 97152 49884 97164
rect 49839 97124 49884 97152
rect 49878 97112 49884 97124
rect 49936 97112 49942 97164
rect 50890 97152 50896 97164
rect 50851 97124 50896 97152
rect 50890 97112 50896 97124
rect 50948 97112 50954 97164
rect 52546 97152 52552 97164
rect 52507 97124 52552 97152
rect 52546 97112 52552 97124
rect 52604 97112 52610 97164
rect 53466 97152 53472 97164
rect 53427 97124 53472 97152
rect 53466 97112 53472 97124
rect 53524 97112 53530 97164
rect 55122 97152 55128 97164
rect 55083 97124 55128 97152
rect 55122 97112 55128 97124
rect 55180 97112 55186 97164
rect 56137 97155 56195 97161
rect 56137 97121 56149 97155
rect 56183 97121 56195 97155
rect 56137 97115 56195 97121
rect 42116 97056 43392 97084
rect 42116 97044 42122 97056
rect 43438 97044 43444 97096
rect 43496 97084 43502 97096
rect 50065 97087 50123 97093
rect 50065 97084 50077 97087
rect 43496 97056 50077 97084
rect 43496 97044 43502 97056
rect 50065 97053 50077 97056
rect 50111 97053 50123 97087
rect 55309 97087 55367 97093
rect 55309 97084 55321 97087
rect 50065 97047 50123 97053
rect 55186 97056 55321 97084
rect 4890 96976 4896 97028
rect 4948 97016 4954 97028
rect 47578 97016 47584 97028
rect 4948 96988 47440 97016
rect 47539 96988 47584 97016
rect 4948 96976 4954 96988
rect 1578 96948 1584 96960
rect 1539 96920 1584 96948
rect 1578 96908 1584 96920
rect 1636 96908 1642 96960
rect 3050 96948 3056 96960
rect 3011 96920 3056 96948
rect 3050 96908 3056 96920
rect 3108 96908 3114 96960
rect 11054 96908 11060 96960
rect 11112 96948 11118 96960
rect 11149 96951 11207 96957
rect 11149 96948 11161 96951
rect 11112 96920 11161 96948
rect 11112 96908 11118 96920
rect 11149 96917 11161 96920
rect 11195 96917 11207 96951
rect 16206 96948 16212 96960
rect 16167 96920 16212 96948
rect 11149 96911 11207 96917
rect 16206 96908 16212 96920
rect 16264 96908 16270 96960
rect 18782 96948 18788 96960
rect 18743 96920 18788 96948
rect 18782 96908 18788 96920
rect 18840 96908 18846 96960
rect 23566 96908 23572 96960
rect 23624 96948 23630 96960
rect 23753 96951 23811 96957
rect 23753 96948 23765 96951
rect 23624 96920 23765 96948
rect 23624 96908 23630 96920
rect 23753 96917 23765 96920
rect 23799 96917 23811 96951
rect 23753 96911 23811 96917
rect 24305 96951 24363 96957
rect 24305 96917 24317 96951
rect 24351 96948 24363 96951
rect 24486 96948 24492 96960
rect 24351 96920 24492 96948
rect 24351 96917 24363 96920
rect 24305 96911 24363 96917
rect 24486 96908 24492 96920
rect 24544 96908 24550 96960
rect 26602 96948 26608 96960
rect 26563 96920 26608 96948
rect 26602 96908 26608 96920
rect 26660 96908 26666 96960
rect 29178 96948 29184 96960
rect 29139 96920 29184 96948
rect 29178 96908 29184 96920
rect 29236 96908 29242 96960
rect 31846 96948 31852 96960
rect 31807 96920 31852 96948
rect 31846 96908 31852 96920
rect 31904 96908 31910 96960
rect 37090 96908 37096 96960
rect 37148 96948 37154 96960
rect 37185 96951 37243 96957
rect 37185 96948 37197 96951
rect 37148 96920 37197 96948
rect 37148 96908 37154 96920
rect 37185 96917 37197 96920
rect 37231 96917 37243 96951
rect 39666 96948 39672 96960
rect 39627 96920 39672 96948
rect 37185 96911 37243 96917
rect 39666 96908 39672 96920
rect 39724 96908 39730 96960
rect 42242 96948 42248 96960
rect 42203 96920 42248 96948
rect 42242 96908 42248 96920
rect 42300 96908 42306 96960
rect 44910 96948 44916 96960
rect 44871 96920 44916 96948
rect 44910 96908 44916 96920
rect 44968 96908 44974 96960
rect 45554 96908 45560 96960
rect 45612 96948 45618 96960
rect 45741 96951 45799 96957
rect 45741 96948 45753 96951
rect 45612 96920 45753 96948
rect 45612 96908 45618 96920
rect 45741 96917 45753 96920
rect 45787 96917 45799 96951
rect 47412 96948 47440 96988
rect 47578 96976 47584 96988
rect 47636 96976 47642 97028
rect 55186 97016 55214 97056
rect 55309 97053 55321 97056
rect 55355 97053 55367 97087
rect 56152 97084 56180 97115
rect 56410 97112 56416 97164
rect 56468 97152 56474 97164
rect 58713 97155 58771 97161
rect 58713 97152 58725 97155
rect 56468 97124 58725 97152
rect 56468 97112 56474 97124
rect 58713 97121 58725 97124
rect 58759 97121 58771 97155
rect 61378 97152 61384 97164
rect 61339 97124 61384 97152
rect 58713 97115 58771 97121
rect 61378 97112 61384 97124
rect 61436 97112 61442 97164
rect 62942 97152 62948 97164
rect 62903 97124 62948 97152
rect 62942 97112 62948 97124
rect 63000 97112 63006 97164
rect 63954 97152 63960 97164
rect 63915 97124 63960 97152
rect 63954 97112 63960 97124
rect 64012 97112 64018 97164
rect 66530 97152 66536 97164
rect 66491 97124 66536 97152
rect 66530 97112 66536 97124
rect 66588 97112 66594 97164
rect 68186 97112 68192 97164
rect 68244 97152 68250 97164
rect 68281 97155 68339 97161
rect 68281 97152 68293 97155
rect 68244 97124 68293 97152
rect 68244 97112 68250 97124
rect 68281 97121 68293 97124
rect 68327 97121 68339 97155
rect 69290 97152 69296 97164
rect 69251 97124 69296 97152
rect 68281 97115 68339 97121
rect 69290 97112 69296 97124
rect 69348 97112 69354 97164
rect 71038 97152 71044 97164
rect 70999 97124 71044 97152
rect 71038 97112 71044 97124
rect 71096 97112 71102 97164
rect 71777 97155 71835 97161
rect 71777 97121 71789 97155
rect 71823 97152 71835 97155
rect 71866 97152 71872 97164
rect 71823 97124 71872 97152
rect 71823 97121 71835 97124
rect 71777 97115 71835 97121
rect 71866 97112 71872 97124
rect 71924 97112 71930 97164
rect 72326 97112 72332 97164
rect 72384 97152 72390 97164
rect 72513 97155 72571 97161
rect 72513 97152 72525 97155
rect 72384 97124 72525 97152
rect 72384 97112 72390 97124
rect 72513 97121 72525 97124
rect 72559 97121 72571 97155
rect 72513 97115 72571 97121
rect 73338 97112 73344 97164
rect 73396 97152 73402 97164
rect 73617 97155 73675 97161
rect 73617 97152 73629 97155
rect 73396 97124 73629 97152
rect 73396 97112 73402 97124
rect 73617 97121 73629 97124
rect 73663 97121 73675 97155
rect 74442 97152 74448 97164
rect 74403 97124 74448 97152
rect 73617 97115 73675 97121
rect 74442 97112 74448 97124
rect 74500 97112 74506 97164
rect 75178 97152 75184 97164
rect 75139 97124 75184 97152
rect 75178 97112 75184 97124
rect 75236 97112 75242 97164
rect 77294 97152 77300 97164
rect 77255 97124 77300 97152
rect 77294 97112 77300 97124
rect 77352 97112 77358 97164
rect 78674 97112 78680 97164
rect 78732 97152 78738 97164
rect 78953 97155 79011 97161
rect 78953 97152 78965 97155
rect 78732 97124 78965 97152
rect 78732 97112 78738 97124
rect 78953 97121 78965 97124
rect 78999 97121 79011 97155
rect 79962 97152 79968 97164
rect 79923 97124 79968 97152
rect 78953 97115 79011 97121
rect 79962 97112 79968 97124
rect 80020 97112 80026 97164
rect 82170 97152 82176 97164
rect 82131 97124 82176 97152
rect 82170 97112 82176 97124
rect 82228 97112 82234 97164
rect 82906 97152 82912 97164
rect 82867 97124 82912 97152
rect 82906 97112 82912 97124
rect 82964 97112 82970 97164
rect 84565 97155 84623 97161
rect 84565 97121 84577 97155
rect 84611 97152 84623 97155
rect 84841 97155 84899 97161
rect 84841 97152 84853 97155
rect 84611 97124 84853 97152
rect 84611 97121 84623 97124
rect 84565 97115 84623 97121
rect 84841 97121 84853 97124
rect 84887 97152 84899 97155
rect 85022 97152 85028 97164
rect 84887 97124 85028 97152
rect 84887 97121 84899 97124
rect 84841 97115 84899 97121
rect 85022 97112 85028 97124
rect 85080 97112 85086 97164
rect 85482 97152 85488 97164
rect 85443 97124 85488 97152
rect 85482 97112 85488 97124
rect 85540 97112 85546 97164
rect 87506 97152 87512 97164
rect 87467 97124 87512 97152
rect 87506 97112 87512 97124
rect 87564 97112 87570 97164
rect 88150 97152 88156 97164
rect 88111 97124 88156 97152
rect 88150 97112 88156 97124
rect 88208 97112 88214 97164
rect 89714 97112 89720 97164
rect 89772 97152 89778 97164
rect 90085 97155 90143 97161
rect 90085 97152 90097 97155
rect 89772 97124 90097 97152
rect 89772 97112 89778 97124
rect 90085 97121 90097 97124
rect 90131 97121 90143 97155
rect 90284 97152 90312 97260
rect 90450 97248 90456 97260
rect 90508 97288 90514 97300
rect 95697 97291 95755 97297
rect 95697 97288 95709 97291
rect 90508 97260 90864 97288
rect 90508 97248 90514 97260
rect 90836 97229 90864 97260
rect 92584 97260 95709 97288
rect 90821 97223 90879 97229
rect 90821 97189 90833 97223
rect 90867 97189 90879 97223
rect 92474 97220 92480 97232
rect 92435 97192 92480 97220
rect 90821 97183 90879 97189
rect 92474 97180 92480 97192
rect 92532 97180 92538 97232
rect 92584 97152 92612 97260
rect 95697 97257 95709 97260
rect 95743 97288 95755 97291
rect 95743 97260 96108 97288
rect 95743 97257 95755 97260
rect 95697 97251 95755 97257
rect 95142 97220 95148 97232
rect 95103 97192 95148 97220
rect 95142 97180 95148 97192
rect 95200 97180 95206 97232
rect 96080 97229 96108 97260
rect 96065 97223 96123 97229
rect 96065 97189 96077 97223
rect 96111 97189 96123 97223
rect 97718 97220 97724 97232
rect 97679 97192 97724 97220
rect 96065 97183 96123 97189
rect 97718 97180 97724 97192
rect 97776 97180 97782 97232
rect 90284 97124 92612 97152
rect 92661 97155 92719 97161
rect 90085 97115 90143 97121
rect 92661 97121 92673 97155
rect 92707 97121 92719 97155
rect 92661 97115 92719 97121
rect 93121 97155 93179 97161
rect 93121 97121 93133 97155
rect 93167 97152 93179 97155
rect 93302 97152 93308 97164
rect 93167 97124 93308 97152
rect 93167 97121 93179 97124
rect 93121 97115 93179 97121
rect 69658 97084 69664 97096
rect 56152 97056 69664 97084
rect 55309 97047 55367 97053
rect 69658 97044 69664 97056
rect 69716 97044 69722 97096
rect 79134 97084 79140 97096
rect 79095 97056 79140 97084
rect 79134 97044 79140 97056
rect 79192 97044 79198 97096
rect 84102 97044 84108 97096
rect 84160 97084 84166 97096
rect 85669 97087 85727 97093
rect 85669 97084 85681 97087
rect 84160 97056 85681 97084
rect 84160 97044 84166 97056
rect 85669 97053 85681 97056
rect 85715 97053 85727 97087
rect 85669 97047 85727 97053
rect 57974 97016 57980 97028
rect 47688 96988 55214 97016
rect 57935 96988 57980 97016
rect 47688 96948 47716 96988
rect 57974 96976 57980 96988
rect 58032 96976 58038 97028
rect 65889 97019 65947 97025
rect 65889 96985 65901 97019
rect 65935 97016 65947 97019
rect 65978 97016 65984 97028
rect 65935 96988 65984 97016
rect 65935 96985 65947 96988
rect 65889 96979 65947 96985
rect 65978 96976 65984 96988
rect 66036 96976 66042 97028
rect 73801 97019 73859 97025
rect 73801 96985 73813 97019
rect 73847 97016 73859 97019
rect 80698 97016 80704 97028
rect 73847 96988 80704 97016
rect 73847 96985 73859 96988
rect 73801 96979 73859 96985
rect 80698 96976 80704 96988
rect 80756 96976 80762 97028
rect 88334 97016 88340 97028
rect 88295 96988 88340 97016
rect 88334 96976 88340 96988
rect 88392 96976 88398 97028
rect 90634 97016 90640 97028
rect 90595 96988 90640 97016
rect 90634 96976 90640 96988
rect 90692 96976 90698 97028
rect 52730 96948 52736 96960
rect 47412 96920 47716 96948
rect 52691 96920 52736 96948
rect 45741 96911 45799 96917
rect 52730 96908 52736 96920
rect 52788 96908 52794 96960
rect 60734 96948 60740 96960
rect 60695 96920 60740 96948
rect 60734 96908 60740 96920
rect 60792 96908 60798 96960
rect 63126 96948 63132 96960
rect 63087 96920 63132 96948
rect 63126 96908 63132 96920
rect 63184 96908 63190 96960
rect 71130 96948 71136 96960
rect 71091 96920 71136 96948
rect 71130 96908 71136 96920
rect 71188 96908 71194 96960
rect 71774 96908 71780 96960
rect 71832 96948 71838 96960
rect 71869 96951 71927 96957
rect 71869 96948 71881 96951
rect 71832 96920 71881 96948
rect 71832 96908 71838 96920
rect 71869 96917 71881 96920
rect 71915 96917 71927 96951
rect 71869 96911 71927 96917
rect 72510 96908 72516 96960
rect 72568 96948 72574 96960
rect 75273 96951 75331 96957
rect 75273 96948 75285 96951
rect 72568 96920 75285 96948
rect 72568 96908 72574 96920
rect 75273 96917 75285 96920
rect 75319 96917 75331 96951
rect 75273 96911 75331 96917
rect 76374 96908 76380 96960
rect 76432 96948 76438 96960
rect 76469 96951 76527 96957
rect 76469 96948 76481 96951
rect 76432 96920 76481 96948
rect 76432 96908 76438 96920
rect 76469 96917 76481 96920
rect 76515 96917 76527 96951
rect 76469 96911 76527 96917
rect 82814 96908 82820 96960
rect 82872 96948 82878 96960
rect 83001 96951 83059 96957
rect 83001 96948 83013 96951
rect 82872 96920 83013 96948
rect 82872 96908 82878 96920
rect 83001 96917 83013 96920
rect 83047 96917 83059 96951
rect 85022 96948 85028 96960
rect 84983 96920 85028 96948
rect 83001 96911 83059 96917
rect 85022 96908 85028 96920
rect 85080 96908 85086 96960
rect 87233 96951 87291 96957
rect 87233 96917 87245 96951
rect 87279 96948 87291 96951
rect 87506 96948 87512 96960
rect 87279 96920 87512 96948
rect 87279 96917 87291 96920
rect 87233 96911 87291 96917
rect 87506 96908 87512 96920
rect 87564 96948 87570 96960
rect 87693 96951 87751 96957
rect 87693 96948 87705 96951
rect 87564 96920 87705 96948
rect 87564 96908 87570 96920
rect 87693 96917 87705 96920
rect 87739 96917 87751 96951
rect 87693 96911 87751 96917
rect 89714 96908 89720 96960
rect 89772 96948 89778 96960
rect 92290 96948 92296 96960
rect 89772 96920 89817 96948
rect 92251 96920 92296 96948
rect 89772 96908 89778 96920
rect 92290 96908 92296 96920
rect 92348 96948 92354 96960
rect 92676 96948 92704 97115
rect 93302 97112 93308 97124
rect 93360 97152 93366 97164
rect 93397 97155 93455 97161
rect 93397 97152 93409 97155
rect 93360 97124 93409 97152
rect 93360 97112 93366 97124
rect 93397 97121 93409 97124
rect 93443 97121 93455 97155
rect 93397 97115 93455 97121
rect 95329 97155 95387 97161
rect 95329 97121 95341 97155
rect 95375 97121 95387 97155
rect 95329 97115 95387 97121
rect 97905 97155 97963 97161
rect 97905 97121 97917 97155
rect 97951 97121 97963 97155
rect 97905 97115 97963 97121
rect 92750 96976 92756 97028
rect 92808 97016 92814 97028
rect 93213 97019 93271 97025
rect 93213 97016 93225 97019
rect 92808 96988 93225 97016
rect 92808 96976 92814 96988
rect 93213 96985 93225 96988
rect 93259 96985 93271 97019
rect 93213 96979 93271 96985
rect 92845 96951 92903 96957
rect 92845 96948 92857 96951
rect 92348 96920 92857 96948
rect 92348 96908 92354 96920
rect 92845 96917 92857 96920
rect 92891 96917 92903 96951
rect 94958 96948 94964 96960
rect 94919 96920 94964 96948
rect 92845 96911 92903 96917
rect 94958 96908 94964 96920
rect 95016 96948 95022 96960
rect 95344 96948 95372 97115
rect 95878 97016 95884 97028
rect 95839 96988 95884 97016
rect 95878 96976 95884 96988
rect 95936 96976 95942 97028
rect 95513 96951 95571 96957
rect 95513 96948 95525 96951
rect 95016 96920 95525 96948
rect 95016 96908 95022 96920
rect 95513 96917 95525 96920
rect 95559 96917 95571 96951
rect 97534 96948 97540 96960
rect 97495 96920 97540 96948
rect 95513 96911 95571 96917
rect 97534 96908 97540 96920
rect 97592 96948 97598 96960
rect 97920 96948 97948 97115
rect 98089 96951 98147 96957
rect 98089 96948 98101 96951
rect 97592 96920 98101 96948
rect 97592 96908 97598 96920
rect 98089 96917 98101 96920
rect 98135 96917 98147 96951
rect 98089 96911 98147 96917
rect 1104 96858 98808 96880
rect 1104 96806 4246 96858
rect 4298 96806 4310 96858
rect 4362 96806 4374 96858
rect 4426 96806 4438 96858
rect 4490 96806 34966 96858
rect 35018 96806 35030 96858
rect 35082 96806 35094 96858
rect 35146 96806 35158 96858
rect 35210 96806 65686 96858
rect 65738 96806 65750 96858
rect 65802 96806 65814 96858
rect 65866 96806 65878 96858
rect 65930 96806 96406 96858
rect 96458 96806 96470 96858
rect 96522 96806 96534 96858
rect 96586 96806 96598 96858
rect 96650 96806 98808 96858
rect 1104 96784 98808 96806
rect 16025 96747 16083 96753
rect 16025 96713 16037 96747
rect 16071 96744 16083 96747
rect 16298 96744 16304 96756
rect 16071 96716 16304 96744
rect 16071 96713 16083 96716
rect 16025 96707 16083 96713
rect 16298 96704 16304 96716
rect 16356 96704 16362 96756
rect 21358 96744 21364 96756
rect 16546 96716 21364 96744
rect 14458 96636 14464 96688
rect 14516 96676 14522 96688
rect 16546 96676 16574 96716
rect 21358 96704 21364 96716
rect 21416 96704 21422 96756
rect 34606 96704 34612 96756
rect 34664 96744 34670 96756
rect 79134 96744 79140 96756
rect 34664 96716 79140 96744
rect 34664 96704 34670 96716
rect 79134 96704 79140 96716
rect 79192 96704 79198 96756
rect 14516 96648 16574 96676
rect 14516 96636 14522 96648
rect 40678 96636 40684 96688
rect 40736 96676 40742 96688
rect 43438 96676 43444 96688
rect 40736 96648 43444 96676
rect 40736 96636 40742 96648
rect 43438 96636 43444 96648
rect 43496 96636 43502 96688
rect 2038 96568 2044 96620
rect 2096 96608 2102 96620
rect 2317 96611 2375 96617
rect 2317 96608 2329 96611
rect 2096 96580 2329 96608
rect 2096 96568 2102 96580
rect 2317 96577 2329 96580
rect 2363 96577 2375 96611
rect 2317 96571 2375 96577
rect 4706 96568 4712 96620
rect 4764 96608 4770 96620
rect 4985 96611 5043 96617
rect 4985 96608 4997 96611
rect 4764 96580 4997 96608
rect 4764 96568 4770 96580
rect 4985 96577 4997 96580
rect 5031 96577 5043 96611
rect 7282 96608 7288 96620
rect 7243 96580 7288 96608
rect 4985 96571 5043 96577
rect 7282 96568 7288 96580
rect 7340 96568 7346 96620
rect 9858 96568 9864 96620
rect 9916 96608 9922 96620
rect 10137 96611 10195 96617
rect 10137 96608 10149 96611
rect 9916 96580 10149 96608
rect 9916 96568 9922 96580
rect 10137 96577 10149 96580
rect 10183 96577 10195 96611
rect 10137 96571 10195 96577
rect 12526 96568 12532 96620
rect 12584 96608 12590 96620
rect 12805 96611 12863 96617
rect 12805 96608 12817 96611
rect 12584 96580 12817 96608
rect 12584 96568 12590 96580
rect 12805 96577 12817 96580
rect 12851 96577 12863 96611
rect 12805 96571 12863 96577
rect 15102 96568 15108 96620
rect 15160 96608 15166 96620
rect 15381 96611 15439 96617
rect 15381 96608 15393 96611
rect 15160 96580 15393 96608
rect 15160 96568 15166 96580
rect 15381 96577 15393 96580
rect 15427 96577 15439 96611
rect 15381 96571 15439 96577
rect 17770 96568 17776 96620
rect 17828 96608 17834 96620
rect 18049 96611 18107 96617
rect 18049 96608 18061 96611
rect 17828 96580 18061 96608
rect 17828 96568 17834 96580
rect 18049 96577 18061 96580
rect 18095 96577 18107 96611
rect 18049 96571 18107 96577
rect 22922 96568 22928 96620
rect 22980 96608 22986 96620
rect 23201 96611 23259 96617
rect 23201 96608 23213 96611
rect 22980 96580 23213 96608
rect 22980 96568 22986 96580
rect 23201 96577 23213 96580
rect 23247 96577 23259 96611
rect 23201 96571 23259 96577
rect 25590 96568 25596 96620
rect 25648 96608 25654 96620
rect 25869 96611 25927 96617
rect 25869 96608 25881 96611
rect 25648 96580 25881 96608
rect 25648 96568 25654 96580
rect 25869 96577 25881 96580
rect 25915 96577 25927 96611
rect 25869 96571 25927 96577
rect 33410 96568 33416 96620
rect 33468 96608 33474 96620
rect 33689 96611 33747 96617
rect 33689 96608 33701 96611
rect 33468 96580 33701 96608
rect 33468 96568 33474 96580
rect 33689 96577 33701 96580
rect 33735 96577 33747 96611
rect 33689 96571 33747 96577
rect 35986 96568 35992 96620
rect 36044 96608 36050 96620
rect 36265 96611 36323 96617
rect 36265 96608 36277 96611
rect 36044 96580 36277 96608
rect 36044 96568 36050 96580
rect 36265 96577 36277 96580
rect 36311 96577 36323 96611
rect 36265 96571 36323 96577
rect 38562 96568 38568 96620
rect 38620 96608 38626 96620
rect 38841 96611 38899 96617
rect 38841 96608 38853 96611
rect 38620 96580 38853 96608
rect 38620 96568 38626 96580
rect 38841 96577 38853 96580
rect 38887 96577 38899 96611
rect 38841 96571 38899 96577
rect 41230 96568 41236 96620
rect 41288 96608 41294 96620
rect 41509 96611 41567 96617
rect 41509 96608 41521 96611
rect 41288 96580 41521 96608
rect 41288 96568 41294 96580
rect 41509 96577 41521 96580
rect 41555 96577 41567 96611
rect 41509 96571 41567 96577
rect 43806 96568 43812 96620
rect 43864 96608 43870 96620
rect 44085 96611 44143 96617
rect 44085 96608 44097 96611
rect 43864 96580 44097 96608
rect 43864 96568 43870 96580
rect 44085 96577 44097 96580
rect 44131 96577 44143 96611
rect 44085 96571 44143 96577
rect 49050 96568 49056 96620
rect 49108 96608 49114 96620
rect 49329 96611 49387 96617
rect 49329 96608 49341 96611
rect 49108 96580 49341 96608
rect 49108 96568 49114 96580
rect 49329 96577 49341 96580
rect 49375 96577 49387 96611
rect 49329 96571 49387 96577
rect 51626 96568 51632 96620
rect 51684 96608 51690 96620
rect 51905 96611 51963 96617
rect 51905 96608 51917 96611
rect 51684 96580 51917 96608
rect 51684 96568 51690 96580
rect 51905 96577 51917 96580
rect 51951 96577 51963 96611
rect 51905 96571 51963 96577
rect 54294 96568 54300 96620
rect 54352 96608 54358 96620
rect 54573 96611 54631 96617
rect 54573 96608 54585 96611
rect 54352 96580 54585 96608
rect 54352 96568 54358 96580
rect 54573 96577 54585 96580
rect 54619 96577 54631 96611
rect 54573 96571 54631 96577
rect 56870 96568 56876 96620
rect 56928 96608 56934 96620
rect 57149 96611 57207 96617
rect 57149 96608 57161 96611
rect 56928 96580 57161 96608
rect 56928 96568 56934 96580
rect 57149 96577 57161 96580
rect 57195 96577 57207 96611
rect 57149 96571 57207 96577
rect 59446 96568 59452 96620
rect 59504 96608 59510 96620
rect 59725 96611 59783 96617
rect 59725 96608 59737 96611
rect 59504 96580 59737 96608
rect 59504 96568 59510 96580
rect 59725 96577 59737 96580
rect 59771 96577 59783 96611
rect 59725 96571 59783 96577
rect 62114 96568 62120 96620
rect 62172 96608 62178 96620
rect 62393 96611 62451 96617
rect 62393 96608 62405 96611
rect 62172 96580 62405 96608
rect 62172 96568 62178 96580
rect 62393 96577 62405 96580
rect 62439 96577 62451 96611
rect 62393 96571 62451 96577
rect 64690 96568 64696 96620
rect 64748 96608 64754 96620
rect 64969 96611 65027 96617
rect 64969 96608 64981 96611
rect 64748 96580 64981 96608
rect 64748 96568 64754 96580
rect 64969 96577 64981 96580
rect 65015 96577 65027 96611
rect 64969 96571 65027 96577
rect 67266 96568 67272 96620
rect 67324 96608 67330 96620
rect 71130 96608 71136 96620
rect 67324 96580 71136 96608
rect 67324 96568 67330 96580
rect 71130 96568 71136 96580
rect 71188 96568 71194 96620
rect 75086 96568 75092 96620
rect 75144 96608 75150 96620
rect 75365 96611 75423 96617
rect 75365 96608 75377 96611
rect 75144 96580 75377 96608
rect 75144 96568 75150 96580
rect 75365 96577 75377 96580
rect 75411 96577 75423 96611
rect 75365 96571 75423 96577
rect 80330 96568 80336 96620
rect 80388 96608 80394 96620
rect 84102 96608 84108 96620
rect 80388 96580 84108 96608
rect 80388 96568 80394 96580
rect 84102 96568 84108 96580
rect 84160 96568 84166 96620
rect 85574 96568 85580 96620
rect 85632 96608 85638 96620
rect 90634 96608 90640 96620
rect 85632 96580 90640 96608
rect 85632 96568 85638 96580
rect 90634 96568 90640 96580
rect 90692 96568 90698 96620
rect 90818 96568 90824 96620
rect 90876 96608 90882 96620
rect 93394 96608 93400 96620
rect 90876 96580 93256 96608
rect 93355 96580 93400 96608
rect 90876 96568 90882 96580
rect 20438 96500 20444 96552
rect 20496 96540 20502 96552
rect 23566 96540 23572 96552
rect 20496 96512 23572 96540
rect 20496 96500 20502 96512
rect 23566 96500 23572 96512
rect 23624 96500 23630 96552
rect 23842 96540 23848 96552
rect 23803 96512 23848 96540
rect 23842 96500 23848 96512
rect 23900 96500 23906 96552
rect 38746 96500 38752 96552
rect 38804 96540 38810 96552
rect 43901 96543 43959 96549
rect 43901 96540 43913 96543
rect 38804 96512 43913 96540
rect 38804 96500 38810 96512
rect 43901 96509 43913 96512
rect 43947 96509 43959 96543
rect 43901 96503 43959 96509
rect 46106 96500 46112 96552
rect 46164 96540 46170 96552
rect 46293 96543 46351 96549
rect 46293 96540 46305 96543
rect 46164 96512 46305 96540
rect 46164 96500 46170 96512
rect 46293 96509 46305 96512
rect 46339 96509 46351 96543
rect 46293 96503 46351 96509
rect 46474 96500 46480 96552
rect 46532 96540 46538 96552
rect 46615 96543 46673 96549
rect 46615 96540 46627 96543
rect 46532 96512 46627 96540
rect 46532 96500 46538 96512
rect 46615 96509 46627 96512
rect 46661 96509 46673 96543
rect 46750 96540 46756 96552
rect 46711 96512 46756 96540
rect 46615 96503 46673 96509
rect 46750 96500 46756 96512
rect 46808 96500 46814 96552
rect 47026 96540 47032 96552
rect 46987 96512 47032 96540
rect 47026 96500 47032 96512
rect 47084 96500 47090 96552
rect 47210 96540 47216 96552
rect 47171 96512 47216 96540
rect 47210 96500 47216 96512
rect 47268 96500 47274 96552
rect 70762 96540 70768 96552
rect 70723 96512 70768 96540
rect 70762 96500 70768 96512
rect 70820 96500 70826 96552
rect 81253 96543 81311 96549
rect 81253 96509 81265 96543
rect 81299 96540 81311 96543
rect 81342 96540 81348 96552
rect 81299 96512 81348 96540
rect 81299 96509 81311 96512
rect 81253 96503 81311 96509
rect 81342 96500 81348 96512
rect 81400 96500 81406 96552
rect 83826 96540 83832 96552
rect 83787 96512 83832 96540
rect 83826 96500 83832 96512
rect 83884 96500 83890 96552
rect 86402 96540 86408 96552
rect 86363 96512 86408 96540
rect 86402 96500 86408 96512
rect 86460 96500 86466 96552
rect 89070 96540 89076 96552
rect 89031 96512 89076 96540
rect 89070 96500 89076 96512
rect 89128 96500 89134 96552
rect 91646 96540 91652 96552
rect 91607 96512 91652 96540
rect 91646 96500 91652 96512
rect 91704 96500 91710 96552
rect 93228 96540 93256 96580
rect 93394 96568 93400 96580
rect 93452 96568 93458 96620
rect 95878 96608 95884 96620
rect 94056 96580 95884 96608
rect 94056 96540 94084 96580
rect 95878 96568 95884 96580
rect 95936 96568 95942 96620
rect 95970 96568 95976 96620
rect 96028 96608 96034 96620
rect 96249 96611 96307 96617
rect 96249 96608 96261 96611
rect 96028 96580 96261 96608
rect 96028 96568 96034 96580
rect 96249 96577 96261 96580
rect 96295 96577 96307 96611
rect 96249 96571 96307 96577
rect 98089 96611 98147 96617
rect 98089 96577 98101 96611
rect 98135 96608 98147 96611
rect 98638 96608 98644 96620
rect 98135 96580 98644 96608
rect 98135 96577 98147 96580
rect 98089 96571 98147 96577
rect 98638 96568 98644 96580
rect 98696 96568 98702 96620
rect 94222 96540 94228 96552
rect 93228 96512 94084 96540
rect 94183 96512 94228 96540
rect 94222 96500 94228 96512
rect 94280 96500 94286 96552
rect 97353 96543 97411 96549
rect 97353 96509 97365 96543
rect 97399 96540 97411 96543
rect 99466 96540 99472 96552
rect 97399 96512 99472 96540
rect 97399 96509 97411 96512
rect 97353 96503 97411 96509
rect 99466 96500 99472 96512
rect 99524 96500 99530 96552
rect 2130 96472 2136 96484
rect 2091 96444 2136 96472
rect 2130 96432 2136 96444
rect 2188 96432 2194 96484
rect 4798 96472 4804 96484
rect 4759 96444 4804 96472
rect 4798 96432 4804 96444
rect 4856 96432 4862 96484
rect 7469 96475 7527 96481
rect 7469 96441 7481 96475
rect 7515 96441 7527 96475
rect 9950 96472 9956 96484
rect 9911 96444 9956 96472
rect 7469 96435 7527 96441
rect 7098 96404 7104 96416
rect 7059 96376 7104 96404
rect 7098 96364 7104 96376
rect 7156 96404 7162 96416
rect 7484 96404 7512 96435
rect 9950 96432 9956 96444
rect 10008 96432 10014 96484
rect 12618 96472 12624 96484
rect 12579 96444 12624 96472
rect 12618 96432 12624 96444
rect 12676 96432 12682 96484
rect 15197 96475 15255 96481
rect 15197 96441 15209 96475
rect 15243 96472 15255 96475
rect 17862 96472 17868 96484
rect 15243 96444 16574 96472
rect 17823 96444 17868 96472
rect 15243 96441 15255 96444
rect 15197 96435 15255 96441
rect 7156 96376 7512 96404
rect 16546 96404 16574 96444
rect 17862 96432 17868 96444
rect 17920 96432 17926 96484
rect 23014 96472 23020 96484
rect 22975 96444 23020 96472
rect 23014 96432 23020 96444
rect 23072 96432 23078 96484
rect 25682 96472 25688 96484
rect 25643 96444 25688 96472
rect 25682 96432 25688 96444
rect 25740 96432 25746 96484
rect 30374 96432 30380 96484
rect 30432 96472 30438 96484
rect 33505 96475 33563 96481
rect 33505 96472 33517 96475
rect 30432 96444 33517 96472
rect 30432 96432 30438 96444
rect 33505 96441 33517 96444
rect 33551 96441 33563 96475
rect 36078 96472 36084 96484
rect 36039 96444 36084 96472
rect 33505 96435 33563 96441
rect 36078 96432 36084 96444
rect 36136 96432 36142 96484
rect 38654 96472 38660 96484
rect 38615 96444 38660 96472
rect 38654 96432 38660 96444
rect 38712 96432 38718 96484
rect 41322 96472 41328 96484
rect 41283 96444 41328 96472
rect 41322 96432 41328 96444
rect 41380 96432 41386 96484
rect 49142 96472 49148 96484
rect 49103 96444 49148 96472
rect 49142 96432 49148 96444
rect 49200 96432 49206 96484
rect 51718 96472 51724 96484
rect 51679 96444 51724 96472
rect 51718 96432 51724 96444
rect 51776 96432 51782 96484
rect 54386 96472 54392 96484
rect 54347 96444 54392 96472
rect 54386 96432 54392 96444
rect 54444 96432 54450 96484
rect 56962 96472 56968 96484
rect 56923 96444 56968 96472
rect 56962 96432 56968 96444
rect 57020 96432 57026 96484
rect 59538 96472 59544 96484
rect 59499 96444 59544 96472
rect 59538 96432 59544 96444
rect 59596 96432 59602 96484
rect 62206 96472 62212 96484
rect 62167 96444 62212 96472
rect 62206 96432 62212 96444
rect 62264 96432 62270 96484
rect 64782 96472 64788 96484
rect 64743 96444 64788 96472
rect 64782 96432 64788 96444
rect 64840 96432 64846 96484
rect 74534 96432 74540 96484
rect 74592 96472 74598 96484
rect 75181 96475 75239 96481
rect 75181 96472 75193 96475
rect 74592 96444 75193 96472
rect 74592 96432 74598 96444
rect 75181 96441 75193 96444
rect 75227 96441 75239 96475
rect 75181 96435 75239 96441
rect 77754 96432 77760 96484
rect 77812 96472 77818 96484
rect 82814 96472 82820 96484
rect 77812 96444 82820 96472
rect 77812 96432 77818 96444
rect 82814 96432 82820 96444
rect 82872 96432 82878 96484
rect 88242 96432 88248 96484
rect 88300 96472 88306 96484
rect 92750 96472 92756 96484
rect 88300 96444 92756 96472
rect 88300 96432 88306 96444
rect 92750 96432 92756 96444
rect 92808 96432 92814 96484
rect 93581 96475 93639 96481
rect 93581 96441 93593 96475
rect 93627 96441 93639 96475
rect 96062 96472 96068 96484
rect 96023 96444 96068 96472
rect 93581 96435 93639 96441
rect 20438 96404 20444 96416
rect 16546 96376 20444 96404
rect 7156 96364 7162 96376
rect 20438 96364 20444 96376
rect 20496 96364 20502 96416
rect 24026 96404 24032 96416
rect 23987 96376 24032 96404
rect 24026 96364 24032 96376
rect 24084 96364 24090 96416
rect 47486 96404 47492 96416
rect 47447 96376 47492 96404
rect 47486 96364 47492 96376
rect 47544 96364 47550 96416
rect 70854 96364 70860 96416
rect 70912 96404 70918 96416
rect 70949 96407 71007 96413
rect 70949 96404 70961 96407
rect 70912 96376 70961 96404
rect 70912 96364 70918 96376
rect 70949 96373 70961 96376
rect 70995 96373 71007 96407
rect 81434 96404 81440 96416
rect 81395 96376 81440 96404
rect 70949 96367 71007 96373
rect 81434 96364 81440 96376
rect 81492 96364 81498 96416
rect 82998 96364 83004 96416
rect 83056 96404 83062 96416
rect 88334 96404 88340 96416
rect 83056 96376 88340 96404
rect 83056 96364 83062 96376
rect 88334 96364 88340 96376
rect 88392 96364 88398 96416
rect 93210 96404 93216 96416
rect 93171 96376 93216 96404
rect 93210 96364 93216 96376
rect 93268 96404 93274 96416
rect 93596 96404 93624 96435
rect 96062 96432 96068 96444
rect 96120 96432 96126 96484
rect 97169 96475 97227 96481
rect 97169 96441 97181 96475
rect 97215 96441 97227 96475
rect 97169 96435 97227 96441
rect 97721 96475 97779 96481
rect 97721 96441 97733 96475
rect 97767 96472 97779 96475
rect 97902 96472 97908 96484
rect 97767 96444 97908 96472
rect 97767 96441 97779 96444
rect 97721 96435 97779 96441
rect 93765 96407 93823 96413
rect 93765 96404 93777 96407
rect 93268 96376 93777 96404
rect 93268 96364 93274 96376
rect 93765 96373 93777 96376
rect 93811 96373 93823 96407
rect 93765 96367 93823 96373
rect 95878 96364 95884 96416
rect 95936 96404 95942 96416
rect 96893 96407 96951 96413
rect 96893 96404 96905 96407
rect 95936 96376 96905 96404
rect 95936 96364 95942 96376
rect 96893 96373 96905 96376
rect 96939 96404 96951 96407
rect 97184 96404 97212 96435
rect 97902 96432 97908 96444
rect 97960 96472 97966 96484
rect 98181 96475 98239 96481
rect 98181 96472 98193 96475
rect 97960 96444 98193 96472
rect 97960 96432 97966 96444
rect 98181 96441 98193 96444
rect 98227 96441 98239 96475
rect 98181 96435 98239 96441
rect 97445 96407 97503 96413
rect 97445 96404 97457 96407
rect 96939 96376 97457 96404
rect 96939 96373 96951 96376
rect 96893 96367 96951 96373
rect 97445 96373 97457 96376
rect 97491 96373 97503 96407
rect 97445 96367 97503 96373
rect 1104 96314 98808 96336
rect 1104 96262 19606 96314
rect 19658 96262 19670 96314
rect 19722 96262 19734 96314
rect 19786 96262 19798 96314
rect 19850 96262 50326 96314
rect 50378 96262 50390 96314
rect 50442 96262 50454 96314
rect 50506 96262 50518 96314
rect 50570 96262 81046 96314
rect 81098 96262 81110 96314
rect 81162 96262 81174 96314
rect 81226 96262 81238 96314
rect 81290 96262 98808 96314
rect 1104 96240 98808 96262
rect 2130 96160 2136 96212
rect 2188 96200 2194 96212
rect 14550 96200 14556 96212
rect 2188 96172 14556 96200
rect 2188 96160 2194 96172
rect 14550 96160 14556 96172
rect 14608 96160 14614 96212
rect 46382 96160 46388 96212
rect 46440 96200 46446 96212
rect 46569 96203 46627 96209
rect 46569 96200 46581 96203
rect 46440 96172 46581 96200
rect 46440 96160 46446 96172
rect 46569 96169 46581 96172
rect 46615 96169 46627 96203
rect 46569 96163 46627 96169
rect 49142 96160 49148 96212
rect 49200 96200 49206 96212
rect 60090 96200 60096 96212
rect 49200 96172 60096 96200
rect 49200 96160 49206 96172
rect 60090 96160 60096 96172
rect 60148 96160 60154 96212
rect 26513 96067 26571 96073
rect 26513 96033 26525 96067
rect 26559 96064 26571 96067
rect 30282 96064 30288 96076
rect 26559 96036 30288 96064
rect 26559 96033 26571 96036
rect 26513 96027 26571 96033
rect 30282 96024 30288 96036
rect 30340 96024 30346 96076
rect 46477 96067 46535 96073
rect 46477 96033 46489 96067
rect 46523 96064 46535 96067
rect 46842 96064 46848 96076
rect 46523 96036 46848 96064
rect 46523 96033 46535 96036
rect 46477 96027 46535 96033
rect 46842 96024 46848 96036
rect 46900 96024 46906 96076
rect 57422 96064 57428 96076
rect 57383 96036 57428 96064
rect 57422 96024 57428 96036
rect 57480 96024 57486 96076
rect 57790 96064 57796 96076
rect 57751 96036 57796 96064
rect 57790 96024 57796 96036
rect 57848 96024 57854 96076
rect 58158 96064 58164 96076
rect 58119 96036 58164 96064
rect 58158 96024 58164 96036
rect 58216 96024 58222 96076
rect 83369 96067 83427 96073
rect 83369 96033 83381 96067
rect 83415 96033 83427 96067
rect 83369 96027 83427 96033
rect 26789 95999 26847 96005
rect 26789 95965 26801 95999
rect 26835 95996 26847 95999
rect 26878 95996 26884 96008
rect 26835 95968 26884 95996
rect 26835 95965 26847 95968
rect 26789 95959 26847 95965
rect 26878 95956 26884 95968
rect 26936 95956 26942 96008
rect 28169 95999 28227 96005
rect 28169 95965 28181 95999
rect 28215 95996 28227 95999
rect 30374 95996 30380 96008
rect 28215 95968 30380 95996
rect 28215 95965 28227 95968
rect 28169 95959 28227 95965
rect 30374 95956 30380 95968
rect 30432 95956 30438 96008
rect 57606 95996 57612 96008
rect 57567 95968 57612 95996
rect 57606 95956 57612 95968
rect 57664 95956 57670 96008
rect 58069 95999 58127 96005
rect 58069 95965 58081 95999
rect 58115 95965 58127 95999
rect 58069 95959 58127 95965
rect 82909 95999 82967 96005
rect 82909 95965 82921 95999
rect 82955 95965 82967 95999
rect 82909 95959 82967 95965
rect 30650 95888 30656 95940
rect 30708 95928 30714 95940
rect 30708 95900 55214 95928
rect 30708 95888 30714 95900
rect 55186 95860 55214 95900
rect 56502 95888 56508 95940
rect 56560 95928 56566 95940
rect 58084 95928 58112 95959
rect 58526 95928 58532 95940
rect 56560 95900 58112 95928
rect 58487 95900 58532 95928
rect 56560 95888 56566 95900
rect 58526 95888 58532 95900
rect 58584 95888 58590 95940
rect 82924 95928 82952 95959
rect 64846 95900 82952 95928
rect 83384 95928 83412 96027
rect 83458 96024 83464 96076
rect 83516 96064 83522 96076
rect 83737 96067 83795 96073
rect 83737 96064 83749 96067
rect 83516 96036 83749 96064
rect 83516 96024 83522 96036
rect 83737 96033 83749 96036
rect 83783 96033 83795 96067
rect 96890 96064 96896 96076
rect 96851 96036 96896 96064
rect 83737 96027 83795 96033
rect 96890 96024 96896 96036
rect 96948 96024 96954 96076
rect 83826 95996 83832 96008
rect 83787 95968 83832 95996
rect 83826 95956 83832 95968
rect 83884 95956 83890 96008
rect 83918 95928 83924 95940
rect 83384 95900 83924 95928
rect 64846 95860 64874 95900
rect 83918 95888 83924 95900
rect 83976 95888 83982 95940
rect 55186 95832 64874 95860
rect 1104 95770 98808 95792
rect 1104 95718 4246 95770
rect 4298 95718 4310 95770
rect 4362 95718 4374 95770
rect 4426 95718 4438 95770
rect 4490 95718 34966 95770
rect 35018 95718 35030 95770
rect 35082 95718 35094 95770
rect 35146 95718 35158 95770
rect 35210 95718 65686 95770
rect 65738 95718 65750 95770
rect 65802 95718 65814 95770
rect 65866 95718 65878 95770
rect 65930 95718 96406 95770
rect 96458 95718 96470 95770
rect 96522 95718 96534 95770
rect 96586 95718 96598 95770
rect 96650 95718 98808 95770
rect 1104 95696 98808 95718
rect 46750 95616 46756 95668
rect 46808 95656 46814 95668
rect 88978 95656 88984 95668
rect 46808 95628 88984 95656
rect 46808 95616 46814 95628
rect 88978 95616 88984 95628
rect 89036 95616 89042 95668
rect 53834 95588 53840 95600
rect 34992 95560 45554 95588
rect 53795 95560 53840 95588
rect 34992 95461 35020 95560
rect 35069 95523 35127 95529
rect 35069 95489 35081 95523
rect 35115 95520 35127 95523
rect 45526 95520 45554 95560
rect 53834 95548 53840 95560
rect 53892 95588 53898 95600
rect 54205 95591 54263 95597
rect 54205 95588 54217 95591
rect 53892 95560 54217 95588
rect 53892 95548 53898 95560
rect 54205 95557 54217 95560
rect 54251 95557 54263 95591
rect 54205 95551 54263 95557
rect 57974 95520 57980 95532
rect 35115 95492 35894 95520
rect 45526 95492 57980 95520
rect 35115 95489 35127 95492
rect 35069 95483 35127 95489
rect 10137 95455 10195 95461
rect 10137 95421 10149 95455
rect 10183 95452 10195 95455
rect 34977 95455 35035 95461
rect 10183 95424 16574 95452
rect 10183 95421 10195 95424
rect 10137 95415 10195 95421
rect 10870 95384 10876 95396
rect 10831 95356 10876 95384
rect 10870 95344 10876 95356
rect 10928 95344 10934 95396
rect 16546 95384 16574 95424
rect 34977 95421 34989 95455
rect 35023 95421 35035 95455
rect 35342 95452 35348 95464
rect 35303 95424 35348 95452
rect 34977 95415 35035 95421
rect 35342 95412 35348 95424
rect 35400 95412 35406 95464
rect 35529 95455 35587 95461
rect 35529 95421 35541 95455
rect 35575 95421 35587 95455
rect 35866 95452 35894 95492
rect 57974 95480 57980 95492
rect 58032 95480 58038 95532
rect 66898 95452 66904 95464
rect 35866 95424 66904 95452
rect 35529 95415 35587 95421
rect 31386 95384 31392 95396
rect 16546 95356 31392 95384
rect 31386 95344 31392 95356
rect 31444 95344 31450 95396
rect 35544 95384 35572 95415
rect 66898 95412 66904 95424
rect 66956 95412 66962 95464
rect 61654 95384 61660 95396
rect 35544 95356 61660 95384
rect 61654 95344 61660 95356
rect 61712 95344 61718 95396
rect 34609 95319 34667 95325
rect 34609 95285 34621 95319
rect 34655 95316 34667 95319
rect 96154 95316 96160 95328
rect 34655 95288 96160 95316
rect 34655 95285 34667 95288
rect 34609 95279 34667 95285
rect 96154 95276 96160 95288
rect 96212 95276 96218 95328
rect 1104 95226 98808 95248
rect 1104 95174 19606 95226
rect 19658 95174 19670 95226
rect 19722 95174 19734 95226
rect 19786 95174 19798 95226
rect 19850 95174 50326 95226
rect 50378 95174 50390 95226
rect 50442 95174 50454 95226
rect 50506 95174 50518 95226
rect 50570 95174 81046 95226
rect 81098 95174 81110 95226
rect 81162 95174 81174 95226
rect 81226 95174 81238 95226
rect 81290 95174 98808 95226
rect 1104 95152 98808 95174
rect 2240 95084 45554 95112
rect 2240 94985 2268 95084
rect 15105 95047 15163 95053
rect 15105 95013 15117 95047
rect 15151 95044 15163 95047
rect 42242 95044 42248 95056
rect 15151 95016 42248 95044
rect 15151 95013 15163 95016
rect 15105 95007 15163 95013
rect 42242 95004 42248 95016
rect 42300 95004 42306 95056
rect 2225 94979 2283 94985
rect 2225 94945 2237 94979
rect 2271 94945 2283 94979
rect 2225 94939 2283 94945
rect 2409 94979 2467 94985
rect 2409 94945 2421 94979
rect 2455 94945 2467 94979
rect 2409 94939 2467 94945
rect 2501 94979 2559 94985
rect 2501 94945 2513 94979
rect 2547 94976 2559 94979
rect 2590 94976 2596 94988
rect 2547 94948 2596 94976
rect 2547 94945 2559 94948
rect 2501 94939 2559 94945
rect 2424 94908 2452 94939
rect 2590 94936 2596 94948
rect 2648 94936 2654 94988
rect 5077 94979 5135 94985
rect 5077 94945 5089 94979
rect 5123 94976 5135 94979
rect 5442 94976 5448 94988
rect 5123 94948 5448 94976
rect 5123 94945 5135 94948
rect 5077 94939 5135 94945
rect 5442 94936 5448 94948
rect 5500 94936 5506 94988
rect 14918 94976 14924 94988
rect 14879 94948 14924 94976
rect 14918 94936 14924 94948
rect 14976 94936 14982 94988
rect 15378 94985 15384 94988
rect 15197 94979 15255 94985
rect 15197 94945 15209 94979
rect 15243 94945 15255 94979
rect 15197 94939 15255 94945
rect 15341 94979 15384 94985
rect 15341 94945 15353 94979
rect 15341 94939 15384 94945
rect 9858 94908 9864 94920
rect 2424 94880 9864 94908
rect 9858 94868 9864 94880
rect 9916 94868 9922 94920
rect 15212 94908 15240 94939
rect 15378 94936 15384 94939
rect 15436 94936 15442 94988
rect 45526 94976 45554 95084
rect 54113 94979 54171 94985
rect 54113 94976 54125 94979
rect 45526 94948 54125 94976
rect 54113 94945 54125 94948
rect 54159 94945 54171 94979
rect 54113 94939 54171 94945
rect 54481 94979 54539 94985
rect 54481 94945 54493 94979
rect 54527 94976 54539 94979
rect 55398 94976 55404 94988
rect 54527 94948 55404 94976
rect 54527 94945 54539 94948
rect 54481 94939 54539 94945
rect 38746 94908 38752 94920
rect 15212 94880 38752 94908
rect 38746 94868 38752 94880
rect 38804 94868 38810 94920
rect 1857 94843 1915 94849
rect 1857 94809 1869 94843
rect 1903 94840 1915 94843
rect 2590 94840 2596 94852
rect 1903 94812 2596 94840
rect 1903 94809 1915 94812
rect 1857 94803 1915 94809
rect 2590 94800 2596 94812
rect 2648 94800 2654 94852
rect 53926 94840 53932 94852
rect 53887 94812 53932 94840
rect 53926 94800 53932 94812
rect 53984 94800 53990 94852
rect 54128 94840 54156 94939
rect 55398 94936 55404 94948
rect 55456 94976 55462 94988
rect 56410 94976 56416 94988
rect 55456 94948 56416 94976
rect 55456 94936 55462 94948
rect 56410 94936 56416 94948
rect 56468 94936 56474 94988
rect 54570 94908 54576 94920
rect 54531 94880 54576 94908
rect 54570 94868 54576 94880
rect 54628 94868 54634 94920
rect 66070 94840 66076 94852
rect 54128 94812 66076 94840
rect 66070 94800 66076 94812
rect 66128 94800 66134 94852
rect 2038 94772 2044 94784
rect 1999 94744 2044 94772
rect 2038 94732 2044 94744
rect 2096 94732 2102 94784
rect 5166 94772 5172 94784
rect 5127 94744 5172 94772
rect 5166 94732 5172 94744
rect 5224 94732 5230 94784
rect 15470 94772 15476 94784
rect 15431 94744 15476 94772
rect 15470 94732 15476 94744
rect 15528 94732 15534 94784
rect 1104 94682 98808 94704
rect 1104 94630 4246 94682
rect 4298 94630 4310 94682
rect 4362 94630 4374 94682
rect 4426 94630 4438 94682
rect 4490 94630 34966 94682
rect 35018 94630 35030 94682
rect 35082 94630 35094 94682
rect 35146 94630 35158 94682
rect 35210 94630 65686 94682
rect 65738 94630 65750 94682
rect 65802 94630 65814 94682
rect 65866 94630 65878 94682
rect 65930 94630 96406 94682
rect 96458 94630 96470 94682
rect 96522 94630 96534 94682
rect 96586 94630 96598 94682
rect 96650 94630 98808 94682
rect 1104 94608 98808 94630
rect 2590 94528 2596 94580
rect 2648 94568 2654 94580
rect 62761 94571 62819 94577
rect 62761 94568 62773 94571
rect 2648 94540 62773 94568
rect 2648 94528 2654 94540
rect 62761 94537 62773 94540
rect 62807 94537 62819 94571
rect 62761 94531 62819 94537
rect 62776 94432 62804 94531
rect 66162 94432 66168 94444
rect 62776 94404 66168 94432
rect 25501 94367 25559 94373
rect 25501 94333 25513 94367
rect 25547 94364 25559 94367
rect 25777 94367 25835 94373
rect 25777 94364 25789 94367
rect 25547 94336 25789 94364
rect 25547 94333 25559 94336
rect 25501 94327 25559 94333
rect 25777 94333 25789 94336
rect 25823 94364 25835 94367
rect 25866 94364 25872 94376
rect 25823 94336 25872 94364
rect 25823 94333 25835 94336
rect 25777 94327 25835 94333
rect 25866 94324 25872 94336
rect 25924 94324 25930 94376
rect 41601 94367 41659 94373
rect 41601 94333 41613 94367
rect 41647 94364 41659 94367
rect 41874 94364 41880 94376
rect 41647 94336 41880 94364
rect 41647 94333 41659 94336
rect 41601 94327 41659 94333
rect 41874 94324 41880 94336
rect 41932 94324 41938 94376
rect 54573 94367 54631 94373
rect 54573 94333 54585 94367
rect 54619 94333 54631 94367
rect 62776 94364 62804 94404
rect 66162 94392 66168 94404
rect 66220 94392 66226 94444
rect 62945 94367 63003 94373
rect 62945 94364 62957 94367
rect 62776 94336 62957 94364
rect 54573 94327 54631 94333
rect 62945 94333 62957 94336
rect 62991 94333 63003 94367
rect 63218 94364 63224 94376
rect 63179 94336 63224 94364
rect 62945 94327 63003 94333
rect 54389 94299 54447 94305
rect 54389 94296 54401 94299
rect 25516 94268 54401 94296
rect 25516 94240 25544 94268
rect 54389 94265 54401 94268
rect 54435 94296 54447 94299
rect 54588 94296 54616 94327
rect 63218 94324 63224 94336
rect 63276 94324 63282 94376
rect 63402 94296 63408 94308
rect 54435 94268 54616 94296
rect 63363 94268 63408 94296
rect 54435 94265 54447 94268
rect 54389 94259 54447 94265
rect 63402 94256 63408 94268
rect 63460 94256 63466 94308
rect 25498 94188 25504 94240
rect 25556 94188 25562 94240
rect 63034 94228 63040 94240
rect 62947 94200 63040 94228
rect 63034 94188 63040 94200
rect 63092 94228 63098 94240
rect 71866 94228 71872 94240
rect 63092 94200 71872 94228
rect 63092 94188 63098 94200
rect 71866 94188 71872 94200
rect 71924 94228 71930 94240
rect 72418 94228 72424 94240
rect 71924 94200 72424 94228
rect 71924 94188 71930 94200
rect 72418 94188 72424 94200
rect 72476 94188 72482 94240
rect 1104 94138 98808 94160
rect 1104 94086 19606 94138
rect 19658 94086 19670 94138
rect 19722 94086 19734 94138
rect 19786 94086 19798 94138
rect 19850 94086 50326 94138
rect 50378 94086 50390 94138
rect 50442 94086 50454 94138
rect 50506 94086 50518 94138
rect 50570 94086 81046 94138
rect 81098 94086 81110 94138
rect 81162 94086 81174 94138
rect 81226 94086 81238 94138
rect 81290 94086 98808 94138
rect 1104 94064 98808 94086
rect 83826 93984 83832 94036
rect 83884 94024 83890 94036
rect 83884 93996 95832 94024
rect 83884 93984 83890 93996
rect 49878 93916 49884 93968
rect 49936 93956 49942 93968
rect 95602 93956 95608 93968
rect 49936 93928 95608 93956
rect 49936 93916 49942 93928
rect 95602 93916 95608 93928
rect 95660 93916 95666 93968
rect 95701 93959 95759 93965
rect 95701 93925 95713 93959
rect 95747 93956 95759 93959
rect 95804 93956 95832 93996
rect 95747 93928 95832 93956
rect 95747 93925 95759 93928
rect 95701 93919 95759 93925
rect 44818 93848 44824 93900
rect 44876 93888 44882 93900
rect 45462 93888 45468 93900
rect 44876 93860 45468 93888
rect 44876 93848 44882 93860
rect 45462 93848 45468 93860
rect 45520 93888 45526 93900
rect 95513 93891 95571 93897
rect 95513 93888 95525 93891
rect 45520 93860 95525 93888
rect 45520 93848 45526 93860
rect 95513 93857 95525 93860
rect 95559 93888 95571 93891
rect 95789 93891 95847 93897
rect 95789 93888 95801 93891
rect 95559 93860 95801 93888
rect 95559 93857 95571 93860
rect 95513 93851 95571 93857
rect 95789 93857 95801 93860
rect 95835 93857 95847 93891
rect 95970 93888 95976 93900
rect 95931 93860 95976 93888
rect 95789 93851 95847 93857
rect 95970 93848 95976 93860
rect 96028 93848 96034 93900
rect 10686 93780 10692 93832
rect 10744 93820 10750 93832
rect 69290 93820 69296 93832
rect 10744 93792 69296 93820
rect 10744 93780 10750 93792
rect 69290 93780 69296 93792
rect 69348 93780 69354 93832
rect 40494 93712 40500 93764
rect 40552 93752 40558 93764
rect 83458 93752 83464 93764
rect 40552 93724 83464 93752
rect 40552 93712 40558 93724
rect 83458 93712 83464 93724
rect 83516 93712 83522 93764
rect 95602 93644 95608 93696
rect 95660 93684 95666 93696
rect 96157 93687 96215 93693
rect 96157 93684 96169 93687
rect 95660 93656 96169 93684
rect 95660 93644 95666 93656
rect 96157 93653 96169 93656
rect 96203 93653 96215 93687
rect 96157 93647 96215 93653
rect 1104 93594 98808 93616
rect 1104 93542 4246 93594
rect 4298 93542 4310 93594
rect 4362 93542 4374 93594
rect 4426 93542 4438 93594
rect 4490 93542 34966 93594
rect 35018 93542 35030 93594
rect 35082 93542 35094 93594
rect 35146 93542 35158 93594
rect 35210 93542 65686 93594
rect 65738 93542 65750 93594
rect 65802 93542 65814 93594
rect 65866 93542 65878 93594
rect 65930 93542 96406 93594
rect 96458 93542 96470 93594
rect 96522 93542 96534 93594
rect 96586 93542 96598 93594
rect 96650 93542 98808 93594
rect 1104 93520 98808 93542
rect 9858 93304 9864 93356
rect 9916 93344 9922 93356
rect 10686 93344 10692 93356
rect 9916 93316 10692 93344
rect 9916 93304 9922 93316
rect 10686 93304 10692 93316
rect 10744 93304 10750 93356
rect 58066 93236 58072 93288
rect 58124 93276 58130 93288
rect 74442 93276 74448 93288
rect 58124 93248 74448 93276
rect 58124 93236 58130 93248
rect 74442 93236 74448 93248
rect 74500 93236 74506 93288
rect 34514 93168 34520 93220
rect 34572 93208 34578 93220
rect 35342 93208 35348 93220
rect 34572 93180 35348 93208
rect 34572 93168 34578 93180
rect 35342 93168 35348 93180
rect 35400 93208 35406 93220
rect 59538 93208 59544 93220
rect 35400 93180 59544 93208
rect 35400 93168 35406 93180
rect 59538 93168 59544 93180
rect 59596 93168 59602 93220
rect 11698 93100 11704 93152
rect 11756 93140 11762 93152
rect 40494 93140 40500 93152
rect 11756 93112 40500 93140
rect 11756 93100 11762 93112
rect 40494 93100 40500 93112
rect 40552 93100 40558 93152
rect 69290 93100 69296 93152
rect 69348 93140 69354 93152
rect 85850 93140 85856 93152
rect 69348 93112 85856 93140
rect 69348 93100 69354 93112
rect 85850 93100 85856 93112
rect 85908 93100 85914 93152
rect 1104 93050 98808 93072
rect 1104 92998 19606 93050
rect 19658 92998 19670 93050
rect 19722 92998 19734 93050
rect 19786 92998 19798 93050
rect 19850 92998 50326 93050
rect 50378 92998 50390 93050
rect 50442 92998 50454 93050
rect 50506 92998 50518 93050
rect 50570 92998 81046 93050
rect 81098 92998 81110 93050
rect 81162 92998 81174 93050
rect 81226 92998 81238 93050
rect 81290 92998 98808 93050
rect 1104 92976 98808 92998
rect 59538 92556 59544 92608
rect 59596 92596 59602 92608
rect 60550 92596 60556 92608
rect 59596 92568 60556 92596
rect 59596 92556 59602 92568
rect 60550 92556 60556 92568
rect 60608 92556 60614 92608
rect 1104 92506 98808 92528
rect 1104 92454 4246 92506
rect 4298 92454 4310 92506
rect 4362 92454 4374 92506
rect 4426 92454 4438 92506
rect 4490 92454 34966 92506
rect 35018 92454 35030 92506
rect 35082 92454 35094 92506
rect 35146 92454 35158 92506
rect 35210 92454 65686 92506
rect 65738 92454 65750 92506
rect 65802 92454 65814 92506
rect 65866 92454 65878 92506
rect 65930 92454 96406 92506
rect 96458 92454 96470 92506
rect 96522 92454 96534 92506
rect 96586 92454 96598 92506
rect 96650 92454 98808 92506
rect 1104 92432 98808 92454
rect 68922 92284 68928 92336
rect 68980 92324 68986 92336
rect 92569 92327 92627 92333
rect 92569 92324 92581 92327
rect 68980 92296 92581 92324
rect 68980 92284 68986 92296
rect 92569 92293 92581 92296
rect 92615 92293 92627 92327
rect 93762 92324 93768 92336
rect 93723 92296 93768 92324
rect 92569 92287 92627 92293
rect 93762 92284 93768 92296
rect 93820 92284 93826 92336
rect 92658 92256 92664 92268
rect 92619 92228 92664 92256
rect 92658 92216 92664 92228
rect 92716 92216 92722 92268
rect 93854 92256 93860 92268
rect 93815 92228 93860 92256
rect 93854 92216 93860 92228
rect 93912 92216 93918 92268
rect 36354 92188 36360 92200
rect 36315 92160 36360 92188
rect 36354 92148 36360 92160
rect 36412 92148 36418 92200
rect 92474 92197 92480 92200
rect 92440 92191 92480 92197
rect 92440 92157 92452 92191
rect 92440 92151 92480 92157
rect 92474 92148 92480 92151
rect 92532 92148 92538 92200
rect 93670 92197 93676 92200
rect 93636 92191 93676 92197
rect 93636 92157 93648 92191
rect 93636 92151 93676 92157
rect 93670 92148 93676 92151
rect 93728 92148 93734 92200
rect 23474 92120 23480 92132
rect 23435 92092 23480 92120
rect 23474 92080 23480 92092
rect 23532 92080 23538 92132
rect 23658 92120 23664 92132
rect 23619 92092 23664 92120
rect 23658 92080 23664 92092
rect 23716 92080 23722 92132
rect 35434 92080 35440 92132
rect 35492 92120 35498 92132
rect 36265 92123 36323 92129
rect 36265 92120 36277 92123
rect 35492 92092 36277 92120
rect 35492 92080 35498 92092
rect 36265 92089 36277 92092
rect 36311 92089 36323 92123
rect 36265 92083 36323 92089
rect 92198 92080 92204 92132
rect 92256 92120 92262 92132
rect 92293 92123 92351 92129
rect 92293 92120 92305 92123
rect 92256 92092 92305 92120
rect 92256 92080 92262 92092
rect 92293 92089 92305 92092
rect 92339 92089 92351 92123
rect 93486 92120 93492 92132
rect 93447 92092 93492 92120
rect 92293 92083 92351 92089
rect 93486 92080 93492 92092
rect 93544 92080 93550 92132
rect 84286 92012 84292 92064
rect 84344 92052 84350 92064
rect 92937 92055 92995 92061
rect 92937 92052 92949 92055
rect 84344 92024 92949 92052
rect 84344 92012 84350 92024
rect 92937 92021 92949 92024
rect 92983 92021 92995 92055
rect 94130 92052 94136 92064
rect 94091 92024 94136 92052
rect 92937 92015 92995 92021
rect 94130 92012 94136 92024
rect 94188 92012 94194 92064
rect 1104 91962 98808 91984
rect 1104 91910 19606 91962
rect 19658 91910 19670 91962
rect 19722 91910 19734 91962
rect 19786 91910 19798 91962
rect 19850 91910 50326 91962
rect 50378 91910 50390 91962
rect 50442 91910 50454 91962
rect 50506 91910 50518 91962
rect 50570 91910 81046 91962
rect 81098 91910 81110 91962
rect 81162 91910 81174 91962
rect 81226 91910 81238 91962
rect 81290 91910 98808 91962
rect 1104 91888 98808 91910
rect 49050 91848 49056 91860
rect 47320 91820 49056 91848
rect 11790 91740 11796 91792
rect 11848 91780 11854 91792
rect 46474 91780 46480 91792
rect 11848 91752 46480 91780
rect 11848 91740 11854 91752
rect 46474 91740 46480 91752
rect 46532 91740 46538 91792
rect 47320 91721 47348 91820
rect 49050 91808 49056 91820
rect 49108 91808 49114 91860
rect 65242 91808 65248 91860
rect 65300 91848 65306 91860
rect 65300 91820 73936 91848
rect 65300 91808 65306 91820
rect 48958 91780 48964 91792
rect 47412 91752 47624 91780
rect 47305 91715 47363 91721
rect 47305 91681 47317 91715
rect 47351 91681 47363 91715
rect 47305 91675 47363 91681
rect 27062 91604 27068 91656
rect 27120 91644 27126 91656
rect 47412 91644 47440 91752
rect 47596 91721 47624 91752
rect 47688 91752 48964 91780
rect 47688 91721 47716 91752
rect 48958 91740 48964 91752
rect 49016 91740 49022 91792
rect 47488 91715 47546 91721
rect 47488 91681 47500 91715
rect 47534 91681 47546 91715
rect 47488 91675 47546 91681
rect 47578 91715 47636 91721
rect 47578 91681 47590 91715
rect 47624 91681 47636 91715
rect 47578 91675 47636 91681
rect 47673 91715 47731 91721
rect 47673 91681 47685 91715
rect 47719 91681 47731 91715
rect 47673 91675 47731 91681
rect 47857 91715 47915 91721
rect 47857 91681 47869 91715
rect 47903 91712 47915 91715
rect 68462 91712 68468 91724
rect 47903 91684 68468 91712
rect 47903 91681 47915 91684
rect 47857 91675 47915 91681
rect 27120 91616 47440 91644
rect 47504 91644 47532 91675
rect 68462 91672 68468 91684
rect 68520 91712 68526 91724
rect 68922 91712 68928 91724
rect 68520 91684 68928 91712
rect 68520 91672 68526 91684
rect 68922 91672 68928 91684
rect 68980 91672 68986 91724
rect 73614 91712 73620 91724
rect 73575 91684 73620 91712
rect 73614 91672 73620 91684
rect 73672 91672 73678 91724
rect 73908 91721 73936 91820
rect 73800 91715 73858 91721
rect 73800 91681 73812 91715
rect 73846 91681 73858 91715
rect 73800 91675 73858 91681
rect 73893 91715 73951 91721
rect 73893 91681 73905 91715
rect 73939 91681 73951 91715
rect 74166 91712 74172 91724
rect 74127 91684 74172 91712
rect 73893 91675 73951 91681
rect 47504 91616 55214 91644
rect 27120 91604 27126 91616
rect 55186 91576 55214 91616
rect 61562 91576 61568 91588
rect 22066 91548 50384 91576
rect 55186 91548 61568 91576
rect 14734 91468 14740 91520
rect 14792 91508 14798 91520
rect 22066 91508 22094 91548
rect 47946 91508 47952 91520
rect 14792 91480 22094 91508
rect 47907 91480 47952 91508
rect 14792 91468 14798 91480
rect 47946 91468 47952 91480
rect 48004 91468 48010 91520
rect 50356 91508 50384 91548
rect 61562 91536 61568 91548
rect 61620 91536 61626 91588
rect 73433 91511 73491 91517
rect 73433 91508 73445 91511
rect 50356 91480 73445 91508
rect 73433 91477 73445 91480
rect 73479 91508 73491 91511
rect 73816 91508 73844 91675
rect 74166 91672 74172 91684
rect 74224 91672 74230 91724
rect 73982 91644 73988 91656
rect 73943 91616 73988 91644
rect 73982 91604 73988 91616
rect 74040 91604 74046 91656
rect 74350 91576 74356 91588
rect 74311 91548 74356 91576
rect 74350 91536 74356 91548
rect 74408 91536 74414 91588
rect 73479 91480 73844 91508
rect 73479 91477 73491 91480
rect 73433 91471 73491 91477
rect 1104 91418 98808 91440
rect 1104 91366 4246 91418
rect 4298 91366 4310 91418
rect 4362 91366 4374 91418
rect 4426 91366 4438 91418
rect 4490 91366 34966 91418
rect 35018 91366 35030 91418
rect 35082 91366 35094 91418
rect 35146 91366 35158 91418
rect 35210 91366 65686 91418
rect 65738 91366 65750 91418
rect 65802 91366 65814 91418
rect 65866 91366 65878 91418
rect 65930 91366 96406 91418
rect 96458 91366 96470 91418
rect 96522 91366 96534 91418
rect 96586 91366 96598 91418
rect 96650 91366 98808 91418
rect 1104 91344 98808 91366
rect 68554 91264 68560 91316
rect 68612 91304 68618 91316
rect 73982 91304 73988 91316
rect 68612 91276 73988 91304
rect 68612 91264 68618 91276
rect 73982 91264 73988 91276
rect 74040 91264 74046 91316
rect 52454 91168 52460 91180
rect 44192 91140 52460 91168
rect 44085 91103 44143 91109
rect 44085 91069 44097 91103
rect 44131 91100 44143 91103
rect 44192 91100 44220 91140
rect 52454 91128 52460 91140
rect 52512 91128 52518 91180
rect 55030 91100 55036 91112
rect 44131 91072 44220 91100
rect 44284 91072 55036 91100
rect 44131 91069 44143 91072
rect 44085 91063 44143 91069
rect 44284 90973 44312 91072
rect 55030 91060 55036 91072
rect 55088 91060 55094 91112
rect 61470 91060 61476 91112
rect 61528 91100 61534 91112
rect 97721 91103 97779 91109
rect 97721 91100 97733 91103
rect 61528 91072 97733 91100
rect 61528 91060 61534 91072
rect 97721 91069 97733 91072
rect 97767 91100 97779 91103
rect 97905 91103 97963 91109
rect 97905 91100 97917 91103
rect 97767 91072 97917 91100
rect 97767 91069 97779 91072
rect 97721 91063 97779 91069
rect 97905 91069 97917 91072
rect 97951 91069 97963 91103
rect 97905 91063 97963 91069
rect 44269 90967 44327 90973
rect 44269 90933 44281 90967
rect 44315 90933 44327 90967
rect 44269 90927 44327 90933
rect 1104 90874 98808 90896
rect 1104 90822 19606 90874
rect 19658 90822 19670 90874
rect 19722 90822 19734 90874
rect 19786 90822 19798 90874
rect 19850 90822 50326 90874
rect 50378 90822 50390 90874
rect 50442 90822 50454 90874
rect 50506 90822 50518 90874
rect 50570 90822 81046 90874
rect 81098 90822 81110 90874
rect 81162 90822 81174 90874
rect 81226 90822 81238 90874
rect 81290 90822 98808 90874
rect 1104 90800 98808 90822
rect 8294 90584 8300 90636
rect 8352 90624 8358 90636
rect 9493 90627 9551 90633
rect 9493 90624 9505 90627
rect 8352 90596 9505 90624
rect 8352 90584 8358 90596
rect 9493 90593 9505 90596
rect 9539 90593 9551 90627
rect 69842 90624 69848 90636
rect 69803 90596 69848 90624
rect 9493 90587 9551 90593
rect 69842 90584 69848 90596
rect 69900 90584 69906 90636
rect 70302 90556 70308 90568
rect 70263 90528 70308 90556
rect 70302 90516 70308 90528
rect 70360 90516 70366 90568
rect 9674 90420 9680 90432
rect 9635 90392 9680 90420
rect 9674 90380 9680 90392
rect 9732 90380 9738 90432
rect 39390 90380 39396 90432
rect 39448 90420 39454 90432
rect 52273 90423 52331 90429
rect 52273 90420 52285 90423
rect 39448 90392 52285 90420
rect 39448 90380 39454 90392
rect 52273 90389 52285 90392
rect 52319 90420 52331 90423
rect 52457 90423 52515 90429
rect 52457 90420 52469 90423
rect 52319 90392 52469 90420
rect 52319 90389 52331 90392
rect 52273 90383 52331 90389
rect 52457 90389 52469 90392
rect 52503 90389 52515 90423
rect 52457 90383 52515 90389
rect 74350 90380 74356 90432
rect 74408 90420 74414 90432
rect 91738 90420 91744 90432
rect 74408 90392 91744 90420
rect 74408 90380 74414 90392
rect 91738 90380 91744 90392
rect 91796 90380 91802 90432
rect 1104 90330 98808 90352
rect 1104 90278 4246 90330
rect 4298 90278 4310 90330
rect 4362 90278 4374 90330
rect 4426 90278 4438 90330
rect 4490 90278 34966 90330
rect 35018 90278 35030 90330
rect 35082 90278 35094 90330
rect 35146 90278 35158 90330
rect 35210 90278 65686 90330
rect 65738 90278 65750 90330
rect 65802 90278 65814 90330
rect 65866 90278 65878 90330
rect 65930 90278 96406 90330
rect 96458 90278 96470 90330
rect 96522 90278 96534 90330
rect 96586 90278 96598 90330
rect 96650 90278 98808 90330
rect 1104 90256 98808 90278
rect 41046 90216 41052 90228
rect 29564 90188 41052 90216
rect 29564 90089 29592 90188
rect 41046 90176 41052 90188
rect 41104 90176 41110 90228
rect 45281 90151 45339 90157
rect 45281 90117 45293 90151
rect 45327 90148 45339 90151
rect 45327 90120 45554 90148
rect 45327 90117 45339 90120
rect 45281 90111 45339 90117
rect 29549 90083 29607 90089
rect 29549 90049 29561 90083
rect 29595 90049 29607 90083
rect 29549 90043 29607 90049
rect 29641 90083 29699 90089
rect 29641 90049 29653 90083
rect 29687 90080 29699 90083
rect 29687 90052 44036 90080
rect 29687 90049 29699 90052
rect 29641 90043 29699 90049
rect 29270 90012 29276 90024
rect 29231 89984 29276 90012
rect 29270 89972 29276 89984
rect 29328 89972 29334 90024
rect 29454 90012 29460 90024
rect 29415 89984 29460 90012
rect 29454 89972 29460 89984
rect 29512 89972 29518 90024
rect 29825 90015 29883 90021
rect 29825 89981 29837 90015
rect 29871 89981 29883 90015
rect 29825 89975 29883 89981
rect 28258 89904 28264 89956
rect 28316 89944 28322 89956
rect 29840 89944 29868 89975
rect 30282 89972 30288 90024
rect 30340 90012 30346 90024
rect 30469 90015 30527 90021
rect 30469 90012 30481 90015
rect 30340 89984 30481 90012
rect 30340 89972 30346 89984
rect 30469 89981 30481 89984
rect 30515 89981 30527 90015
rect 30742 90012 30748 90024
rect 30703 89984 30748 90012
rect 30469 89975 30527 89981
rect 28316 89916 29868 89944
rect 28316 89904 28322 89916
rect 4062 89836 4068 89888
rect 4120 89876 4126 89888
rect 29917 89879 29975 89885
rect 29917 89876 29929 89879
rect 4120 89848 29929 89876
rect 4120 89836 4126 89848
rect 29917 89845 29929 89848
rect 29963 89845 29975 89879
rect 30484 89876 30512 89975
rect 30742 89972 30748 89984
rect 30800 89972 30806 90024
rect 43901 90015 43959 90021
rect 43901 90012 43913 90015
rect 31726 89984 43913 90012
rect 31726 89876 31754 89984
rect 43901 89981 43913 89984
rect 43947 89981 43959 90015
rect 44008 90012 44036 90052
rect 44450 90012 44456 90024
rect 44008 89984 44456 90012
rect 43901 89975 43959 89981
rect 44450 89972 44456 89984
rect 44508 89972 44514 90024
rect 45526 90012 45554 90120
rect 49970 90108 49976 90160
rect 50028 90148 50034 90160
rect 75089 90151 75147 90157
rect 75089 90148 75101 90151
rect 50028 90120 75101 90148
rect 50028 90108 50034 90120
rect 75089 90117 75101 90120
rect 75135 90117 75147 90151
rect 75089 90111 75147 90117
rect 74721 90083 74779 90089
rect 74721 90049 74733 90083
rect 74767 90080 74779 90083
rect 74905 90083 74963 90089
rect 74905 90080 74917 90083
rect 74767 90052 74917 90080
rect 74767 90049 74779 90052
rect 74721 90043 74779 90049
rect 74905 90049 74917 90052
rect 74951 90080 74963 90083
rect 74951 90052 75500 90080
rect 74951 90049 74963 90052
rect 74905 90043 74963 90049
rect 63034 90012 63040 90024
rect 45526 89984 63040 90012
rect 63034 89972 63040 89984
rect 63092 89972 63098 90024
rect 75270 90021 75276 90024
rect 75268 89975 75276 90021
rect 75328 90012 75334 90024
rect 75472 90021 75500 90052
rect 75457 90015 75515 90021
rect 75328 89984 75368 90012
rect 75270 89972 75276 89975
rect 75328 89972 75334 89984
rect 75457 89981 75469 90015
rect 75503 89981 75515 90015
rect 75457 89975 75515 89981
rect 75641 90015 75699 90021
rect 75641 89981 75653 90015
rect 75687 90012 75699 90015
rect 75822 90012 75828 90024
rect 75687 89984 75828 90012
rect 75687 89981 75699 89984
rect 75641 89975 75699 89981
rect 75822 89972 75828 89984
rect 75880 89972 75886 90024
rect 44174 89953 44180 89956
rect 44168 89907 44180 89953
rect 44232 89944 44238 89956
rect 44232 89916 44268 89944
rect 44174 89904 44180 89907
rect 44232 89904 44238 89916
rect 46842 89904 46848 89956
rect 46900 89944 46906 89956
rect 75365 89947 75423 89953
rect 75365 89944 75377 89947
rect 46900 89916 75377 89944
rect 46900 89904 46906 89916
rect 75365 89913 75377 89916
rect 75411 89944 75423 89947
rect 76190 89944 76196 89956
rect 75411 89916 75592 89944
rect 76151 89916 76196 89944
rect 75411 89913 75423 89916
rect 75365 89907 75423 89913
rect 30484 89848 31754 89876
rect 29917 89839 29975 89845
rect 31938 89836 31944 89888
rect 31996 89876 32002 89888
rect 32033 89879 32091 89885
rect 32033 89876 32045 89879
rect 31996 89848 32045 89876
rect 31996 89836 32002 89848
rect 32033 89845 32045 89848
rect 32079 89845 32091 89879
rect 32033 89839 32091 89845
rect 44910 89836 44916 89888
rect 44968 89876 44974 89888
rect 74721 89879 74779 89885
rect 74721 89876 74733 89879
rect 44968 89848 74733 89876
rect 44968 89836 44974 89848
rect 74721 89845 74733 89848
rect 74767 89845 74779 89879
rect 75564 89876 75592 89916
rect 76190 89904 76196 89916
rect 76248 89904 76254 89956
rect 75730 89876 75736 89888
rect 75564 89848 75736 89876
rect 74721 89839 74779 89845
rect 75730 89836 75736 89848
rect 75788 89836 75794 89888
rect 76282 89876 76288 89888
rect 76243 89848 76288 89876
rect 76282 89836 76288 89848
rect 76340 89836 76346 89888
rect 1104 89786 98808 89808
rect 1104 89734 19606 89786
rect 19658 89734 19670 89786
rect 19722 89734 19734 89786
rect 19786 89734 19798 89786
rect 19850 89734 50326 89786
rect 50378 89734 50390 89786
rect 50442 89734 50454 89786
rect 50506 89734 50518 89786
rect 50570 89734 81046 89786
rect 81098 89734 81110 89786
rect 81162 89734 81174 89786
rect 81226 89734 81238 89786
rect 81290 89734 98808 89786
rect 1104 89712 98808 89734
rect 48958 89564 48964 89616
rect 49016 89604 49022 89616
rect 49016 89576 74580 89604
rect 49016 89564 49022 89576
rect 31110 89496 31116 89548
rect 31168 89536 31174 89548
rect 73798 89536 73804 89548
rect 31168 89508 60734 89536
rect 73759 89508 73804 89536
rect 31168 89496 31174 89508
rect 60706 89468 60734 89508
rect 73798 89496 73804 89508
rect 73856 89496 73862 89548
rect 74552 89545 74580 89576
rect 87966 89564 87972 89616
rect 88024 89604 88030 89616
rect 88150 89604 88156 89616
rect 88024 89576 88156 89604
rect 88024 89564 88030 89576
rect 88150 89564 88156 89576
rect 88208 89604 88214 89616
rect 88208 89576 89208 89604
rect 88208 89564 88214 89576
rect 74169 89539 74227 89545
rect 74169 89536 74181 89539
rect 73908 89508 74181 89536
rect 73908 89468 73936 89508
rect 74169 89505 74181 89508
rect 74215 89505 74227 89539
rect 74169 89499 74227 89505
rect 74537 89539 74595 89545
rect 74537 89505 74549 89539
rect 74583 89505 74595 89539
rect 74537 89499 74595 89505
rect 81434 89496 81440 89548
rect 81492 89536 81498 89548
rect 89180 89545 89208 89576
rect 88797 89539 88855 89545
rect 88797 89536 88809 89539
rect 81492 89508 88809 89536
rect 81492 89496 81498 89508
rect 88797 89505 88809 89508
rect 88843 89505 88855 89539
rect 88797 89499 88855 89505
rect 89165 89539 89223 89545
rect 89165 89505 89177 89539
rect 89211 89505 89223 89539
rect 89165 89499 89223 89505
rect 60706 89440 73936 89468
rect 73985 89471 74043 89477
rect 73985 89437 73997 89471
rect 74031 89437 74043 89471
rect 74626 89468 74632 89480
rect 74587 89440 74632 89468
rect 73985 89431 74043 89437
rect 70762 89360 70768 89412
rect 70820 89400 70826 89412
rect 74000 89400 74028 89431
rect 74626 89428 74632 89440
rect 74684 89428 74690 89480
rect 88242 89468 88248 89480
rect 88203 89440 88248 89468
rect 88242 89428 88248 89440
rect 88300 89428 88306 89480
rect 88610 89468 88616 89480
rect 88571 89440 88616 89468
rect 88610 89428 88616 89440
rect 88668 89428 88674 89480
rect 89073 89471 89131 89477
rect 89073 89437 89085 89471
rect 89119 89437 89131 89471
rect 89073 89431 89131 89437
rect 74902 89400 74908 89412
rect 70820 89372 74028 89400
rect 74863 89372 74908 89400
rect 70820 89360 70826 89372
rect 74902 89360 74908 89372
rect 74960 89360 74966 89412
rect 52454 89292 52460 89344
rect 52512 89332 52518 89344
rect 53190 89332 53196 89344
rect 52512 89304 53196 89332
rect 52512 89292 52518 89304
rect 53190 89292 53196 89304
rect 53248 89332 53254 89344
rect 89088 89332 89116 89431
rect 53248 89304 89116 89332
rect 53248 89292 53254 89304
rect 1104 89242 98808 89264
rect 1104 89190 4246 89242
rect 4298 89190 4310 89242
rect 4362 89190 4374 89242
rect 4426 89190 4438 89242
rect 4490 89190 34966 89242
rect 35018 89190 35030 89242
rect 35082 89190 35094 89242
rect 35146 89190 35158 89242
rect 35210 89190 65686 89242
rect 65738 89190 65750 89242
rect 65802 89190 65814 89242
rect 65866 89190 65878 89242
rect 65930 89190 96406 89242
rect 96458 89190 96470 89242
rect 96522 89190 96534 89242
rect 96586 89190 96598 89242
rect 96650 89190 98808 89242
rect 1104 89168 98808 89190
rect 8297 89131 8355 89137
rect 8297 89097 8309 89131
rect 8343 89128 8355 89131
rect 53742 89128 53748 89140
rect 8343 89100 53748 89128
rect 8343 89097 8355 89100
rect 8297 89091 8355 89097
rect 53742 89088 53748 89100
rect 53800 89128 53806 89140
rect 53800 89100 55214 89128
rect 53800 89088 53806 89100
rect 3881 89063 3939 89069
rect 3881 89029 3893 89063
rect 3927 89060 3939 89063
rect 5074 89060 5080 89072
rect 3927 89032 5080 89060
rect 3927 89029 3939 89032
rect 3881 89023 3939 89029
rect 5074 89020 5080 89032
rect 5132 89060 5138 89072
rect 5132 89032 16574 89060
rect 5132 89020 5138 89032
rect 6733 88995 6791 89001
rect 6733 88961 6745 88995
rect 6779 88992 6791 88995
rect 8297 88995 8355 89001
rect 8297 88992 8309 88995
rect 6779 88964 8309 88992
rect 6779 88961 6791 88964
rect 6733 88955 6791 88961
rect 2501 88927 2559 88933
rect 2501 88893 2513 88927
rect 2547 88924 2559 88927
rect 2590 88924 2596 88936
rect 2547 88896 2596 88924
rect 2547 88893 2559 88896
rect 2501 88887 2559 88893
rect 2590 88884 2596 88896
rect 2648 88884 2654 88936
rect 2768 88927 2826 88933
rect 2768 88893 2780 88927
rect 2814 88924 2826 88927
rect 4062 88924 4068 88936
rect 2814 88896 4068 88924
rect 2814 88893 2826 88896
rect 2768 88887 2826 88893
rect 4062 88884 4068 88896
rect 4120 88884 4126 88936
rect 7285 88927 7343 88933
rect 7285 88924 7297 88927
rect 7116 88896 7297 88924
rect 6914 88788 6920 88800
rect 6875 88760 6920 88788
rect 6914 88748 6920 88760
rect 6972 88748 6978 88800
rect 7116 88788 7144 88896
rect 7285 88893 7297 88896
rect 7331 88893 7343 88927
rect 7558 88924 7564 88936
rect 7519 88896 7564 88924
rect 7285 88887 7343 88893
rect 7558 88884 7564 88896
rect 7616 88884 7622 88936
rect 7653 88927 7711 88933
rect 7653 88893 7665 88927
rect 7699 88924 7711 88927
rect 7742 88924 7748 88936
rect 7699 88896 7748 88924
rect 7699 88893 7711 88896
rect 7653 88887 7711 88893
rect 7742 88884 7748 88896
rect 7800 88884 7806 88936
rect 7944 88933 7972 88964
rect 8297 88961 8309 88964
rect 8343 88961 8355 88995
rect 16546 88992 16574 89032
rect 28166 88992 28172 89004
rect 16546 88964 28172 88992
rect 8297 88955 8355 88961
rect 28166 88952 28172 88964
rect 28224 88952 28230 89004
rect 55186 88992 55214 89100
rect 82170 88992 82176 89004
rect 55186 88964 82176 88992
rect 82170 88952 82176 88964
rect 82228 88952 82234 89004
rect 7929 88927 7987 88933
rect 7929 88893 7941 88927
rect 7975 88893 7987 88927
rect 7929 88887 7987 88893
rect 8205 88927 8263 88933
rect 8205 88893 8217 88927
rect 8251 88924 8263 88927
rect 16298 88924 16304 88936
rect 8251 88896 16304 88924
rect 8251 88893 8263 88896
rect 8205 88887 8263 88893
rect 16298 88884 16304 88896
rect 16356 88884 16362 88936
rect 17681 88927 17739 88933
rect 17681 88924 17693 88927
rect 16546 88896 17693 88924
rect 13814 88816 13820 88868
rect 13872 88856 13878 88868
rect 15102 88856 15108 88868
rect 13872 88828 15108 88856
rect 13872 88816 13878 88828
rect 15102 88816 15108 88828
rect 15160 88856 15166 88868
rect 16546 88856 16574 88896
rect 17681 88893 17693 88896
rect 17727 88893 17739 88927
rect 17954 88924 17960 88936
rect 17915 88896 17960 88924
rect 17681 88887 17739 88893
rect 17954 88884 17960 88896
rect 18012 88884 18018 88936
rect 55030 88924 55036 88936
rect 54991 88896 55036 88924
rect 55030 88884 55036 88896
rect 55088 88884 55094 88936
rect 55861 88859 55919 88865
rect 15160 88828 16574 88856
rect 18892 88828 26234 88856
rect 15160 88816 15166 88828
rect 18892 88788 18920 88828
rect 19058 88788 19064 88800
rect 7116 88760 18920 88788
rect 19019 88760 19064 88788
rect 19058 88748 19064 88760
rect 19116 88748 19122 88800
rect 26206 88788 26234 88828
rect 55861 88825 55873 88859
rect 55907 88856 55919 88859
rect 71130 88856 71136 88868
rect 55907 88828 71136 88856
rect 55907 88825 55919 88828
rect 55861 88819 55919 88825
rect 71130 88816 71136 88828
rect 71188 88816 71194 88868
rect 50062 88788 50068 88800
rect 26206 88760 50068 88788
rect 50062 88748 50068 88760
rect 50120 88748 50126 88800
rect 1104 88698 98808 88720
rect 1104 88646 19606 88698
rect 19658 88646 19670 88698
rect 19722 88646 19734 88698
rect 19786 88646 19798 88698
rect 19850 88646 50326 88698
rect 50378 88646 50390 88698
rect 50442 88646 50454 88698
rect 50506 88646 50518 88698
rect 50570 88646 81046 88698
rect 81098 88646 81110 88698
rect 81162 88646 81174 88698
rect 81226 88646 81238 88698
rect 81290 88646 98808 88698
rect 1104 88624 98808 88646
rect 16025 88587 16083 88593
rect 16025 88553 16037 88587
rect 16071 88584 16083 88587
rect 16114 88584 16120 88596
rect 16071 88556 16120 88584
rect 16071 88553 16083 88556
rect 16025 88547 16083 88553
rect 16114 88544 16120 88556
rect 16172 88544 16178 88596
rect 16298 88544 16304 88596
rect 16356 88584 16362 88596
rect 49694 88584 49700 88596
rect 16356 88556 49700 88584
rect 16356 88544 16362 88556
rect 49694 88544 49700 88556
rect 49752 88544 49758 88596
rect 7742 88476 7748 88528
rect 7800 88516 7806 88528
rect 43806 88516 43812 88528
rect 7800 88488 43812 88516
rect 7800 88476 7806 88488
rect 43806 88476 43812 88488
rect 43864 88476 43870 88528
rect 2590 88408 2596 88460
rect 2648 88448 2654 88460
rect 13814 88448 13820 88460
rect 2648 88420 13820 88448
rect 2648 88408 2654 88420
rect 13814 88408 13820 88420
rect 13872 88408 13878 88460
rect 15838 88448 15844 88460
rect 15799 88420 15844 88448
rect 15838 88408 15844 88420
rect 15896 88408 15902 88460
rect 67269 88383 67327 88389
rect 67269 88349 67281 88383
rect 67315 88380 67327 88383
rect 67545 88383 67603 88389
rect 67545 88380 67557 88383
rect 67315 88352 67557 88380
rect 67315 88349 67327 88352
rect 67269 88343 67327 88349
rect 67545 88349 67557 88352
rect 67591 88380 67603 88383
rect 68278 88380 68284 88392
rect 67591 88352 68284 88380
rect 67591 88349 67603 88352
rect 67545 88343 67603 88349
rect 68278 88340 68284 88352
rect 68336 88340 68342 88392
rect 77478 88204 77484 88256
rect 77536 88244 77542 88256
rect 83826 88244 83832 88256
rect 77536 88216 83832 88244
rect 77536 88204 77542 88216
rect 83826 88204 83832 88216
rect 83884 88204 83890 88256
rect 1104 88154 98808 88176
rect 1104 88102 4246 88154
rect 4298 88102 4310 88154
rect 4362 88102 4374 88154
rect 4426 88102 4438 88154
rect 4490 88102 34966 88154
rect 35018 88102 35030 88154
rect 35082 88102 35094 88154
rect 35146 88102 35158 88154
rect 35210 88102 65686 88154
rect 65738 88102 65750 88154
rect 65802 88102 65814 88154
rect 65866 88102 65878 88154
rect 65930 88102 96406 88154
rect 96458 88102 96470 88154
rect 96522 88102 96534 88154
rect 96586 88102 96598 88154
rect 96650 88102 98808 88154
rect 1104 88080 98808 88102
rect 41046 88000 41052 88052
rect 41104 88040 41110 88052
rect 90266 88040 90272 88052
rect 41104 88012 90272 88040
rect 41104 88000 41110 88012
rect 90266 88000 90272 88012
rect 90324 88000 90330 88052
rect 77573 87975 77631 87981
rect 77573 87941 77585 87975
rect 77619 87972 77631 87975
rect 77662 87972 77668 87984
rect 77619 87944 77668 87972
rect 77619 87941 77631 87944
rect 77573 87935 77631 87941
rect 77662 87932 77668 87944
rect 77720 87932 77726 87984
rect 32490 87864 32496 87916
rect 32548 87904 32554 87916
rect 89622 87904 89628 87916
rect 32548 87876 89628 87904
rect 32548 87864 32554 87876
rect 89622 87864 89628 87876
rect 89680 87864 89686 87916
rect 8294 87836 8300 87848
rect 8255 87808 8300 87836
rect 8294 87796 8300 87808
rect 8352 87796 8358 87848
rect 8573 87839 8631 87845
rect 8573 87805 8585 87839
rect 8619 87836 8631 87839
rect 15657 87839 15715 87845
rect 15657 87836 15669 87839
rect 8619 87808 15669 87836
rect 8619 87805 8631 87808
rect 8573 87799 8631 87805
rect 15657 87805 15669 87808
rect 15703 87836 15715 87839
rect 77478 87836 77484 87848
rect 15703 87808 77484 87836
rect 15703 87805 15715 87808
rect 15657 87799 15715 87805
rect 77478 87796 77484 87808
rect 77536 87796 77542 87848
rect 77570 87796 77576 87848
rect 77628 87836 77634 87848
rect 77665 87839 77723 87845
rect 77665 87836 77677 87839
rect 77628 87808 77677 87836
rect 77628 87796 77634 87808
rect 77665 87805 77677 87808
rect 77711 87805 77723 87839
rect 77665 87799 77723 87805
rect 77754 87796 77760 87848
rect 77812 87836 77818 87848
rect 77941 87839 77999 87845
rect 77941 87836 77953 87839
rect 77812 87808 77953 87836
rect 77812 87796 77818 87808
rect 77941 87805 77953 87808
rect 77987 87805 77999 87839
rect 77941 87799 77999 87805
rect 15746 87728 15752 87780
rect 15804 87768 15810 87780
rect 15933 87771 15991 87777
rect 15933 87768 15945 87771
rect 15804 87740 15945 87768
rect 15804 87728 15810 87740
rect 15933 87737 15945 87740
rect 15979 87737 15991 87771
rect 15933 87731 15991 87737
rect 22094 87728 22100 87780
rect 22152 87768 22158 87780
rect 23382 87768 23388 87780
rect 22152 87740 23388 87768
rect 22152 87728 22158 87740
rect 23382 87728 23388 87740
rect 23440 87768 23446 87780
rect 34790 87768 34796 87780
rect 23440 87740 34796 87768
rect 23440 87728 23446 87740
rect 34790 87728 34796 87740
rect 34848 87728 34854 87780
rect 69750 87728 69756 87780
rect 69808 87768 69814 87780
rect 69808 87740 77616 87768
rect 69808 87728 69814 87740
rect 29270 87660 29276 87712
rect 29328 87700 29334 87712
rect 54478 87700 54484 87712
rect 29328 87672 54484 87700
rect 29328 87660 29334 87672
rect 54478 87660 54484 87672
rect 54536 87660 54542 87712
rect 77588 87700 77616 87740
rect 79045 87703 79103 87709
rect 79045 87700 79057 87703
rect 77588 87672 79057 87700
rect 79045 87669 79057 87672
rect 79091 87669 79103 87703
rect 79045 87663 79103 87669
rect 1104 87610 98808 87632
rect 1104 87558 19606 87610
rect 19658 87558 19670 87610
rect 19722 87558 19734 87610
rect 19786 87558 19798 87610
rect 19850 87558 50326 87610
rect 50378 87558 50390 87610
rect 50442 87558 50454 87610
rect 50506 87558 50518 87610
rect 50570 87558 81046 87610
rect 81098 87558 81110 87610
rect 81162 87558 81174 87610
rect 81226 87558 81238 87610
rect 81290 87558 98808 87610
rect 1104 87536 98808 87558
rect 2056 87468 12434 87496
rect 2056 87369 2084 87468
rect 10778 87428 10784 87440
rect 2424 87400 10784 87428
rect 2424 87369 2452 87400
rect 10778 87388 10784 87400
rect 10836 87388 10842 87440
rect 12406 87428 12434 87468
rect 77570 87456 77576 87508
rect 77628 87496 77634 87508
rect 84562 87496 84568 87508
rect 77628 87468 84568 87496
rect 77628 87456 77634 87468
rect 84562 87456 84568 87468
rect 84620 87456 84626 87508
rect 89622 87456 89628 87508
rect 89680 87496 89686 87508
rect 89806 87496 89812 87508
rect 89680 87468 89812 87496
rect 89680 87456 89686 87468
rect 89806 87456 89812 87468
rect 89864 87456 89870 87508
rect 22094 87428 22100 87440
rect 12406 87400 22100 87428
rect 22094 87388 22100 87400
rect 22152 87388 22158 87440
rect 44450 87388 44456 87440
rect 44508 87428 44514 87440
rect 45094 87428 45100 87440
rect 44508 87400 45100 87428
rect 44508 87388 44514 87400
rect 45094 87388 45100 87400
rect 45152 87428 45158 87440
rect 45152 87400 90680 87428
rect 45152 87388 45158 87400
rect 2041 87363 2099 87369
rect 2041 87329 2053 87363
rect 2087 87329 2099 87363
rect 2041 87323 2099 87329
rect 2410 87363 2468 87369
rect 2410 87329 2422 87363
rect 2456 87329 2468 87363
rect 2410 87323 2468 87329
rect 2593 87363 2651 87369
rect 2593 87329 2605 87363
rect 2639 87329 2651 87363
rect 27890 87360 27896 87372
rect 27851 87332 27896 87360
rect 2593 87323 2651 87329
rect 2225 87295 2283 87301
rect 2225 87261 2237 87295
rect 2271 87261 2283 87295
rect 2225 87255 2283 87261
rect 1765 87227 1823 87233
rect 1765 87193 1777 87227
rect 1811 87224 1823 87227
rect 2240 87224 2268 87255
rect 2314 87252 2320 87304
rect 2372 87292 2378 87304
rect 2372 87264 2417 87292
rect 2372 87252 2378 87264
rect 2406 87224 2412 87236
rect 1811 87196 2176 87224
rect 2240 87196 2412 87224
rect 1811 87193 1823 87196
rect 1765 87187 1823 87193
rect 1946 87156 1952 87168
rect 1907 87128 1952 87156
rect 1946 87116 1952 87128
rect 2004 87116 2010 87168
rect 2148 87156 2176 87196
rect 2406 87184 2412 87196
rect 2464 87184 2470 87236
rect 2608 87224 2636 87323
rect 27890 87320 27896 87332
rect 27948 87320 27954 87372
rect 29270 87360 29276 87372
rect 28276 87332 29276 87360
rect 28276 87292 28304 87332
rect 29270 87320 29276 87332
rect 29328 87320 29334 87372
rect 59906 87320 59912 87372
rect 59964 87360 59970 87372
rect 73157 87363 73215 87369
rect 73157 87360 73169 87363
rect 59964 87332 73169 87360
rect 59964 87320 59970 87332
rect 73157 87329 73169 87332
rect 73203 87329 73215 87363
rect 73522 87360 73528 87372
rect 73483 87332 73528 87360
rect 73157 87323 73215 87329
rect 73522 87320 73528 87332
rect 73580 87320 73586 87372
rect 73890 87360 73896 87372
rect 73851 87332 73896 87360
rect 73890 87320 73896 87332
rect 73948 87320 73954 87372
rect 74077 87363 74135 87369
rect 74077 87329 74089 87363
rect 74123 87360 74135 87363
rect 74534 87360 74540 87372
rect 74123 87332 74540 87360
rect 74123 87329 74135 87332
rect 74077 87323 74135 87329
rect 74534 87320 74540 87332
rect 74592 87360 74598 87372
rect 75362 87360 75368 87372
rect 74592 87332 75368 87360
rect 74592 87320 74598 87332
rect 75362 87320 75368 87332
rect 75420 87320 75426 87372
rect 89898 87360 89904 87372
rect 89859 87332 89904 87360
rect 89898 87320 89904 87332
rect 89956 87320 89962 87372
rect 90266 87360 90272 87372
rect 90227 87332 90272 87360
rect 90266 87320 90272 87332
rect 90324 87320 90330 87372
rect 90652 87369 90680 87400
rect 90637 87363 90695 87369
rect 90637 87329 90649 87363
rect 90683 87329 90695 87363
rect 90637 87323 90695 87329
rect 28442 87292 28448 87304
rect 2746 87264 28304 87292
rect 28403 87264 28448 87292
rect 2746 87224 2774 87264
rect 28442 87252 28448 87264
rect 28500 87252 28506 87304
rect 73617 87295 73675 87301
rect 57946 87264 67634 87292
rect 2608 87196 2774 87224
rect 2608 87156 2636 87196
rect 10134 87184 10140 87236
rect 10192 87224 10198 87236
rect 57946 87224 57974 87264
rect 10192 87196 57974 87224
rect 67606 87224 67634 87264
rect 70366 87264 73292 87292
rect 70366 87224 70394 87264
rect 67606 87196 70394 87224
rect 73264 87224 73292 87264
rect 73617 87261 73629 87295
rect 73663 87292 73675 87295
rect 73706 87292 73712 87304
rect 73663 87264 73712 87292
rect 73663 87261 73675 87264
rect 73617 87255 73675 87261
rect 73706 87252 73712 87264
rect 73764 87252 73770 87304
rect 90082 87292 90088 87304
rect 90043 87264 90088 87292
rect 90082 87252 90088 87264
rect 90140 87252 90146 87304
rect 90545 87295 90603 87301
rect 90545 87261 90557 87295
rect 90591 87261 90603 87295
rect 90545 87255 90603 87261
rect 74261 87227 74319 87233
rect 74261 87224 74273 87227
rect 73264 87196 74273 87224
rect 10192 87184 10198 87196
rect 74261 87193 74273 87196
rect 74307 87193 74319 87227
rect 89806 87224 89812 87236
rect 89719 87196 89812 87224
rect 74261 87187 74319 87193
rect 89806 87184 89812 87196
rect 89864 87224 89870 87236
rect 90560 87224 90588 87255
rect 91002 87224 91008 87236
rect 89864 87196 90588 87224
rect 90963 87196 91008 87224
rect 89864 87184 89870 87196
rect 91002 87184 91008 87196
rect 91060 87184 91066 87236
rect 2148 87128 2636 87156
rect 35250 87116 35256 87168
rect 35308 87156 35314 87168
rect 59906 87156 59912 87168
rect 35308 87128 59912 87156
rect 35308 87116 35314 87128
rect 59906 87116 59912 87128
rect 59964 87116 59970 87168
rect 1104 87066 98808 87088
rect 1104 87014 4246 87066
rect 4298 87014 4310 87066
rect 4362 87014 4374 87066
rect 4426 87014 4438 87066
rect 4490 87014 34966 87066
rect 35018 87014 35030 87066
rect 35082 87014 35094 87066
rect 35146 87014 35158 87066
rect 35210 87014 65686 87066
rect 65738 87014 65750 87066
rect 65802 87014 65814 87066
rect 65866 87014 65878 87066
rect 65930 87014 96406 87066
rect 96458 87014 96470 87066
rect 96522 87014 96534 87066
rect 96586 87014 96598 87066
rect 96650 87014 98808 87066
rect 1104 86992 98808 87014
rect 29362 86912 29368 86964
rect 29420 86952 29426 86964
rect 30190 86952 30196 86964
rect 29420 86924 30196 86952
rect 29420 86912 29426 86924
rect 30190 86912 30196 86924
rect 30248 86912 30254 86964
rect 12526 86884 12532 86896
rect 12452 86856 12532 86884
rect 12345 86819 12403 86825
rect 12345 86785 12357 86819
rect 12391 86816 12403 86819
rect 12452 86816 12480 86856
rect 12526 86844 12532 86856
rect 12584 86844 12590 86896
rect 12391 86788 12480 86816
rect 12897 86819 12955 86825
rect 12391 86785 12403 86788
rect 12345 86779 12403 86785
rect 12897 86785 12909 86819
rect 12943 86816 12955 86819
rect 34514 86816 34520 86828
rect 12943 86788 34520 86816
rect 12943 86785 12955 86788
rect 12897 86779 12955 86785
rect 34514 86776 34520 86788
rect 34572 86776 34578 86828
rect 12066 86748 12072 86760
rect 12027 86720 12072 86748
rect 12066 86708 12072 86720
rect 12124 86708 12130 86760
rect 12437 86751 12495 86757
rect 12437 86717 12449 86751
rect 12483 86717 12495 86751
rect 12802 86748 12808 86760
rect 12763 86720 12808 86748
rect 12437 86711 12495 86717
rect 12452 86680 12480 86711
rect 12802 86708 12808 86720
rect 12860 86708 12866 86760
rect 29362 86708 29368 86760
rect 29420 86748 29426 86760
rect 29457 86751 29515 86757
rect 29457 86748 29469 86751
rect 29420 86720 29469 86748
rect 29420 86708 29426 86720
rect 29457 86717 29469 86720
rect 29503 86717 29515 86751
rect 29730 86748 29736 86760
rect 29691 86720 29736 86748
rect 29457 86711 29515 86717
rect 29730 86708 29736 86720
rect 29788 86708 29794 86760
rect 55861 86751 55919 86757
rect 55861 86717 55873 86751
rect 55907 86748 55919 86751
rect 56137 86751 56195 86757
rect 56137 86748 56149 86751
rect 55907 86720 56149 86748
rect 55907 86717 55919 86720
rect 55861 86711 55919 86717
rect 56137 86717 56149 86720
rect 56183 86748 56195 86751
rect 64138 86748 64144 86760
rect 56183 86720 64144 86748
rect 56183 86717 56195 86720
rect 56137 86711 56195 86717
rect 64138 86708 64144 86720
rect 64196 86708 64202 86760
rect 24210 86680 24216 86692
rect 12452 86652 24216 86680
rect 24210 86640 24216 86652
rect 24268 86640 24274 86692
rect 31113 86683 31171 86689
rect 30760 86652 30972 86680
rect 13265 86615 13323 86621
rect 13265 86581 13277 86615
rect 13311 86612 13323 86615
rect 30760 86612 30788 86652
rect 13311 86584 30788 86612
rect 30944 86612 30972 86652
rect 31113 86649 31125 86683
rect 31159 86680 31171 86683
rect 46842 86680 46848 86692
rect 31159 86652 46848 86680
rect 31159 86649 31171 86652
rect 31113 86643 31171 86649
rect 46842 86640 46848 86652
rect 46900 86640 46906 86692
rect 55186 86652 60734 86680
rect 55186 86612 55214 86652
rect 30944 86584 55214 86612
rect 60706 86612 60734 86652
rect 90542 86612 90548 86624
rect 60706 86584 90548 86612
rect 13311 86581 13323 86584
rect 13265 86575 13323 86581
rect 90542 86572 90548 86584
rect 90600 86572 90606 86624
rect 1104 86522 98808 86544
rect 1104 86470 19606 86522
rect 19658 86470 19670 86522
rect 19722 86470 19734 86522
rect 19786 86470 19798 86522
rect 19850 86470 50326 86522
rect 50378 86470 50390 86522
rect 50442 86470 50454 86522
rect 50506 86470 50518 86522
rect 50570 86470 81046 86522
rect 81098 86470 81110 86522
rect 81162 86470 81174 86522
rect 81226 86470 81238 86522
rect 81290 86470 98808 86522
rect 1104 86448 98808 86470
rect 12066 86300 12072 86352
rect 12124 86340 12130 86352
rect 46290 86340 46296 86352
rect 12124 86312 46296 86340
rect 12124 86300 12130 86312
rect 46290 86300 46296 86312
rect 46348 86300 46354 86352
rect 54662 86300 54668 86352
rect 54720 86340 54726 86352
rect 74626 86340 74632 86352
rect 54720 86312 74632 86340
rect 54720 86300 54726 86312
rect 74626 86300 74632 86312
rect 74684 86300 74690 86352
rect 43530 86272 43536 86284
rect 43491 86244 43536 86272
rect 43530 86232 43536 86244
rect 43588 86232 43594 86284
rect 49050 86232 49056 86284
rect 49108 86272 49114 86284
rect 73798 86272 73804 86284
rect 49108 86244 73804 86272
rect 49108 86232 49114 86244
rect 73798 86232 73804 86244
rect 73856 86232 73862 86284
rect 44177 86207 44235 86213
rect 44177 86173 44189 86207
rect 44223 86204 44235 86207
rect 44910 86204 44916 86216
rect 44223 86176 44916 86204
rect 44223 86173 44235 86176
rect 44177 86167 44235 86173
rect 44910 86164 44916 86176
rect 44968 86164 44974 86216
rect 82817 86207 82875 86213
rect 82817 86173 82829 86207
rect 82863 86204 82875 86207
rect 83090 86204 83096 86216
rect 82863 86176 83096 86204
rect 82863 86173 82875 86176
rect 82817 86167 82875 86173
rect 83090 86164 83096 86176
rect 83148 86204 83154 86216
rect 84289 86207 84347 86213
rect 84289 86204 84301 86207
rect 83148 86176 84301 86204
rect 83148 86164 83154 86176
rect 84289 86173 84301 86176
rect 84335 86173 84347 86207
rect 84562 86204 84568 86216
rect 84523 86176 84568 86204
rect 84289 86167 84347 86173
rect 84562 86164 84568 86176
rect 84620 86164 84626 86216
rect 82814 86028 82820 86080
rect 82872 86068 82878 86080
rect 83001 86071 83059 86077
rect 83001 86068 83013 86071
rect 82872 86040 83013 86068
rect 82872 86028 82878 86040
rect 83001 86037 83013 86040
rect 83047 86037 83059 86071
rect 83001 86031 83059 86037
rect 89809 86071 89867 86077
rect 89809 86037 89821 86071
rect 89855 86068 89867 86071
rect 89901 86071 89959 86077
rect 89901 86068 89913 86071
rect 89855 86040 89913 86068
rect 89855 86037 89867 86040
rect 89809 86031 89867 86037
rect 89901 86037 89913 86040
rect 89947 86068 89959 86071
rect 90266 86068 90272 86080
rect 89947 86040 90272 86068
rect 89947 86037 89959 86040
rect 89901 86031 89959 86037
rect 90266 86028 90272 86040
rect 90324 86028 90330 86080
rect 97445 86071 97503 86077
rect 97445 86037 97457 86071
rect 97491 86068 97503 86071
rect 97626 86068 97632 86080
rect 97491 86040 97632 86068
rect 97491 86037 97503 86040
rect 97445 86031 97503 86037
rect 97626 86028 97632 86040
rect 97684 86068 97690 86080
rect 97721 86071 97779 86077
rect 97721 86068 97733 86071
rect 97684 86040 97733 86068
rect 97684 86028 97690 86040
rect 97721 86037 97733 86040
rect 97767 86037 97779 86071
rect 97721 86031 97779 86037
rect 1104 85978 98808 86000
rect 1104 85926 4246 85978
rect 4298 85926 4310 85978
rect 4362 85926 4374 85978
rect 4426 85926 4438 85978
rect 4490 85926 34966 85978
rect 35018 85926 35030 85978
rect 35082 85926 35094 85978
rect 35146 85926 35158 85978
rect 35210 85926 65686 85978
rect 65738 85926 65750 85978
rect 65802 85926 65814 85978
rect 65866 85926 65878 85978
rect 65930 85926 96406 85978
rect 96458 85926 96470 85978
rect 96522 85926 96534 85978
rect 96586 85926 96598 85978
rect 96650 85926 98808 85978
rect 1104 85904 98808 85926
rect 80977 85663 81035 85669
rect 80977 85629 80989 85663
rect 81023 85660 81035 85663
rect 81253 85663 81311 85669
rect 81253 85660 81265 85663
rect 81023 85632 81265 85660
rect 81023 85629 81035 85632
rect 80977 85623 81035 85629
rect 81253 85629 81265 85632
rect 81299 85660 81311 85663
rect 82078 85660 82084 85672
rect 81299 85632 82084 85660
rect 81299 85629 81311 85632
rect 81253 85623 81311 85629
rect 82078 85620 82084 85632
rect 82136 85620 82142 85672
rect 87233 85663 87291 85669
rect 87233 85629 87245 85663
rect 87279 85629 87291 85663
rect 87233 85623 87291 85629
rect 23658 85592 23664 85604
rect 23619 85564 23664 85592
rect 23658 85552 23664 85564
rect 23716 85552 23722 85604
rect 24394 85592 24400 85604
rect 24355 85564 24400 85592
rect 24394 85552 24400 85564
rect 24452 85552 24458 85604
rect 45002 85552 45008 85604
rect 45060 85592 45066 85604
rect 87049 85595 87107 85601
rect 87049 85592 87061 85595
rect 45060 85564 87061 85592
rect 45060 85552 45066 85564
rect 87049 85561 87061 85564
rect 87095 85592 87107 85595
rect 87248 85592 87276 85623
rect 87095 85564 87276 85592
rect 87095 85561 87107 85564
rect 87049 85555 87107 85561
rect 30374 85484 30380 85536
rect 30432 85524 30438 85536
rect 31294 85524 31300 85536
rect 30432 85496 31300 85524
rect 30432 85484 30438 85496
rect 31294 85484 31300 85496
rect 31352 85484 31358 85536
rect 1104 85434 98808 85456
rect 1104 85382 19606 85434
rect 19658 85382 19670 85434
rect 19722 85382 19734 85434
rect 19786 85382 19798 85434
rect 19850 85382 50326 85434
rect 50378 85382 50390 85434
rect 50442 85382 50454 85434
rect 50506 85382 50518 85434
rect 50570 85382 81046 85434
rect 81098 85382 81110 85434
rect 81162 85382 81174 85434
rect 81226 85382 81238 85434
rect 81290 85382 98808 85434
rect 1104 85360 98808 85382
rect 10502 85280 10508 85332
rect 10560 85320 10566 85332
rect 10560 85292 14044 85320
rect 10560 85280 10566 85292
rect 10594 85252 10600 85264
rect 4724 85224 10600 85252
rect 4724 85193 4752 85224
rect 10594 85212 10600 85224
rect 10652 85212 10658 85264
rect 4709 85187 4767 85193
rect 4709 85153 4721 85187
rect 4755 85153 4767 85187
rect 5074 85184 5080 85196
rect 5035 85156 5080 85184
rect 4709 85147 4767 85153
rect 5074 85144 5080 85156
rect 5132 85144 5138 85196
rect 10042 85144 10048 85196
rect 10100 85184 10106 85196
rect 10137 85187 10195 85193
rect 10137 85184 10149 85187
rect 10100 85156 10149 85184
rect 10100 85144 10106 85156
rect 10137 85153 10149 85156
rect 10183 85153 10195 85187
rect 10137 85147 10195 85153
rect 10502 85144 10508 85196
rect 10560 85184 10566 85196
rect 14016 85184 14044 85292
rect 14642 85280 14648 85332
rect 14700 85320 14706 85332
rect 31846 85320 31852 85332
rect 14700 85292 31852 85320
rect 14700 85280 14706 85292
rect 31846 85280 31852 85292
rect 31904 85280 31910 85332
rect 45462 85280 45468 85332
rect 45520 85320 45526 85332
rect 45520 85292 46704 85320
rect 45520 85280 45526 85292
rect 14185 85255 14243 85261
rect 14185 85221 14197 85255
rect 14231 85252 14243 85255
rect 23658 85252 23664 85264
rect 14231 85224 23664 85252
rect 14231 85221 14243 85224
rect 14185 85215 14243 85221
rect 23658 85212 23664 85224
rect 23716 85212 23722 85264
rect 30006 85212 30012 85264
rect 30064 85252 30070 85264
rect 30064 85224 46520 85252
rect 30064 85212 30070 85224
rect 31849 85187 31907 85193
rect 10560 85156 10605 85184
rect 14016 85156 19334 85184
rect 10560 85144 10566 85156
rect 5169 85119 5227 85125
rect 5169 85085 5181 85119
rect 5215 85116 5227 85119
rect 6454 85116 6460 85128
rect 5215 85088 6460 85116
rect 5215 85085 5227 85088
rect 5169 85079 5227 85085
rect 6454 85076 6460 85088
rect 6512 85076 6518 85128
rect 9582 85116 9588 85128
rect 9543 85088 9588 85116
rect 9582 85076 9588 85088
rect 9640 85076 9646 85128
rect 10226 85116 10232 85128
rect 9784 85088 9996 85116
rect 10187 85088 10232 85116
rect 4525 85051 4583 85057
rect 4525 85017 4537 85051
rect 4571 85048 4583 85051
rect 9784 85048 9812 85088
rect 4571 85020 9812 85048
rect 9968 85048 9996 85088
rect 10226 85076 10232 85088
rect 10284 85076 10290 85128
rect 10318 85076 10324 85128
rect 10376 85116 10382 85128
rect 10413 85119 10471 85125
rect 10413 85116 10425 85119
rect 10376 85088 10425 85116
rect 10376 85076 10382 85088
rect 10413 85085 10425 85088
rect 10459 85085 10471 85119
rect 19306 85116 19334 85156
rect 31849 85153 31861 85187
rect 31895 85184 31907 85187
rect 32582 85184 32588 85196
rect 31895 85156 32588 85184
rect 31895 85153 31907 85156
rect 31849 85147 31907 85153
rect 32582 85144 32588 85156
rect 32640 85144 32646 85196
rect 46290 85184 46296 85196
rect 46251 85156 46296 85184
rect 46290 85144 46296 85156
rect 46348 85144 46354 85196
rect 46492 85193 46520 85224
rect 46676 85193 46704 85292
rect 50154 85280 50160 85332
rect 50212 85320 50218 85332
rect 74902 85320 74908 85332
rect 50212 85292 74908 85320
rect 50212 85280 50218 85292
rect 74902 85280 74908 85292
rect 74960 85280 74966 85332
rect 53926 85212 53932 85264
rect 53984 85252 53990 85264
rect 95694 85252 95700 85264
rect 53984 85224 95700 85252
rect 53984 85212 53990 85224
rect 95694 85212 95700 85224
rect 95752 85212 95758 85264
rect 46476 85187 46534 85193
rect 46476 85153 46488 85187
rect 46522 85153 46534 85187
rect 46476 85147 46534 85153
rect 46661 85187 46719 85193
rect 46661 85153 46673 85187
rect 46707 85153 46719 85187
rect 46661 85147 46719 85153
rect 46750 85144 46756 85196
rect 46808 85184 46814 85196
rect 46845 85187 46903 85193
rect 46845 85184 46857 85187
rect 46808 85156 46857 85184
rect 46808 85144 46814 85156
rect 46845 85153 46857 85156
rect 46891 85184 46903 85187
rect 56962 85184 56968 85196
rect 46891 85156 56968 85184
rect 46891 85153 46903 85156
rect 46845 85147 46903 85153
rect 56962 85144 56968 85156
rect 57020 85144 57026 85196
rect 72510 85184 72516 85196
rect 72471 85156 72516 85184
rect 72510 85144 72516 85156
rect 72568 85144 72574 85196
rect 30374 85116 30380 85128
rect 19306 85088 30380 85116
rect 10413 85079 10471 85085
rect 30374 85076 30380 85088
rect 30432 85076 30438 85128
rect 32493 85119 32551 85125
rect 32493 85085 32505 85119
rect 32539 85116 32551 85119
rect 45186 85116 45192 85128
rect 32539 85088 45192 85116
rect 32539 85085 32551 85088
rect 32493 85079 32551 85085
rect 45186 85076 45192 85088
rect 45244 85076 45250 85128
rect 46566 85116 46572 85128
rect 46527 85088 46572 85116
rect 46566 85076 46572 85088
rect 46624 85076 46630 85128
rect 46934 85076 46940 85128
rect 46992 85116 46998 85128
rect 47029 85119 47087 85125
rect 47029 85116 47041 85119
rect 46992 85088 47041 85116
rect 46992 85076 46998 85088
rect 47029 85085 47041 85088
rect 47075 85085 47087 85119
rect 47029 85079 47087 85085
rect 73065 85119 73123 85125
rect 73065 85085 73077 85119
rect 73111 85116 73123 85119
rect 79502 85116 79508 85128
rect 73111 85088 79508 85116
rect 73111 85085 73123 85088
rect 73065 85079 73123 85085
rect 79502 85076 79508 85088
rect 79560 85076 79566 85128
rect 82630 85048 82636 85060
rect 9968 85020 46612 85048
rect 4571 85017 4583 85020
rect 4525 85011 4583 85017
rect 10594 84940 10600 84992
rect 10652 84980 10658 84992
rect 14185 84983 14243 84989
rect 14185 84980 14197 84983
rect 10652 84952 14197 84980
rect 10652 84940 10658 84952
rect 14185 84949 14197 84952
rect 14231 84949 14243 84983
rect 14185 84943 14243 84949
rect 34146 84940 34152 84992
rect 34204 84980 34210 84992
rect 46474 84980 46480 84992
rect 34204 84952 46480 84980
rect 34204 84940 34210 84952
rect 46474 84940 46480 84952
rect 46532 84940 46538 84992
rect 46584 84980 46612 85020
rect 46860 85020 82636 85048
rect 46860 84980 46888 85020
rect 82630 85008 82636 85020
rect 82688 85008 82694 85060
rect 46584 84952 46888 84980
rect 61102 84940 61108 84992
rect 61160 84980 61166 84992
rect 61749 84983 61807 84989
rect 61749 84980 61761 84983
rect 61160 84952 61761 84980
rect 61160 84940 61166 84952
rect 61749 84949 61761 84952
rect 61795 84980 61807 84983
rect 61933 84983 61991 84989
rect 61933 84980 61945 84983
rect 61795 84952 61945 84980
rect 61795 84949 61807 84952
rect 61749 84943 61807 84949
rect 61933 84949 61945 84952
rect 61979 84949 61991 84983
rect 61933 84943 61991 84949
rect 1104 84890 98808 84912
rect 1104 84838 4246 84890
rect 4298 84838 4310 84890
rect 4362 84838 4374 84890
rect 4426 84838 4438 84890
rect 4490 84838 34966 84890
rect 35018 84838 35030 84890
rect 35082 84838 35094 84890
rect 35146 84838 35158 84890
rect 35210 84838 65686 84890
rect 65738 84838 65750 84890
rect 65802 84838 65814 84890
rect 65866 84838 65878 84890
rect 65930 84838 96406 84890
rect 96458 84838 96470 84890
rect 96522 84838 96534 84890
rect 96586 84838 96598 84890
rect 96650 84838 98808 84890
rect 1104 84816 98808 84838
rect 38473 84779 38531 84785
rect 38473 84745 38485 84779
rect 38519 84776 38531 84779
rect 42058 84776 42064 84788
rect 38519 84748 42064 84776
rect 38519 84745 38531 84748
rect 38473 84739 38531 84745
rect 42058 84736 42064 84748
rect 42116 84736 42122 84788
rect 39850 84668 39856 84720
rect 39908 84708 39914 84720
rect 50154 84708 50160 84720
rect 39908 84680 50160 84708
rect 39908 84668 39914 84680
rect 50154 84668 50160 84680
rect 50212 84668 50218 84720
rect 62025 84575 62083 84581
rect 62025 84541 62037 84575
rect 62071 84572 62083 84575
rect 62298 84572 62304 84584
rect 62071 84544 62304 84572
rect 62071 84541 62083 84544
rect 62025 84535 62083 84541
rect 62298 84532 62304 84544
rect 62356 84532 62362 84584
rect 85758 84572 85764 84584
rect 85719 84544 85764 84572
rect 85758 84532 85764 84544
rect 85816 84532 85822 84584
rect 85942 84436 85948 84448
rect 85903 84408 85948 84436
rect 85942 84396 85948 84408
rect 86000 84396 86006 84448
rect 1104 84346 98808 84368
rect 1104 84294 19606 84346
rect 19658 84294 19670 84346
rect 19722 84294 19734 84346
rect 19786 84294 19798 84346
rect 19850 84294 50326 84346
rect 50378 84294 50390 84346
rect 50442 84294 50454 84346
rect 50506 84294 50518 84346
rect 50570 84294 81046 84346
rect 81098 84294 81110 84346
rect 81162 84294 81174 84346
rect 81226 84294 81238 84346
rect 81290 84294 98808 84346
rect 1104 84272 98808 84294
rect 87601 84235 87659 84241
rect 87601 84201 87613 84235
rect 87647 84232 87659 84235
rect 96341 84235 96399 84241
rect 96341 84232 96353 84235
rect 87647 84204 96353 84232
rect 87647 84201 87659 84204
rect 87601 84195 87659 84201
rect 96341 84201 96353 84204
rect 96387 84201 96399 84235
rect 96341 84195 96399 84201
rect 65978 84124 65984 84176
rect 66036 84164 66042 84176
rect 66036 84136 85896 84164
rect 66036 84124 66042 84136
rect 47578 84056 47584 84108
rect 47636 84096 47642 84108
rect 85868 84105 85896 84136
rect 85960 84136 97212 84164
rect 85853 84099 85911 84105
rect 47636 84068 85804 84096
rect 47636 84056 47642 84068
rect 60366 83988 60372 84040
rect 60424 84028 60430 84040
rect 79318 84028 79324 84040
rect 60424 84000 79324 84028
rect 60424 83988 60430 84000
rect 79318 83988 79324 84000
rect 79376 83988 79382 84040
rect 85298 84028 85304 84040
rect 85259 84000 85304 84028
rect 85298 83988 85304 84000
rect 85356 83988 85362 84040
rect 85666 84028 85672 84040
rect 85627 84000 85672 84028
rect 85666 83988 85672 84000
rect 85724 83988 85730 84040
rect 85776 84028 85804 84068
rect 85853 84065 85865 84099
rect 85899 84065 85911 84099
rect 85853 84059 85911 84065
rect 85960 84028 85988 84136
rect 86218 84096 86224 84108
rect 86179 84068 86224 84096
rect 86218 84056 86224 84068
rect 86276 84056 86282 84108
rect 97184 84105 97212 84136
rect 97169 84099 97227 84105
rect 89686 84068 97120 84096
rect 86126 84028 86132 84040
rect 85776 84000 85988 84028
rect 86087 84000 86132 84028
rect 86126 83988 86132 84000
rect 86184 83988 86190 84040
rect 88518 83988 88524 84040
rect 88576 84028 88582 84040
rect 89686 84028 89714 84068
rect 96985 84031 97043 84037
rect 96985 84028 96997 84031
rect 88576 84000 89714 84028
rect 91296 84000 96997 84028
rect 88576 83988 88582 84000
rect 62022 83920 62028 83972
rect 62080 83960 62086 83972
rect 87601 83963 87659 83969
rect 87601 83960 87613 83963
rect 62080 83932 87613 83960
rect 62080 83920 62086 83932
rect 87601 83929 87613 83932
rect 87647 83929 87659 83963
rect 87601 83923 87659 83929
rect 34517 83895 34575 83901
rect 34517 83861 34529 83895
rect 34563 83892 34575 83895
rect 34793 83895 34851 83901
rect 34793 83892 34805 83895
rect 34563 83864 34805 83892
rect 34563 83861 34575 83864
rect 34517 83855 34575 83861
rect 34793 83861 34805 83864
rect 34839 83892 34851 83895
rect 65518 83892 65524 83904
rect 34839 83864 65524 83892
rect 34839 83861 34851 83864
rect 34793 83855 34851 83861
rect 65518 83852 65524 83864
rect 65576 83852 65582 83904
rect 66898 83852 66904 83904
rect 66956 83892 66962 83904
rect 67542 83892 67548 83904
rect 66956 83864 67548 83892
rect 66956 83852 66962 83864
rect 67542 83852 67548 83864
rect 67600 83892 67606 83904
rect 91296 83892 91324 84000
rect 96985 83997 96997 84000
rect 97031 83997 97043 84031
rect 97092 84028 97120 84068
rect 97169 84065 97181 84099
rect 97215 84065 97227 84099
rect 97537 84099 97595 84105
rect 97537 84096 97549 84099
rect 97169 84059 97227 84065
rect 97276 84068 97549 84096
rect 97276 84028 97304 84068
rect 97537 84065 97549 84068
rect 97583 84065 97595 84099
rect 97537 84059 97595 84065
rect 97092 84000 97304 84028
rect 97445 84031 97503 84037
rect 96985 83991 97043 83997
rect 97445 83997 97457 84031
rect 97491 83997 97503 84031
rect 97445 83991 97503 83997
rect 96341 83963 96399 83969
rect 96341 83929 96353 83963
rect 96387 83960 96399 83963
rect 97460 83960 97488 83991
rect 96387 83932 97488 83960
rect 96387 83929 96399 83932
rect 96341 83923 96399 83929
rect 67600 83864 91324 83892
rect 96801 83895 96859 83901
rect 67600 83852 67606 83864
rect 96801 83861 96813 83895
rect 96847 83892 96859 83895
rect 96890 83892 96896 83904
rect 96847 83864 96896 83892
rect 96847 83861 96859 83864
rect 96801 83855 96859 83861
rect 96890 83852 96896 83864
rect 96948 83852 96954 83904
rect 1104 83802 98808 83824
rect 1104 83750 4246 83802
rect 4298 83750 4310 83802
rect 4362 83750 4374 83802
rect 4426 83750 4438 83802
rect 4490 83750 34966 83802
rect 35018 83750 35030 83802
rect 35082 83750 35094 83802
rect 35146 83750 35158 83802
rect 35210 83750 65686 83802
rect 65738 83750 65750 83802
rect 65802 83750 65814 83802
rect 65866 83750 65878 83802
rect 65930 83750 96406 83802
rect 96458 83750 96470 83802
rect 96522 83750 96534 83802
rect 96586 83750 96598 83802
rect 96650 83750 98808 83802
rect 1104 83728 98808 83750
rect 71038 83648 71044 83700
rect 71096 83688 71102 83700
rect 71096 83660 79180 83688
rect 71096 83648 71102 83660
rect 12802 83580 12808 83632
rect 12860 83620 12866 83632
rect 21082 83620 21088 83632
rect 12860 83592 21088 83620
rect 12860 83580 12866 83592
rect 21082 83580 21088 83592
rect 21140 83580 21146 83632
rect 20346 83512 20352 83564
rect 20404 83552 20410 83564
rect 31202 83552 31208 83564
rect 20404 83524 31208 83552
rect 20404 83512 20410 83524
rect 31202 83512 31208 83524
rect 31260 83512 31266 83564
rect 79152 83552 79180 83660
rect 79318 83648 79324 83700
rect 79376 83688 79382 83700
rect 88518 83688 88524 83700
rect 79376 83660 88524 83688
rect 79376 83648 79382 83660
rect 88518 83648 88524 83660
rect 88576 83648 88582 83700
rect 86218 83552 86224 83564
rect 79152 83524 86224 83552
rect 86218 83512 86224 83524
rect 86276 83512 86282 83564
rect 19337 83487 19395 83493
rect 19337 83453 19349 83487
rect 19383 83484 19395 83487
rect 19613 83487 19671 83493
rect 19613 83484 19625 83487
rect 19383 83456 19625 83484
rect 19383 83453 19395 83456
rect 19337 83447 19395 83453
rect 19613 83453 19625 83456
rect 19659 83484 19671 83487
rect 64322 83484 64328 83496
rect 19659 83456 64328 83484
rect 19659 83453 19671 83456
rect 19613 83447 19671 83453
rect 64322 83444 64328 83456
rect 64380 83444 64386 83496
rect 71130 83444 71136 83496
rect 71188 83484 71194 83496
rect 86126 83484 86132 83496
rect 71188 83456 86132 83484
rect 71188 83444 71194 83456
rect 86126 83444 86132 83456
rect 86184 83444 86190 83496
rect 97166 83376 97172 83428
rect 97224 83416 97230 83428
rect 97905 83419 97963 83425
rect 97905 83416 97917 83419
rect 97224 83388 97917 83416
rect 97224 83376 97230 83388
rect 97905 83385 97917 83388
rect 97951 83385 97963 83419
rect 97905 83379 97963 83385
rect 97994 83348 98000 83360
rect 97955 83320 98000 83348
rect 97994 83308 98000 83320
rect 98052 83308 98058 83360
rect 1104 83258 98808 83280
rect 1104 83206 19606 83258
rect 19658 83206 19670 83258
rect 19722 83206 19734 83258
rect 19786 83206 19798 83258
rect 19850 83206 50326 83258
rect 50378 83206 50390 83258
rect 50442 83206 50454 83258
rect 50506 83206 50518 83258
rect 50570 83206 81046 83258
rect 81098 83206 81110 83258
rect 81162 83206 81174 83258
rect 81226 83206 81238 83258
rect 81290 83206 98808 83258
rect 1104 83184 98808 83206
rect 26602 82968 26608 83020
rect 26660 83008 26666 83020
rect 76193 83011 76251 83017
rect 76193 83008 76205 83011
rect 26660 82980 76205 83008
rect 26660 82968 26666 82980
rect 76193 82977 76205 82980
rect 76239 82977 76251 83011
rect 76558 83008 76564 83020
rect 76519 82980 76564 83008
rect 76193 82971 76251 82977
rect 76558 82968 76564 82980
rect 76616 82968 76622 83020
rect 75638 82940 75644 82952
rect 75599 82912 75644 82940
rect 75638 82900 75644 82912
rect 75696 82900 75702 82952
rect 76006 82940 76012 82952
rect 75967 82912 76012 82940
rect 76006 82900 76012 82912
rect 76064 82900 76070 82952
rect 76466 82940 76472 82952
rect 76427 82912 76472 82940
rect 76466 82900 76472 82912
rect 76524 82900 76530 82952
rect 1104 82714 98808 82736
rect 1104 82662 4246 82714
rect 4298 82662 4310 82714
rect 4362 82662 4374 82714
rect 4426 82662 4438 82714
rect 4490 82662 34966 82714
rect 35018 82662 35030 82714
rect 35082 82662 35094 82714
rect 35146 82662 35158 82714
rect 35210 82662 65686 82714
rect 65738 82662 65750 82714
rect 65802 82662 65814 82714
rect 65866 82662 65878 82714
rect 65930 82662 96406 82714
rect 96458 82662 96470 82714
rect 96522 82662 96534 82714
rect 96586 82662 96598 82714
rect 96650 82662 98808 82714
rect 1104 82640 98808 82662
rect 53834 82424 53840 82476
rect 53892 82464 53898 82476
rect 68830 82464 68836 82476
rect 53892 82436 68836 82464
rect 53892 82424 53898 82436
rect 68830 82424 68836 82436
rect 68888 82424 68894 82476
rect 61194 82396 61200 82408
rect 60706 82368 61200 82396
rect 6914 82288 6920 82340
rect 6972 82328 6978 82340
rect 39482 82328 39488 82340
rect 6972 82300 39488 82328
rect 6972 82288 6978 82300
rect 39482 82288 39488 82300
rect 39540 82288 39546 82340
rect 41874 82288 41880 82340
rect 41932 82328 41938 82340
rect 60706 82328 60734 82368
rect 61194 82356 61200 82368
rect 61252 82356 61258 82408
rect 65337 82399 65395 82405
rect 65337 82365 65349 82399
rect 65383 82396 65395 82399
rect 65613 82399 65671 82405
rect 65613 82396 65625 82399
rect 65383 82368 65625 82396
rect 65383 82365 65395 82368
rect 65337 82359 65395 82365
rect 65613 82365 65625 82368
rect 65659 82396 65671 82399
rect 65978 82396 65984 82408
rect 65659 82368 65984 82396
rect 65659 82365 65671 82368
rect 65613 82359 65671 82365
rect 65978 82356 65984 82368
rect 66036 82356 66042 82408
rect 41932 82300 60734 82328
rect 61028 82300 70394 82328
rect 41932 82288 41938 82300
rect 14642 82220 14648 82272
rect 14700 82260 14706 82272
rect 61028 82260 61056 82300
rect 14700 82232 61056 82260
rect 70366 82260 70394 82300
rect 71038 82260 71044 82272
rect 70366 82232 71044 82260
rect 14700 82220 14706 82232
rect 71038 82220 71044 82232
rect 71096 82220 71102 82272
rect 1104 82170 98808 82192
rect 1104 82118 19606 82170
rect 19658 82118 19670 82170
rect 19722 82118 19734 82170
rect 19786 82118 19798 82170
rect 19850 82118 50326 82170
rect 50378 82118 50390 82170
rect 50442 82118 50454 82170
rect 50506 82118 50518 82170
rect 50570 82118 81046 82170
rect 81098 82118 81110 82170
rect 81162 82118 81174 82170
rect 81226 82118 81238 82170
rect 81290 82118 98808 82170
rect 1104 82096 98808 82118
rect 91738 82016 91744 82068
rect 91796 82056 91802 82068
rect 93673 82059 93731 82065
rect 93673 82056 93685 82059
rect 91796 82028 93685 82056
rect 91796 82016 91802 82028
rect 93673 82025 93685 82028
rect 93719 82025 93731 82059
rect 93673 82019 93731 82025
rect 73798 81948 73804 82000
rect 73856 81988 73862 82000
rect 73856 81960 78260 81988
rect 73856 81948 73862 81960
rect 74074 81920 74080 81932
rect 74035 81892 74080 81920
rect 74074 81880 74080 81892
rect 74132 81920 74138 81932
rect 74132 81892 78168 81920
rect 74132 81880 74138 81892
rect 54294 81812 54300 81864
rect 54352 81852 54358 81864
rect 54478 81852 54484 81864
rect 54352 81824 54484 81852
rect 54352 81812 54358 81824
rect 54478 81812 54484 81824
rect 54536 81852 54542 81864
rect 74445 81855 74503 81861
rect 74445 81852 74457 81855
rect 54536 81824 74457 81852
rect 54536 81812 54542 81824
rect 74445 81821 74457 81824
rect 74491 81821 74503 81855
rect 74445 81815 74503 81821
rect 78140 81784 78168 81892
rect 78232 81852 78260 81960
rect 82998 81920 83004 81932
rect 82959 81892 83004 81920
rect 82998 81880 83004 81892
rect 83056 81880 83062 81932
rect 93688 81920 93716 82019
rect 94133 81923 94191 81929
rect 94133 81920 94145 81923
rect 93688 81892 94145 81920
rect 94133 81889 94145 81892
rect 94179 81889 94191 81923
rect 94133 81883 94191 81889
rect 83277 81855 83335 81861
rect 83277 81852 83289 81855
rect 78232 81824 83289 81852
rect 83277 81821 83289 81824
rect 83323 81821 83335 81855
rect 83277 81815 83335 81821
rect 92566 81812 92572 81864
rect 92624 81852 92630 81864
rect 93857 81855 93915 81861
rect 93857 81852 93869 81855
rect 92624 81824 93869 81852
rect 92624 81812 92630 81824
rect 93857 81821 93869 81824
rect 93903 81821 93915 81855
rect 93857 81815 93915 81821
rect 89898 81784 89904 81796
rect 78140 81756 89904 81784
rect 89898 81744 89904 81756
rect 89956 81744 89962 81796
rect 41233 81719 41291 81725
rect 41233 81685 41245 81719
rect 41279 81716 41291 81719
rect 89714 81716 89720 81728
rect 41279 81688 89720 81716
rect 41279 81685 41291 81688
rect 41233 81679 41291 81685
rect 89714 81676 89720 81688
rect 89772 81676 89778 81728
rect 95234 81716 95240 81728
rect 95195 81688 95240 81716
rect 95234 81676 95240 81688
rect 95292 81676 95298 81728
rect 1104 81626 98808 81648
rect 1104 81574 4246 81626
rect 4298 81574 4310 81626
rect 4362 81574 4374 81626
rect 4426 81574 4438 81626
rect 4490 81574 34966 81626
rect 35018 81574 35030 81626
rect 35082 81574 35094 81626
rect 35146 81574 35158 81626
rect 35210 81574 65686 81626
rect 65738 81574 65750 81626
rect 65802 81574 65814 81626
rect 65866 81574 65878 81626
rect 65930 81574 96406 81626
rect 96458 81574 96470 81626
rect 96522 81574 96534 81626
rect 96586 81574 96598 81626
rect 96650 81574 98808 81626
rect 1104 81552 98808 81574
rect 73798 81472 73804 81524
rect 73856 81512 73862 81524
rect 74166 81512 74172 81524
rect 73856 81484 74172 81512
rect 73856 81472 73862 81484
rect 74166 81472 74172 81484
rect 74224 81512 74230 81524
rect 95234 81512 95240 81524
rect 74224 81484 95240 81512
rect 74224 81472 74230 81484
rect 95234 81472 95240 81484
rect 95292 81472 95298 81524
rect 7006 81336 7012 81388
rect 7064 81376 7070 81388
rect 8202 81376 8208 81388
rect 7064 81348 8208 81376
rect 7064 81336 7070 81348
rect 8202 81336 8208 81348
rect 8260 81336 8266 81388
rect 27801 81311 27859 81317
rect 27801 81308 27813 81311
rect 27632 81280 27813 81308
rect 27632 81184 27660 81280
rect 27801 81277 27813 81280
rect 27847 81277 27859 81311
rect 27801 81271 27859 81277
rect 29825 81243 29883 81249
rect 29825 81209 29837 81243
rect 29871 81240 29883 81243
rect 32490 81240 32496 81252
rect 29871 81212 32496 81240
rect 29871 81209 29883 81212
rect 29825 81203 29883 81209
rect 32490 81200 32496 81212
rect 32548 81200 32554 81252
rect 32582 81200 32588 81252
rect 32640 81240 32646 81252
rect 82449 81243 82507 81249
rect 82449 81240 82461 81243
rect 32640 81212 82461 81240
rect 32640 81200 32646 81212
rect 82449 81209 82461 81212
rect 82495 81240 82507 81243
rect 82725 81243 82783 81249
rect 82725 81240 82737 81243
rect 82495 81212 82737 81240
rect 82495 81209 82507 81212
rect 82449 81203 82507 81209
rect 82725 81209 82737 81212
rect 82771 81209 82783 81243
rect 82725 81203 82783 81209
rect 82998 81200 83004 81252
rect 83056 81240 83062 81252
rect 83093 81243 83151 81249
rect 83093 81240 83105 81243
rect 83056 81212 83105 81240
rect 83056 81200 83062 81212
rect 83093 81209 83105 81212
rect 83139 81240 83151 81243
rect 83642 81240 83648 81252
rect 83139 81212 83648 81240
rect 83139 81209 83151 81212
rect 83093 81203 83151 81209
rect 83642 81200 83648 81212
rect 83700 81200 83706 81252
rect 27614 81172 27620 81184
rect 27575 81144 27620 81172
rect 27614 81132 27620 81144
rect 27672 81132 27678 81184
rect 29914 81172 29920 81184
rect 29875 81144 29920 81172
rect 29914 81132 29920 81144
rect 29972 81132 29978 81184
rect 1104 81082 98808 81104
rect 1104 81030 19606 81082
rect 19658 81030 19670 81082
rect 19722 81030 19734 81082
rect 19786 81030 19798 81082
rect 19850 81030 50326 81082
rect 50378 81030 50390 81082
rect 50442 81030 50454 81082
rect 50506 81030 50518 81082
rect 50570 81030 81046 81082
rect 81098 81030 81110 81082
rect 81162 81030 81174 81082
rect 81226 81030 81238 81082
rect 81290 81030 98808 81082
rect 1104 81008 98808 81030
rect 74074 80900 74080 80912
rect 74035 80872 74080 80900
rect 74074 80860 74080 80872
rect 74132 80860 74138 80912
rect 84286 80900 84292 80912
rect 84247 80872 84292 80900
rect 84286 80860 84292 80872
rect 84344 80860 84350 80912
rect 73893 80835 73951 80841
rect 73893 80801 73905 80835
rect 73939 80801 73951 80835
rect 73893 80795 73951 80801
rect 10226 80588 10232 80640
rect 10284 80628 10290 80640
rect 12894 80628 12900 80640
rect 10284 80600 12900 80628
rect 10284 80588 10290 80600
rect 12894 80588 12900 80600
rect 12952 80588 12958 80640
rect 31386 80588 31392 80640
rect 31444 80628 31450 80640
rect 73617 80631 73675 80637
rect 73617 80628 73629 80631
rect 31444 80600 73629 80628
rect 31444 80588 31450 80600
rect 73617 80597 73629 80600
rect 73663 80628 73675 80631
rect 73908 80628 73936 80795
rect 84378 80724 84384 80776
rect 84436 80724 84442 80776
rect 84654 80764 84660 80776
rect 84615 80736 84660 80764
rect 84654 80724 84660 80736
rect 84712 80724 84718 80776
rect 84396 80696 84424 80724
rect 84565 80699 84623 80705
rect 84565 80696 84577 80699
rect 84396 80668 84577 80696
rect 84565 80665 84577 80668
rect 84611 80665 84623 80699
rect 84565 80659 84623 80665
rect 84470 80637 84476 80640
rect 73663 80600 73936 80628
rect 84454 80631 84476 80637
rect 73663 80597 73675 80600
rect 73617 80591 73675 80597
rect 84454 80597 84466 80631
rect 84454 80591 84476 80597
rect 84470 80588 84476 80591
rect 84528 80588 84534 80640
rect 84746 80628 84752 80640
rect 84707 80600 84752 80628
rect 84746 80588 84752 80600
rect 84804 80588 84810 80640
rect 1104 80538 98808 80560
rect 1104 80486 4246 80538
rect 4298 80486 4310 80538
rect 4362 80486 4374 80538
rect 4426 80486 4438 80538
rect 4490 80486 34966 80538
rect 35018 80486 35030 80538
rect 35082 80486 35094 80538
rect 35146 80486 35158 80538
rect 35210 80486 65686 80538
rect 65738 80486 65750 80538
rect 65802 80486 65814 80538
rect 65866 80486 65878 80538
rect 65930 80486 96406 80538
rect 96458 80486 96470 80538
rect 96522 80486 96534 80538
rect 96586 80486 96598 80538
rect 96650 80486 98808 80538
rect 1104 80464 98808 80486
rect 8202 80248 8208 80300
rect 8260 80288 8266 80300
rect 50249 80291 50307 80297
rect 50249 80288 50261 80291
rect 8260 80260 50261 80288
rect 8260 80248 8266 80260
rect 50249 80257 50261 80260
rect 50295 80257 50307 80291
rect 50249 80251 50307 80257
rect 29089 80223 29147 80229
rect 29089 80189 29101 80223
rect 29135 80189 29147 80223
rect 29089 80183 29147 80189
rect 29365 80223 29423 80229
rect 29365 80189 29377 80223
rect 29411 80220 29423 80223
rect 29638 80220 29644 80232
rect 29411 80192 29644 80220
rect 29411 80189 29423 80192
rect 29365 80183 29423 80189
rect 29104 80084 29132 80183
rect 29638 80180 29644 80192
rect 29696 80180 29702 80232
rect 49602 80220 49608 80232
rect 49563 80192 49608 80220
rect 49602 80180 49608 80192
rect 49660 80180 49666 80232
rect 49786 80220 49792 80232
rect 49747 80192 49792 80220
rect 49786 80180 49792 80192
rect 49844 80180 49850 80232
rect 49973 80223 50031 80229
rect 49973 80189 49985 80223
rect 50019 80220 50031 80223
rect 50062 80220 50068 80232
rect 50019 80192 50068 80220
rect 50019 80189 50031 80192
rect 49973 80183 50031 80189
rect 30834 80152 30840 80164
rect 30024 80124 30840 80152
rect 29362 80084 29368 80096
rect 29104 80056 29368 80084
rect 29362 80044 29368 80056
rect 29420 80084 29426 80096
rect 30024 80084 30052 80124
rect 30834 80112 30840 80124
rect 30892 80112 30898 80164
rect 49694 80112 49700 80164
rect 49752 80152 49758 80164
rect 49988 80152 50016 80183
rect 50062 80180 50068 80192
rect 50120 80180 50126 80232
rect 50154 80180 50160 80232
rect 50212 80220 50218 80232
rect 50341 80223 50399 80229
rect 50341 80220 50353 80223
rect 50212 80192 50353 80220
rect 50212 80180 50218 80192
rect 50341 80189 50353 80192
rect 50387 80189 50399 80223
rect 50341 80183 50399 80189
rect 49752 80124 50016 80152
rect 50356 80152 50384 80183
rect 50706 80152 50712 80164
rect 50356 80124 50712 80152
rect 49752 80112 49758 80124
rect 50706 80112 50712 80124
rect 50764 80112 50770 80164
rect 29420 80056 30052 80084
rect 30653 80087 30711 80093
rect 29420 80044 29426 80056
rect 30653 80053 30665 80087
rect 30699 80084 30711 80087
rect 40770 80084 40776 80096
rect 30699 80056 40776 80084
rect 30699 80053 30711 80056
rect 30653 80047 30711 80053
rect 40770 80044 40776 80056
rect 40828 80084 40834 80096
rect 41322 80084 41328 80096
rect 40828 80056 41328 80084
rect 40828 80044 40834 80056
rect 41322 80044 41328 80056
rect 41380 80044 41386 80096
rect 50798 80084 50804 80096
rect 50759 80056 50804 80084
rect 50798 80044 50804 80056
rect 50856 80044 50862 80096
rect 75638 80044 75644 80096
rect 75696 80084 75702 80096
rect 82170 80084 82176 80096
rect 75696 80056 82176 80084
rect 75696 80044 75702 80056
rect 82170 80044 82176 80056
rect 82228 80044 82234 80096
rect 1104 79994 98808 80016
rect 1104 79942 19606 79994
rect 19658 79942 19670 79994
rect 19722 79942 19734 79994
rect 19786 79942 19798 79994
rect 19850 79942 50326 79994
rect 50378 79942 50390 79994
rect 50442 79942 50454 79994
rect 50506 79942 50518 79994
rect 50570 79942 81046 79994
rect 81098 79942 81110 79994
rect 81162 79942 81174 79994
rect 81226 79942 81238 79994
rect 81290 79942 98808 79994
rect 1104 79920 98808 79942
rect 31018 79840 31024 79892
rect 31076 79880 31082 79892
rect 31076 79852 42932 79880
rect 31076 79840 31082 79852
rect 42904 79824 42932 79852
rect 42886 79812 42892 79824
rect 38626 79784 42748 79812
rect 42799 79784 42892 79812
rect 29178 79704 29184 79756
rect 29236 79744 29242 79756
rect 38626 79744 38654 79784
rect 42610 79744 42616 79756
rect 29236 79716 38654 79744
rect 42571 79716 42616 79744
rect 29236 79704 29242 79716
rect 42610 79704 42616 79716
rect 42668 79704 42674 79756
rect 42720 79744 42748 79784
rect 42886 79772 42892 79784
rect 42944 79772 42950 79824
rect 84166 79784 89484 79812
rect 42797 79747 42855 79753
rect 42797 79744 42809 79747
rect 42720 79716 42809 79744
rect 42797 79713 42809 79716
rect 42843 79713 42855 79747
rect 42797 79707 42855 79713
rect 42986 79747 43044 79753
rect 42986 79713 42998 79747
rect 43032 79713 43044 79747
rect 42986 79707 43044 79713
rect 30466 79636 30472 79688
rect 30524 79676 30530 79688
rect 42628 79676 42656 79704
rect 30524 79648 42656 79676
rect 30524 79636 30530 79648
rect 3970 79500 3976 79552
rect 4028 79540 4034 79552
rect 29178 79540 29184 79552
rect 4028 79512 29184 79540
rect 4028 79500 4034 79512
rect 29178 79500 29184 79512
rect 29236 79500 29242 79552
rect 30374 79500 30380 79552
rect 30432 79540 30438 79552
rect 42521 79543 42579 79549
rect 42521 79540 42533 79543
rect 30432 79512 42533 79540
rect 30432 79500 30438 79512
rect 42521 79509 42533 79512
rect 42567 79540 42579 79543
rect 42996 79540 43024 79707
rect 43162 79704 43168 79756
rect 43220 79753 43226 79756
rect 43220 79747 43240 79753
rect 43228 79713 43240 79747
rect 76466 79744 76472 79756
rect 43220 79707 43240 79713
rect 48286 79716 76472 79744
rect 43220 79704 43226 79707
rect 48286 79676 48314 79716
rect 76466 79704 76472 79716
rect 76524 79704 76530 79756
rect 43180 79648 48314 79676
rect 43180 79608 43208 79648
rect 78122 79636 78128 79688
rect 78180 79676 78186 79688
rect 84166 79676 84194 79784
rect 89073 79747 89131 79753
rect 89073 79713 89085 79747
rect 89119 79713 89131 79747
rect 89073 79707 89131 79713
rect 78180 79648 84194 79676
rect 78180 79636 78186 79648
rect 43088 79580 43208 79608
rect 43088 79540 43116 79580
rect 46290 79568 46296 79620
rect 46348 79608 46354 79620
rect 62114 79608 62120 79620
rect 46348 79580 62120 79608
rect 46348 79568 46354 79580
rect 62114 79568 62120 79580
rect 62172 79568 62178 79620
rect 80790 79568 80796 79620
rect 80848 79608 80854 79620
rect 89088 79608 89116 79707
rect 89162 79704 89168 79756
rect 89220 79753 89226 79756
rect 89456 79753 89484 79784
rect 89220 79747 89279 79753
rect 89220 79713 89233 79747
rect 89267 79713 89279 79747
rect 89220 79707 89279 79713
rect 89441 79747 89499 79753
rect 89441 79713 89453 79747
rect 89487 79713 89499 79747
rect 89622 79744 89628 79756
rect 89583 79716 89628 79744
rect 89441 79707 89499 79713
rect 89220 79704 89226 79707
rect 89622 79704 89628 79716
rect 89680 79704 89686 79756
rect 89346 79676 89352 79688
rect 89307 79648 89352 79676
rect 89346 79636 89352 79648
rect 89404 79636 89410 79688
rect 89806 79608 89812 79620
rect 80848 79580 89116 79608
rect 89767 79580 89812 79608
rect 80848 79568 80854 79580
rect 89806 79568 89812 79580
rect 89864 79568 89870 79620
rect 43438 79540 43444 79552
rect 42567 79512 43116 79540
rect 43351 79512 43444 79540
rect 42567 79509 42579 79512
rect 42521 79503 42579 79509
rect 43438 79500 43444 79512
rect 43496 79540 43502 79552
rect 76006 79540 76012 79552
rect 43496 79512 76012 79540
rect 43496 79500 43502 79512
rect 76006 79500 76012 79512
rect 76064 79500 76070 79552
rect 88981 79543 89039 79549
rect 88981 79509 88993 79543
rect 89027 79540 89039 79543
rect 89162 79540 89168 79552
rect 89027 79512 89168 79540
rect 89027 79509 89039 79512
rect 88981 79503 89039 79509
rect 89162 79500 89168 79512
rect 89220 79500 89226 79552
rect 89346 79500 89352 79552
rect 89404 79540 89410 79552
rect 89901 79543 89959 79549
rect 89901 79540 89913 79543
rect 89404 79512 89913 79540
rect 89404 79500 89410 79512
rect 89901 79509 89913 79512
rect 89947 79509 89959 79543
rect 89901 79503 89959 79509
rect 1104 79450 98808 79472
rect 1104 79398 4246 79450
rect 4298 79398 4310 79450
rect 4362 79398 4374 79450
rect 4426 79398 4438 79450
rect 4490 79398 34966 79450
rect 35018 79398 35030 79450
rect 35082 79398 35094 79450
rect 35146 79398 35158 79450
rect 35210 79398 65686 79450
rect 65738 79398 65750 79450
rect 65802 79398 65814 79450
rect 65866 79398 65878 79450
rect 65930 79398 96406 79450
rect 96458 79398 96470 79450
rect 96522 79398 96534 79450
rect 96586 79398 96598 79450
rect 96650 79398 98808 79450
rect 1104 79376 98808 79398
rect 6822 79336 6828 79348
rect 4080 79308 6828 79336
rect 4080 79209 4108 79308
rect 6822 79296 6828 79308
rect 6880 79336 6886 79348
rect 82814 79336 82820 79348
rect 6880 79308 82820 79336
rect 6880 79296 6886 79308
rect 82814 79296 82820 79308
rect 82872 79296 82878 79348
rect 10318 79228 10324 79280
rect 10376 79268 10382 79280
rect 30374 79268 30380 79280
rect 10376 79240 30380 79268
rect 10376 79228 10382 79240
rect 30374 79228 30380 79240
rect 30432 79228 30438 79280
rect 3237 79203 3295 79209
rect 3237 79169 3249 79203
rect 3283 79200 3295 79203
rect 4065 79203 4123 79209
rect 4065 79200 4077 79203
rect 3283 79172 4077 79200
rect 3283 79169 3295 79172
rect 3237 79163 3295 79169
rect 4065 79169 4077 79172
rect 4111 79169 4123 79203
rect 4065 79163 4123 79169
rect 4433 79203 4491 79209
rect 4433 79169 4445 79203
rect 4479 79200 4491 79203
rect 6270 79200 6276 79212
rect 4479 79172 6276 79200
rect 4479 79169 4491 79172
rect 4433 79163 4491 79169
rect 6270 79160 6276 79172
rect 6328 79160 6334 79212
rect 12894 79160 12900 79212
rect 12952 79200 12958 79212
rect 30466 79200 30472 79212
rect 12952 79172 30472 79200
rect 12952 79160 12958 79172
rect 30466 79160 30472 79172
rect 30524 79160 30530 79212
rect 86218 79160 86224 79212
rect 86276 79200 86282 79212
rect 97353 79203 97411 79209
rect 97353 79200 97365 79203
rect 86276 79172 97365 79200
rect 86276 79160 86282 79172
rect 97353 79169 97365 79172
rect 97399 79169 97411 79203
rect 97353 79163 97411 79169
rect 3970 79132 3976 79144
rect 3931 79104 3976 79132
rect 3970 79092 3976 79104
rect 4028 79092 4034 79144
rect 4341 79135 4399 79141
rect 4341 79101 4353 79135
rect 4387 79132 4399 79135
rect 4522 79132 4528 79144
rect 4387 79104 4528 79132
rect 4387 79101 4399 79104
rect 4341 79095 4399 79101
rect 4522 79092 4528 79104
rect 4580 79092 4586 79144
rect 4706 79132 4712 79144
rect 4667 79104 4712 79132
rect 4706 79092 4712 79104
rect 4764 79092 4770 79144
rect 28169 79135 28227 79141
rect 28169 79101 28181 79135
rect 28215 79132 28227 79135
rect 28445 79135 28503 79141
rect 28445 79132 28457 79135
rect 28215 79104 28457 79132
rect 28215 79101 28227 79104
rect 28169 79095 28227 79101
rect 28445 79101 28457 79104
rect 28491 79132 28503 79135
rect 28534 79132 28540 79144
rect 28491 79104 28540 79132
rect 28491 79101 28503 79104
rect 28445 79095 28503 79101
rect 28534 79092 28540 79104
rect 28592 79092 28598 79144
rect 62114 79092 62120 79144
rect 62172 79132 62178 79144
rect 62850 79132 62856 79144
rect 62172 79104 62856 79132
rect 62172 79092 62178 79104
rect 62850 79092 62856 79104
rect 62908 79132 62914 79144
rect 96709 79135 96767 79141
rect 96709 79132 96721 79135
rect 62908 79104 96721 79132
rect 62908 79092 62914 79104
rect 96709 79101 96721 79104
rect 96755 79101 96767 79135
rect 96890 79132 96896 79144
rect 96851 79104 96896 79132
rect 96709 79095 96767 79101
rect 96890 79092 96896 79104
rect 96948 79092 96954 79144
rect 97074 79132 97080 79144
rect 97035 79104 97080 79132
rect 97074 79092 97080 79104
rect 97132 79092 97138 79144
rect 97442 79132 97448 79144
rect 97403 79104 97448 79132
rect 97442 79092 97448 79104
rect 97500 79092 97506 79144
rect 3421 79067 3479 79073
rect 3421 79033 3433 79067
rect 3467 79064 3479 79067
rect 83090 79064 83096 79076
rect 3467 79036 83096 79064
rect 3467 79033 3479 79036
rect 3421 79027 3479 79033
rect 83090 79024 83096 79036
rect 83148 79024 83154 79076
rect 11606 78956 11612 79008
rect 11664 78996 11670 79008
rect 97905 78999 97963 79005
rect 97905 78996 97917 78999
rect 11664 78968 97917 78996
rect 11664 78956 11670 78968
rect 97905 78965 97917 78968
rect 97951 78965 97963 78999
rect 97905 78959 97963 78965
rect 1104 78906 98808 78928
rect 1104 78854 19606 78906
rect 19658 78854 19670 78906
rect 19722 78854 19734 78906
rect 19786 78854 19798 78906
rect 19850 78854 50326 78906
rect 50378 78854 50390 78906
rect 50442 78854 50454 78906
rect 50506 78854 50518 78906
rect 50570 78854 81046 78906
rect 81098 78854 81110 78906
rect 81162 78854 81174 78906
rect 81226 78854 81238 78906
rect 81290 78854 98808 78906
rect 1104 78832 98808 78854
rect 4706 78752 4712 78804
rect 4764 78792 4770 78804
rect 20714 78792 20720 78804
rect 4764 78764 20720 78792
rect 4764 78752 4770 78764
rect 20714 78752 20720 78764
rect 20772 78752 20778 78804
rect 25774 78752 25780 78804
rect 25832 78792 25838 78804
rect 25832 78764 30788 78792
rect 25832 78752 25838 78764
rect 17052 78696 17540 78724
rect 17052 78668 17080 78696
rect 11057 78659 11115 78665
rect 11057 78625 11069 78659
rect 11103 78656 11115 78659
rect 11514 78656 11520 78668
rect 11103 78628 11520 78656
rect 11103 78625 11115 78628
rect 11057 78619 11115 78625
rect 11514 78616 11520 78628
rect 11572 78616 11578 78668
rect 17034 78616 17040 78668
rect 17092 78616 17098 78668
rect 17126 78616 17132 78668
rect 17184 78656 17190 78668
rect 17512 78665 17540 78696
rect 17586 78684 17592 78736
rect 17644 78724 17650 78736
rect 30760 78733 30788 78764
rect 30745 78727 30803 78733
rect 17644 78696 18184 78724
rect 17644 78684 17650 78696
rect 17770 78665 17776 78668
rect 17313 78659 17371 78665
rect 17313 78656 17325 78659
rect 17184 78628 17325 78656
rect 17184 78616 17190 78628
rect 17313 78625 17325 78628
rect 17359 78625 17371 78659
rect 17313 78619 17371 78625
rect 17497 78659 17555 78665
rect 17497 78625 17509 78659
rect 17543 78625 17555 78659
rect 17497 78619 17555 78625
rect 17717 78659 17776 78665
rect 17717 78625 17729 78659
rect 17763 78625 17776 78659
rect 17717 78619 17776 78625
rect 17770 78616 17776 78619
rect 17828 78616 17834 78668
rect 17865 78659 17923 78665
rect 17865 78625 17877 78659
rect 17911 78656 17923 78659
rect 17911 78628 18000 78656
rect 17911 78625 17923 78628
rect 17865 78619 17923 78625
rect 11241 78591 11299 78597
rect 11241 78557 11253 78591
rect 11287 78588 11299 78591
rect 17402 78588 17408 78600
rect 11287 78560 17408 78588
rect 11287 78557 11299 78560
rect 11241 78551 11299 78557
rect 17402 78548 17408 78560
rect 17460 78548 17466 78600
rect 17589 78591 17647 78597
rect 17589 78588 17601 78591
rect 17512 78560 17601 78588
rect 3878 78480 3884 78532
rect 3936 78520 3942 78532
rect 17512 78520 17540 78560
rect 17589 78557 17601 78560
rect 17635 78557 17647 78591
rect 17589 78551 17647 78557
rect 3936 78492 17540 78520
rect 17972 78520 18000 78628
rect 18156 78588 18184 78696
rect 30300 78696 30604 78724
rect 24026 78616 24032 78668
rect 24084 78656 24090 78668
rect 30300 78656 30328 78696
rect 30466 78656 30472 78668
rect 24084 78628 30328 78656
rect 30427 78628 30472 78656
rect 24084 78616 24090 78628
rect 30466 78616 30472 78628
rect 30524 78616 30530 78668
rect 30576 78656 30604 78696
rect 30745 78693 30757 78727
rect 30791 78693 30803 78727
rect 30745 78687 30803 78693
rect 30653 78659 30711 78665
rect 30653 78656 30665 78659
rect 30576 78628 30665 78656
rect 30653 78625 30665 78628
rect 30699 78625 30711 78659
rect 30653 78619 30711 78625
rect 30842 78659 30900 78665
rect 30842 78625 30854 78659
rect 30888 78625 30900 78659
rect 30842 78619 30900 78625
rect 27890 78588 27896 78600
rect 18156 78560 27896 78588
rect 27890 78548 27896 78560
rect 27948 78548 27954 78600
rect 30374 78588 30380 78600
rect 30335 78560 30380 78588
rect 30374 78548 30380 78560
rect 30432 78588 30438 78600
rect 30852 78588 30880 78619
rect 82722 78616 82728 78668
rect 82780 78656 82786 78668
rect 83093 78659 83151 78665
rect 83093 78656 83105 78659
rect 82780 78628 83105 78656
rect 82780 78616 82786 78628
rect 83093 78625 83105 78628
rect 83139 78656 83151 78659
rect 97994 78656 98000 78668
rect 83139 78628 98000 78656
rect 83139 78625 83151 78628
rect 83093 78619 83151 78625
rect 97994 78616 98000 78628
rect 98052 78616 98058 78668
rect 30432 78560 30880 78588
rect 30432 78548 30438 78560
rect 66070 78548 66076 78600
rect 66128 78588 66134 78600
rect 83277 78591 83335 78597
rect 83277 78588 83289 78591
rect 66128 78560 83289 78588
rect 66128 78548 66134 78560
rect 83277 78557 83289 78560
rect 83323 78557 83335 78591
rect 83277 78551 83335 78557
rect 18049 78523 18107 78529
rect 18049 78520 18061 78523
rect 17972 78492 18061 78520
rect 3936 78480 3942 78492
rect 18049 78489 18061 78492
rect 18095 78520 18107 78523
rect 49050 78520 49056 78532
rect 18095 78492 49056 78520
rect 18095 78489 18107 78492
rect 18049 78483 18107 78489
rect 49050 78480 49056 78492
rect 49108 78480 49114 78532
rect 17034 78452 17040 78464
rect 16995 78424 17040 78452
rect 17034 78412 17040 78424
rect 17092 78412 17098 78464
rect 17218 78452 17224 78464
rect 17179 78424 17224 78452
rect 17218 78412 17224 78424
rect 17276 78412 17282 78464
rect 31021 78455 31079 78461
rect 31021 78421 31033 78455
rect 31067 78452 31079 78455
rect 31110 78452 31116 78464
rect 31067 78424 31116 78452
rect 31067 78421 31079 78424
rect 31021 78415 31079 78421
rect 31110 78412 31116 78424
rect 31168 78412 31174 78464
rect 84289 78455 84347 78461
rect 84289 78421 84301 78455
rect 84335 78452 84347 78455
rect 84565 78455 84623 78461
rect 84565 78452 84577 78455
rect 84335 78424 84577 78452
rect 84335 78421 84347 78424
rect 84289 78415 84347 78421
rect 84565 78421 84577 78424
rect 84611 78452 84623 78455
rect 90358 78452 90364 78464
rect 84611 78424 90364 78452
rect 84611 78421 84623 78424
rect 84565 78415 84623 78421
rect 90358 78412 90364 78424
rect 90416 78412 90422 78464
rect 1104 78362 98808 78384
rect 1104 78310 4246 78362
rect 4298 78310 4310 78362
rect 4362 78310 4374 78362
rect 4426 78310 4438 78362
rect 4490 78310 34966 78362
rect 35018 78310 35030 78362
rect 35082 78310 35094 78362
rect 35146 78310 35158 78362
rect 35210 78310 65686 78362
rect 65738 78310 65750 78362
rect 65802 78310 65814 78362
rect 65866 78310 65878 78362
rect 65930 78310 96406 78362
rect 96458 78310 96470 78362
rect 96522 78310 96534 78362
rect 96586 78310 96598 78362
rect 96650 78310 98808 78362
rect 1104 78288 98808 78310
rect 66162 78208 66168 78260
rect 66220 78248 66226 78260
rect 66220 78220 82952 78248
rect 66220 78208 66226 78220
rect 11514 78140 11520 78192
rect 11572 78180 11578 78192
rect 58618 78180 58624 78192
rect 11572 78152 58624 78180
rect 11572 78140 11578 78152
rect 58618 78140 58624 78152
rect 58676 78140 58682 78192
rect 17034 78072 17040 78124
rect 17092 78112 17098 78124
rect 48958 78112 48964 78124
rect 17092 78084 48964 78112
rect 17092 78072 17098 78084
rect 48958 78072 48964 78084
rect 49016 78072 49022 78124
rect 23385 78047 23443 78053
rect 23385 78013 23397 78047
rect 23431 78044 23443 78047
rect 23658 78044 23664 78056
rect 23431 78016 23664 78044
rect 23431 78013 23443 78016
rect 23385 78007 23443 78013
rect 23658 78004 23664 78016
rect 23716 78004 23722 78056
rect 78401 78047 78459 78053
rect 78401 78044 78413 78047
rect 77312 78016 78413 78044
rect 77021 77979 77079 77985
rect 77021 77976 77033 77979
rect 64846 77948 77033 77976
rect 50890 77868 50896 77920
rect 50948 77908 50954 77920
rect 53650 77908 53656 77920
rect 50948 77880 53656 77908
rect 50948 77868 50954 77880
rect 53650 77868 53656 77880
rect 53708 77908 53714 77920
rect 64846 77908 64874 77948
rect 77021 77945 77033 77948
rect 77067 77945 77079 77979
rect 77021 77939 77079 77945
rect 53708 77880 64874 77908
rect 53708 77868 53714 77880
rect 76742 77868 76748 77920
rect 76800 77908 76806 77920
rect 76837 77911 76895 77917
rect 76837 77908 76849 77911
rect 76800 77880 76849 77908
rect 76800 77868 76806 77880
rect 76837 77877 76849 77880
rect 76883 77908 76895 77911
rect 77312 77908 77340 78016
rect 78401 78013 78413 78016
rect 78447 78013 78459 78047
rect 78401 78007 78459 78013
rect 78677 78047 78735 78053
rect 78677 78013 78689 78047
rect 78723 78044 78735 78047
rect 82722 78044 82728 78056
rect 78723 78016 82400 78044
rect 82683 78016 82728 78044
rect 78723 78013 78735 78016
rect 78677 78007 78735 78013
rect 82262 77976 82268 77988
rect 82223 77948 82268 77976
rect 82262 77936 82268 77948
rect 82320 77936 82326 77988
rect 82372 77976 82400 78016
rect 82722 78004 82728 78016
rect 82780 78004 82786 78056
rect 82924 78053 82952 78220
rect 82909 78047 82967 78053
rect 82909 78013 82921 78047
rect 82955 78013 82967 78047
rect 83090 78044 83096 78056
rect 83051 78016 83096 78044
rect 82909 78007 82967 78013
rect 83090 78004 83096 78016
rect 83148 78004 83154 78056
rect 84194 77976 84200 77988
rect 82372 77948 84200 77976
rect 84194 77936 84200 77948
rect 84252 77976 84258 77988
rect 84562 77976 84568 77988
rect 84252 77948 84568 77976
rect 84252 77936 84258 77948
rect 84562 77936 84568 77948
rect 84620 77976 84626 77988
rect 92566 77976 92572 77988
rect 84620 77948 92572 77976
rect 84620 77936 84626 77948
rect 92566 77936 92572 77948
rect 92624 77936 92630 77988
rect 76883 77880 77340 77908
rect 76883 77877 76895 77880
rect 76837 77871 76895 77877
rect 1104 77818 98808 77840
rect 1104 77766 19606 77818
rect 19658 77766 19670 77818
rect 19722 77766 19734 77818
rect 19786 77766 19798 77818
rect 19850 77766 50326 77818
rect 50378 77766 50390 77818
rect 50442 77766 50454 77818
rect 50506 77766 50518 77818
rect 50570 77766 81046 77818
rect 81098 77766 81110 77818
rect 81162 77766 81174 77818
rect 81226 77766 81238 77818
rect 81290 77766 98808 77818
rect 1104 77744 98808 77766
rect 28442 77704 28448 77716
rect 26344 77676 28448 77704
rect 20714 77636 20720 77648
rect 20675 77608 20720 77636
rect 20714 77596 20720 77608
rect 20772 77596 20778 77648
rect 25958 77568 25964 77580
rect 25919 77540 25964 77568
rect 25958 77528 25964 77540
rect 26016 77528 26022 77580
rect 26142 77528 26148 77580
rect 26200 77568 26206 77580
rect 26344 77577 26372 77676
rect 28442 77664 28448 77676
rect 28500 77664 28506 77716
rect 61378 77664 61384 77716
rect 61436 77704 61442 77716
rect 62758 77704 62764 77716
rect 61436 77676 62764 77704
rect 61436 77664 61442 77676
rect 62758 77664 62764 77676
rect 62816 77704 62822 77716
rect 83090 77704 83096 77716
rect 62816 77676 83096 77704
rect 62816 77664 62822 77676
rect 83090 77664 83096 77676
rect 83148 77664 83154 77716
rect 96798 77636 96804 77648
rect 26436 77608 96804 77636
rect 26329 77571 26387 77577
rect 26200 77540 26244 77568
rect 26200 77528 26206 77540
rect 26329 77537 26341 77571
rect 26375 77537 26387 77571
rect 26329 77531 26387 77537
rect 21545 77503 21603 77509
rect 21545 77469 21557 77503
rect 21591 77500 21603 77503
rect 23382 77500 23388 77512
rect 21591 77472 23388 77500
rect 21591 77469 21603 77472
rect 21545 77463 21603 77469
rect 23382 77460 23388 77472
rect 23440 77460 23446 77512
rect 26237 77503 26295 77509
rect 26237 77469 26249 77503
rect 26283 77469 26295 77503
rect 26237 77463 26295 77469
rect 26252 77432 26280 77463
rect 26436 77432 26464 77608
rect 96798 77596 96804 77608
rect 96856 77596 96862 77648
rect 26510 77528 26516 77580
rect 26568 77568 26574 77580
rect 93762 77568 93768 77580
rect 26568 77540 93768 77568
rect 26568 77528 26574 77540
rect 93762 77528 93768 77540
rect 93820 77528 93826 77580
rect 26252 77404 26464 77432
rect 25869 77367 25927 77373
rect 25869 77333 25881 77367
rect 25915 77364 25927 77367
rect 26418 77364 26424 77376
rect 25915 77336 26424 77364
rect 25915 77333 25927 77336
rect 25869 77327 25927 77333
rect 26418 77324 26424 77336
rect 26476 77324 26482 77376
rect 26602 77364 26608 77376
rect 26563 77336 26608 77364
rect 26602 77324 26608 77336
rect 26660 77324 26666 77376
rect 1104 77274 98808 77296
rect 1104 77222 4246 77274
rect 4298 77222 4310 77274
rect 4362 77222 4374 77274
rect 4426 77222 4438 77274
rect 4490 77222 34966 77274
rect 35018 77222 35030 77274
rect 35082 77222 35094 77274
rect 35146 77222 35158 77274
rect 35210 77222 65686 77274
rect 65738 77222 65750 77274
rect 65802 77222 65814 77274
rect 65866 77222 65878 77274
rect 65930 77222 96406 77274
rect 96458 77222 96470 77274
rect 96522 77222 96534 77274
rect 96586 77222 96598 77274
rect 96650 77222 98808 77274
rect 1104 77200 98808 77222
rect 23382 77120 23388 77172
rect 23440 77160 23446 77172
rect 28261 77163 28319 77169
rect 28261 77160 28273 77163
rect 23440 77132 28273 77160
rect 23440 77120 23446 77132
rect 28261 77129 28273 77132
rect 28307 77129 28319 77163
rect 28261 77123 28319 77129
rect 20714 77092 20720 77104
rect 20675 77064 20720 77092
rect 20714 77052 20720 77064
rect 20772 77052 20778 77104
rect 28276 77092 28304 77123
rect 36354 77120 36360 77172
rect 36412 77160 36418 77172
rect 43257 77163 43315 77169
rect 43257 77160 43269 77163
rect 36412 77132 43269 77160
rect 36412 77120 36418 77132
rect 43257 77129 43269 77132
rect 43303 77160 43315 77163
rect 43349 77163 43407 77169
rect 43349 77160 43361 77163
rect 43303 77132 43361 77160
rect 43303 77129 43315 77132
rect 43257 77123 43315 77129
rect 43349 77129 43361 77132
rect 43395 77129 43407 77163
rect 43349 77123 43407 77129
rect 80790 77092 80796 77104
rect 28276 77064 80796 77092
rect 28276 76956 28304 77064
rect 80790 77052 80796 77064
rect 80848 77052 80854 77104
rect 78122 77024 78128 77036
rect 29196 76996 78128 77024
rect 29196 76968 29224 76996
rect 78122 76984 78128 76996
rect 78180 76984 78186 77036
rect 28445 76959 28503 76965
rect 28445 76956 28457 76959
rect 28276 76928 28457 76956
rect 28445 76925 28457 76928
rect 28491 76925 28503 76959
rect 28445 76919 28503 76925
rect 28629 76959 28687 76965
rect 28629 76925 28641 76959
rect 28675 76925 28687 76959
rect 28810 76956 28816 76968
rect 28771 76928 28816 76956
rect 28629 76919 28687 76925
rect 20533 76891 20591 76897
rect 20533 76857 20545 76891
rect 20579 76857 20591 76891
rect 20533 76851 20591 76857
rect 20548 76820 20576 76851
rect 21358 76848 21364 76900
rect 21416 76888 21422 76900
rect 28644 76888 28672 76919
rect 28810 76916 28816 76928
rect 28868 76916 28874 76968
rect 29178 76956 29184 76968
rect 29139 76928 29184 76956
rect 29178 76916 29184 76928
rect 29236 76916 29242 76968
rect 29362 76956 29368 76968
rect 29323 76928 29368 76956
rect 29362 76916 29368 76928
rect 29420 76916 29426 76968
rect 43257 76959 43315 76965
rect 43257 76925 43269 76959
rect 43303 76956 43315 76959
rect 43533 76959 43591 76965
rect 43533 76956 43545 76959
rect 43303 76928 43545 76956
rect 43303 76925 43315 76928
rect 43257 76919 43315 76925
rect 43533 76925 43545 76928
rect 43579 76925 43591 76959
rect 43806 76956 43812 76968
rect 43767 76928 43812 76956
rect 43533 76919 43591 76925
rect 43806 76916 43812 76928
rect 43864 76916 43870 76968
rect 54205 76959 54263 76965
rect 54205 76925 54217 76959
rect 54251 76956 54263 76959
rect 54478 76956 54484 76968
rect 54251 76928 54484 76956
rect 54251 76925 54263 76928
rect 54205 76919 54263 76925
rect 54478 76916 54484 76928
rect 54536 76916 54542 76968
rect 93121 76959 93179 76965
rect 93121 76925 93133 76959
rect 93167 76925 93179 76959
rect 93121 76919 93179 76925
rect 32582 76888 32588 76900
rect 21416 76860 28672 76888
rect 28736 76860 32588 76888
rect 21416 76848 21422 76860
rect 21266 76820 21272 76832
rect 20548 76792 21272 76820
rect 21266 76780 21272 76792
rect 21324 76820 21330 76832
rect 28736 76820 28764 76860
rect 32582 76848 32588 76860
rect 32640 76848 32646 76900
rect 29638 76820 29644 76832
rect 21324 76792 28764 76820
rect 29599 76792 29644 76820
rect 21324 76780 21330 76792
rect 29638 76780 29644 76792
rect 29696 76780 29702 76832
rect 79410 76780 79416 76832
rect 79468 76820 79474 76832
rect 92937 76823 92995 76829
rect 92937 76820 92949 76823
rect 79468 76792 92949 76820
rect 79468 76780 79474 76792
rect 92937 76789 92949 76792
rect 92983 76820 92995 76823
rect 93136 76820 93164 76919
rect 92983 76792 93164 76820
rect 92983 76789 92995 76792
rect 92937 76783 92995 76789
rect 1104 76730 98808 76752
rect 1104 76678 19606 76730
rect 19658 76678 19670 76730
rect 19722 76678 19734 76730
rect 19786 76678 19798 76730
rect 19850 76678 50326 76730
rect 50378 76678 50390 76730
rect 50442 76678 50454 76730
rect 50506 76678 50518 76730
rect 50570 76678 81046 76730
rect 81098 76678 81110 76730
rect 81162 76678 81174 76730
rect 81226 76678 81238 76730
rect 81290 76678 98808 76730
rect 1104 76656 98808 76678
rect 24486 76576 24492 76628
rect 24544 76616 24550 76628
rect 55582 76616 55588 76628
rect 24544 76588 55588 76616
rect 24544 76576 24550 76588
rect 55582 76576 55588 76588
rect 55640 76616 55646 76628
rect 56226 76616 56232 76628
rect 55640 76588 56232 76616
rect 55640 76576 55646 76588
rect 56226 76576 56232 76588
rect 56284 76576 56290 76628
rect 58066 76616 58072 76628
rect 58027 76588 58072 76616
rect 58066 76576 58072 76588
rect 58124 76616 58130 76628
rect 58342 76616 58348 76628
rect 58124 76588 58348 76616
rect 58124 76576 58130 76588
rect 58342 76576 58348 76588
rect 58400 76576 58406 76628
rect 71774 76508 71780 76560
rect 71832 76548 71838 76560
rect 72510 76548 72516 76560
rect 71832 76520 72516 76548
rect 71832 76508 71838 76520
rect 72510 76508 72516 76520
rect 72568 76548 72574 76560
rect 79778 76548 79784 76560
rect 72568 76520 79784 76548
rect 72568 76508 72574 76520
rect 79778 76508 79784 76520
rect 79836 76508 79842 76560
rect 3326 76440 3332 76492
rect 3384 76480 3390 76492
rect 21358 76480 21364 76492
rect 3384 76452 21364 76480
rect 3384 76440 3390 76452
rect 21358 76440 21364 76452
rect 21416 76440 21422 76492
rect 25593 76483 25651 76489
rect 25593 76449 25605 76483
rect 25639 76480 25651 76483
rect 26145 76483 26203 76489
rect 26145 76480 26157 76483
rect 25639 76452 26157 76480
rect 25639 76449 25651 76452
rect 25593 76443 25651 76449
rect 26145 76449 26157 76452
rect 26191 76449 26203 76483
rect 30558 76480 30564 76492
rect 30471 76452 30564 76480
rect 26145 76443 26203 76449
rect 30558 76440 30564 76452
rect 30616 76480 30622 76492
rect 31386 76480 31392 76492
rect 30616 76452 31392 76480
rect 30616 76440 30622 76452
rect 31386 76440 31392 76452
rect 31444 76440 31450 76492
rect 47670 76440 47676 76492
rect 47728 76480 47734 76492
rect 56965 76483 57023 76489
rect 56965 76480 56977 76483
rect 47728 76452 56977 76480
rect 47728 76440 47734 76452
rect 56965 76449 56977 76452
rect 57011 76449 57023 76483
rect 56965 76443 57023 76449
rect 93578 76440 93584 76492
rect 93636 76480 93642 76492
rect 94041 76483 94099 76489
rect 94041 76480 94053 76483
rect 93636 76452 94053 76480
rect 93636 76440 93642 76452
rect 94041 76449 94053 76452
rect 94087 76449 94099 76483
rect 94041 76443 94099 76449
rect 13814 76372 13820 76424
rect 13872 76412 13878 76424
rect 15102 76412 15108 76424
rect 13872 76384 15108 76412
rect 13872 76372 13878 76384
rect 15102 76372 15108 76384
rect 15160 76412 15166 76424
rect 25869 76415 25927 76421
rect 25869 76412 25881 76415
rect 15160 76384 25881 76412
rect 15160 76372 15166 76384
rect 25869 76381 25881 76384
rect 25915 76381 25927 76415
rect 31110 76412 31116 76424
rect 31071 76384 31116 76412
rect 25869 76375 25927 76381
rect 31110 76372 31116 76384
rect 31168 76372 31174 76424
rect 56686 76412 56692 76424
rect 56647 76384 56692 76412
rect 56686 76372 56692 76384
rect 56744 76372 56750 76424
rect 92566 76372 92572 76424
rect 92624 76412 92630 76424
rect 93765 76415 93823 76421
rect 93765 76412 93777 76415
rect 92624 76384 93777 76412
rect 92624 76372 92630 76384
rect 93765 76381 93777 76384
rect 93811 76381 93823 76415
rect 93765 76375 93823 76381
rect 24118 76304 24124 76356
rect 24176 76344 24182 76356
rect 24176 76316 25820 76344
rect 24176 76304 24182 76316
rect 8938 76236 8944 76288
rect 8996 76276 9002 76288
rect 25593 76279 25651 76285
rect 25593 76276 25605 76279
rect 8996 76248 25605 76276
rect 8996 76236 9002 76248
rect 25593 76245 25605 76248
rect 25639 76276 25651 76279
rect 25685 76279 25743 76285
rect 25685 76276 25697 76279
rect 25639 76248 25697 76276
rect 25639 76245 25651 76248
rect 25593 76239 25651 76245
rect 25685 76245 25697 76248
rect 25731 76245 25743 76279
rect 25792 76276 25820 76316
rect 27249 76279 27307 76285
rect 27249 76276 27261 76279
rect 25792 76248 27261 76276
rect 25685 76239 25743 76245
rect 27249 76245 27261 76248
rect 27295 76245 27307 76279
rect 27249 76239 27307 76245
rect 37461 76279 37519 76285
rect 37461 76245 37473 76279
rect 37507 76276 37519 76279
rect 37550 76276 37556 76288
rect 37507 76248 37556 76276
rect 37507 76245 37519 76248
rect 37461 76239 37519 76245
rect 37550 76236 37556 76248
rect 37608 76236 37614 76288
rect 93578 76276 93584 76288
rect 93539 76248 93584 76276
rect 93578 76236 93584 76248
rect 93636 76236 93642 76288
rect 95142 76276 95148 76288
rect 95103 76248 95148 76276
rect 95142 76236 95148 76248
rect 95200 76236 95206 76288
rect 1104 76186 98808 76208
rect 1104 76134 4246 76186
rect 4298 76134 4310 76186
rect 4362 76134 4374 76186
rect 4426 76134 4438 76186
rect 4490 76134 34966 76186
rect 35018 76134 35030 76186
rect 35082 76134 35094 76186
rect 35146 76134 35158 76186
rect 35210 76134 65686 76186
rect 65738 76134 65750 76186
rect 65802 76134 65814 76186
rect 65866 76134 65878 76186
rect 65930 76134 96406 76186
rect 96458 76134 96470 76186
rect 96522 76134 96534 76186
rect 96586 76134 96598 76186
rect 96650 76134 98808 76186
rect 1104 76112 98808 76134
rect 56226 76032 56232 76084
rect 56284 76072 56290 76084
rect 95142 76072 95148 76084
rect 56284 76044 95148 76072
rect 56284 76032 56290 76044
rect 95142 76032 95148 76044
rect 95200 76032 95206 76084
rect 4893 76007 4951 76013
rect 4893 75973 4905 76007
rect 4939 76004 4951 76007
rect 5350 76004 5356 76016
rect 4939 75976 5356 76004
rect 4939 75973 4951 75976
rect 4893 75967 4951 75973
rect 5350 75964 5356 75976
rect 5408 75964 5414 76016
rect 44545 75939 44603 75945
rect 44545 75905 44557 75939
rect 44591 75936 44603 75939
rect 71774 75936 71780 75948
rect 44591 75908 71780 75936
rect 44591 75905 44603 75908
rect 44545 75899 44603 75905
rect 71774 75896 71780 75908
rect 71832 75896 71838 75948
rect 5074 75868 5080 75880
rect 5035 75840 5080 75868
rect 5074 75828 5080 75840
rect 5132 75828 5138 75880
rect 5261 75871 5319 75877
rect 5261 75837 5273 75871
rect 5307 75837 5319 75871
rect 5261 75831 5319 75837
rect 5445 75871 5503 75877
rect 5445 75837 5457 75871
rect 5491 75868 5503 75871
rect 15010 75868 15016 75880
rect 5491 75840 15016 75868
rect 5491 75837 5503 75840
rect 5445 75831 5503 75837
rect 5276 75800 5304 75831
rect 15010 75828 15016 75840
rect 15068 75828 15074 75880
rect 30009 75871 30067 75877
rect 30009 75837 30021 75871
rect 30055 75868 30067 75871
rect 35434 75868 35440 75880
rect 30055 75840 35440 75868
rect 30055 75837 30067 75840
rect 30009 75831 30067 75837
rect 35434 75828 35440 75840
rect 35492 75828 35498 75880
rect 38010 75828 38016 75880
rect 38068 75868 38074 75880
rect 38654 75868 38660 75880
rect 38068 75840 38660 75868
rect 38068 75828 38074 75840
rect 38654 75828 38660 75840
rect 38712 75828 38718 75880
rect 44082 75868 44088 75880
rect 44043 75840 44088 75868
rect 44082 75828 44088 75840
rect 44140 75828 44146 75880
rect 9674 75800 9680 75812
rect 5276 75772 9680 75800
rect 9674 75760 9680 75772
rect 9732 75760 9738 75812
rect 30285 75803 30343 75809
rect 30285 75769 30297 75803
rect 30331 75800 30343 75803
rect 30558 75800 30564 75812
rect 30331 75772 30564 75800
rect 30331 75769 30343 75772
rect 30285 75763 30343 75769
rect 30558 75760 30564 75772
rect 30616 75760 30622 75812
rect 1104 75642 98808 75664
rect 1104 75590 19606 75642
rect 19658 75590 19670 75642
rect 19722 75590 19734 75642
rect 19786 75590 19798 75642
rect 19850 75590 50326 75642
rect 50378 75590 50390 75642
rect 50442 75590 50454 75642
rect 50506 75590 50518 75642
rect 50570 75590 81046 75642
rect 81098 75590 81110 75642
rect 81162 75590 81174 75642
rect 81226 75590 81238 75642
rect 81290 75590 98808 75642
rect 1104 75568 98808 75590
rect 57514 75420 57520 75472
rect 57572 75460 57578 75472
rect 68554 75460 68560 75472
rect 57572 75432 68560 75460
rect 57572 75420 57578 75432
rect 68554 75420 68560 75432
rect 68612 75420 68618 75472
rect 12434 75352 12440 75404
rect 12492 75392 12498 75404
rect 12618 75392 12624 75404
rect 12492 75364 12624 75392
rect 12492 75352 12498 75364
rect 12618 75352 12624 75364
rect 12676 75392 12682 75404
rect 43438 75392 43444 75404
rect 12676 75364 43444 75392
rect 12676 75352 12682 75364
rect 43438 75352 43444 75364
rect 43496 75352 43502 75404
rect 54478 75352 54484 75404
rect 54536 75392 54542 75404
rect 94498 75392 94504 75404
rect 54536 75364 94504 75392
rect 54536 75352 54542 75364
rect 94498 75352 94504 75364
rect 94556 75352 94562 75404
rect 17770 75284 17776 75336
rect 17828 75324 17834 75336
rect 68370 75324 68376 75336
rect 17828 75296 68376 75324
rect 17828 75284 17834 75296
rect 68370 75284 68376 75296
rect 68428 75284 68434 75336
rect 28534 75216 28540 75268
rect 28592 75256 28598 75268
rect 87874 75256 87880 75268
rect 28592 75228 87880 75256
rect 28592 75216 28598 75228
rect 87874 75216 87880 75228
rect 87932 75216 87938 75268
rect 25866 75148 25872 75200
rect 25924 75188 25930 75200
rect 91094 75188 91100 75200
rect 25924 75160 91100 75188
rect 25924 75148 25930 75160
rect 91094 75148 91100 75160
rect 91152 75148 91158 75200
rect 93946 75148 93952 75200
rect 94004 75188 94010 75200
rect 94961 75191 95019 75197
rect 94961 75188 94973 75191
rect 94004 75160 94973 75188
rect 94004 75148 94010 75160
rect 94961 75157 94973 75160
rect 95007 75188 95019 75191
rect 95145 75191 95203 75197
rect 95145 75188 95157 75191
rect 95007 75160 95157 75188
rect 95007 75157 95019 75160
rect 94961 75151 95019 75157
rect 95145 75157 95157 75160
rect 95191 75157 95203 75191
rect 95145 75151 95203 75157
rect 1104 75098 98808 75120
rect 1104 75046 4246 75098
rect 4298 75046 4310 75098
rect 4362 75046 4374 75098
rect 4426 75046 4438 75098
rect 4490 75046 34966 75098
rect 35018 75046 35030 75098
rect 35082 75046 35094 75098
rect 35146 75046 35158 75098
rect 35210 75046 65686 75098
rect 65738 75046 65750 75098
rect 65802 75046 65814 75098
rect 65866 75046 65878 75098
rect 65930 75046 96406 75098
rect 96458 75046 96470 75098
rect 96522 75046 96534 75098
rect 96586 75046 96598 75098
rect 96650 75046 98808 75098
rect 1104 75024 98808 75046
rect 2593 74851 2651 74857
rect 2593 74817 2605 74851
rect 2639 74848 2651 74851
rect 13722 74848 13728 74860
rect 2639 74820 13728 74848
rect 2639 74817 2651 74820
rect 2593 74811 2651 74817
rect 13722 74808 13728 74820
rect 13780 74808 13786 74860
rect 72418 74808 72424 74860
rect 72476 74848 72482 74860
rect 72476 74820 73200 74848
rect 72476 74808 72482 74820
rect 2866 74780 2872 74792
rect 2827 74752 2872 74780
rect 2866 74740 2872 74752
rect 2924 74740 2930 74792
rect 72234 74740 72240 74792
rect 72292 74780 72298 74792
rect 72605 74783 72663 74789
rect 72605 74780 72617 74783
rect 72292 74752 72617 74780
rect 72292 74740 72298 74752
rect 72605 74749 72617 74752
rect 72651 74749 72663 74783
rect 72605 74743 72663 74749
rect 72694 74740 72700 74792
rect 72752 74789 72758 74792
rect 72752 74783 72811 74789
rect 72752 74749 72765 74783
rect 72799 74749 72811 74783
rect 72878 74780 72884 74792
rect 72839 74752 72884 74780
rect 72752 74743 72811 74749
rect 72752 74740 72758 74743
rect 72878 74740 72884 74752
rect 72936 74740 72942 74792
rect 72970 74740 72976 74792
rect 73028 74780 73034 74792
rect 73172 74789 73200 74820
rect 73157 74783 73215 74789
rect 73028 74752 73073 74780
rect 73028 74740 73034 74752
rect 73157 74749 73169 74783
rect 73203 74749 73215 74783
rect 73157 74743 73215 74749
rect 77941 74715 77999 74721
rect 77941 74681 77953 74715
rect 77987 74712 77999 74715
rect 79318 74712 79324 74724
rect 77987 74684 79324 74712
rect 77987 74681 77999 74684
rect 77941 74675 77999 74681
rect 79318 74672 79324 74684
rect 79376 74672 79382 74724
rect 4157 74647 4215 74653
rect 4157 74613 4169 74647
rect 4203 74644 4215 74647
rect 12434 74644 12440 74656
rect 4203 74616 12440 74644
rect 4203 74613 4215 74616
rect 4157 74607 4215 74613
rect 12434 74604 12440 74616
rect 12492 74604 12498 74656
rect 44174 74604 44180 74656
rect 44232 74644 44238 74656
rect 73249 74647 73307 74653
rect 73249 74644 73261 74647
rect 44232 74616 73261 74644
rect 44232 74604 44238 74616
rect 73249 74613 73261 74616
rect 73295 74613 73307 74647
rect 73249 74607 73307 74613
rect 78033 74647 78091 74653
rect 78033 74613 78045 74647
rect 78079 74644 78091 74647
rect 78306 74644 78312 74656
rect 78079 74616 78312 74644
rect 78079 74613 78091 74616
rect 78033 74607 78091 74613
rect 78306 74604 78312 74616
rect 78364 74644 78370 74656
rect 97074 74644 97080 74656
rect 78364 74616 97080 74644
rect 78364 74604 78370 74616
rect 97074 74604 97080 74616
rect 97132 74604 97138 74656
rect 1104 74554 98808 74576
rect 1104 74502 19606 74554
rect 19658 74502 19670 74554
rect 19722 74502 19734 74554
rect 19786 74502 19798 74554
rect 19850 74502 50326 74554
rect 50378 74502 50390 74554
rect 50442 74502 50454 74554
rect 50506 74502 50518 74554
rect 50570 74502 81046 74554
rect 81098 74502 81110 74554
rect 81162 74502 81174 74554
rect 81226 74502 81238 74554
rect 81290 74502 98808 74554
rect 1104 74480 98808 74502
rect 32490 74400 32496 74452
rect 32548 74440 32554 74452
rect 44082 74440 44088 74452
rect 32548 74412 44088 74440
rect 32548 74400 32554 74412
rect 44082 74400 44088 74412
rect 44140 74400 44146 74452
rect 53282 74440 53288 74452
rect 51644 74412 53288 74440
rect 51442 74304 51448 74316
rect 51403 74276 51448 74304
rect 51442 74264 51448 74276
rect 51500 74264 51506 74316
rect 51644 74313 51672 74412
rect 53282 74400 53288 74412
rect 53340 74400 53346 74452
rect 53374 74372 53380 74384
rect 51736 74344 53380 74372
rect 51736 74313 51764 74344
rect 53374 74332 53380 74344
rect 53432 74332 53438 74384
rect 76561 74375 76619 74381
rect 76561 74341 76573 74375
rect 76607 74372 76619 74375
rect 76607 74344 84194 74372
rect 76607 74341 76619 74344
rect 76561 74335 76619 74341
rect 51628 74307 51686 74313
rect 51628 74273 51640 74307
rect 51674 74273 51686 74307
rect 51628 74267 51686 74273
rect 51721 74307 51779 74313
rect 51721 74273 51733 74307
rect 51767 74273 51779 74307
rect 51994 74304 52000 74316
rect 51955 74276 52000 74304
rect 51721 74267 51779 74273
rect 51994 74264 52000 74276
rect 52052 74264 52058 74316
rect 56686 74304 56692 74316
rect 56599 74276 56692 74304
rect 56686 74264 56692 74276
rect 56744 74304 56750 74316
rect 61930 74304 61936 74316
rect 56744 74276 61936 74304
rect 56744 74264 56750 74276
rect 61930 74264 61936 74276
rect 61988 74264 61994 74316
rect 78306 74304 78312 74316
rect 78267 74276 78312 74304
rect 78306 74264 78312 74276
rect 78364 74264 78370 74316
rect 51813 74239 51871 74245
rect 51813 74205 51825 74239
rect 51859 74236 51871 74239
rect 52454 74236 52460 74248
rect 51859 74208 52460 74236
rect 51859 74205 51871 74208
rect 51813 74199 51871 74205
rect 52454 74196 52460 74208
rect 52512 74196 52518 74248
rect 56962 74236 56968 74248
rect 56923 74208 56968 74236
rect 56962 74196 56968 74208
rect 57020 74196 57026 74248
rect 78490 74236 78496 74248
rect 78451 74208 78496 74236
rect 78490 74196 78496 74208
rect 78548 74196 78554 74248
rect 84166 74236 84194 74344
rect 96062 74236 96068 74248
rect 84166 74208 96068 74236
rect 96062 74196 96068 74208
rect 96120 74196 96126 74248
rect 41386 74140 55214 74168
rect 25038 74060 25044 74112
rect 25096 74100 25102 74112
rect 26786 74100 26792 74112
rect 25096 74072 26792 74100
rect 25096 74060 25102 74072
rect 26786 74060 26792 74072
rect 26844 74100 26850 74112
rect 41386 74100 41414 74140
rect 52086 74100 52092 74112
rect 26844 74072 41414 74100
rect 52047 74072 52092 74100
rect 26844 74060 26850 74072
rect 52086 74060 52092 74072
rect 52144 74060 52150 74112
rect 55186 74100 55214 74140
rect 58069 74103 58127 74109
rect 58069 74100 58081 74103
rect 55186 74072 58081 74100
rect 58069 74069 58081 74072
rect 58115 74069 58127 74103
rect 58069 74063 58127 74069
rect 1104 74010 98808 74032
rect 1104 73958 4246 74010
rect 4298 73958 4310 74010
rect 4362 73958 4374 74010
rect 4426 73958 4438 74010
rect 4490 73958 34966 74010
rect 35018 73958 35030 74010
rect 35082 73958 35094 74010
rect 35146 73958 35158 74010
rect 35210 73958 65686 74010
rect 65738 73958 65750 74010
rect 65802 73958 65814 74010
rect 65866 73958 65878 74010
rect 65930 73958 96406 74010
rect 96458 73958 96470 74010
rect 96522 73958 96534 74010
rect 96586 73958 96598 74010
rect 96650 73958 98808 74010
rect 1104 73936 98808 73958
rect 16298 73856 16304 73908
rect 16356 73896 16362 73908
rect 17862 73896 17868 73908
rect 16356 73868 17868 73896
rect 16356 73856 16362 73868
rect 17862 73856 17868 73868
rect 17920 73896 17926 73908
rect 25038 73896 25044 73908
rect 17920 73868 25044 73896
rect 17920 73856 17926 73868
rect 25038 73856 25044 73868
rect 25096 73856 25102 73908
rect 39574 73856 39580 73908
rect 39632 73896 39638 73908
rect 56962 73896 56968 73908
rect 39632 73868 56968 73896
rect 39632 73856 39638 73868
rect 56962 73856 56968 73868
rect 57020 73856 57026 73908
rect 26050 73788 26056 73840
rect 26108 73828 26114 73840
rect 38838 73828 38844 73840
rect 26108 73800 38844 73828
rect 26108 73788 26114 73800
rect 38838 73788 38844 73800
rect 38896 73828 38902 73840
rect 39942 73828 39948 73840
rect 38896 73800 39948 73828
rect 38896 73788 38902 73800
rect 39942 73788 39948 73800
rect 40000 73788 40006 73840
rect 45278 73788 45284 73840
rect 45336 73828 45342 73840
rect 52086 73828 52092 73840
rect 45336 73800 52092 73828
rect 45336 73788 45342 73800
rect 52086 73788 52092 73800
rect 52144 73788 52150 73840
rect 24210 73720 24216 73772
rect 24268 73760 24274 73772
rect 78490 73760 78496 73772
rect 24268 73732 78496 73760
rect 24268 73720 24274 73732
rect 78490 73720 78496 73732
rect 78548 73720 78554 73772
rect 44082 73584 44088 73636
rect 44140 73624 44146 73636
rect 76834 73624 76840 73636
rect 44140 73596 76840 73624
rect 44140 73584 44146 73596
rect 76834 73584 76840 73596
rect 76892 73584 76898 73636
rect 76926 73556 76932 73568
rect 76887 73528 76932 73556
rect 76926 73516 76932 73528
rect 76984 73516 76990 73568
rect 1104 73466 98808 73488
rect 1104 73414 19606 73466
rect 19658 73414 19670 73466
rect 19722 73414 19734 73466
rect 19786 73414 19798 73466
rect 19850 73414 50326 73466
rect 50378 73414 50390 73466
rect 50442 73414 50454 73466
rect 50506 73414 50518 73466
rect 50570 73414 81046 73466
rect 81098 73414 81110 73466
rect 81162 73414 81174 73466
rect 81226 73414 81238 73466
rect 81290 73414 98808 73466
rect 1104 73392 98808 73414
rect 39942 73244 39948 73296
rect 40000 73284 40006 73296
rect 76558 73284 76564 73296
rect 40000 73256 76564 73284
rect 40000 73244 40006 73256
rect 76558 73244 76564 73256
rect 76616 73244 76622 73296
rect 27890 73176 27896 73228
rect 27948 73216 27954 73228
rect 46201 73219 46259 73225
rect 46201 73216 46213 73219
rect 27948 73188 46213 73216
rect 27948 73176 27954 73188
rect 46201 73185 46213 73188
rect 46247 73185 46259 73219
rect 46201 73179 46259 73185
rect 47029 73219 47087 73225
rect 47029 73185 47041 73219
rect 47075 73216 47087 73219
rect 70210 73216 70216 73228
rect 47075 73188 70216 73216
rect 47075 73185 47087 73188
rect 47029 73179 47087 73185
rect 70210 73176 70216 73188
rect 70268 73176 70274 73228
rect 43806 73108 43812 73160
rect 43864 73148 43870 73160
rect 48774 73148 48780 73160
rect 43864 73120 48780 73148
rect 43864 73108 43870 73120
rect 48774 73108 48780 73120
rect 48832 73108 48838 73160
rect 1104 72922 98808 72944
rect 1104 72870 4246 72922
rect 4298 72870 4310 72922
rect 4362 72870 4374 72922
rect 4426 72870 4438 72922
rect 4490 72870 34966 72922
rect 35018 72870 35030 72922
rect 35082 72870 35094 72922
rect 35146 72870 35158 72922
rect 35210 72870 65686 72922
rect 65738 72870 65750 72922
rect 65802 72870 65814 72922
rect 65866 72870 65878 72922
rect 65930 72870 96406 72922
rect 96458 72870 96470 72922
rect 96522 72870 96534 72922
rect 96586 72870 96598 72922
rect 96650 72870 98808 72922
rect 1104 72848 98808 72870
rect 84194 72808 84200 72820
rect 82924 72780 84200 72808
rect 13265 72675 13323 72681
rect 13265 72641 13277 72675
rect 13311 72672 13323 72675
rect 13722 72672 13728 72684
rect 13311 72644 13728 72672
rect 13311 72641 13323 72644
rect 13265 72635 13323 72641
rect 13722 72632 13728 72644
rect 13780 72632 13786 72684
rect 82924 72681 82952 72780
rect 84194 72768 84200 72780
rect 84252 72808 84258 72820
rect 84562 72808 84568 72820
rect 84252 72780 84568 72808
rect 84252 72768 84258 72780
rect 84562 72768 84568 72780
rect 84620 72768 84626 72820
rect 82909 72675 82967 72681
rect 82909 72641 82921 72675
rect 82955 72641 82967 72675
rect 82909 72635 82967 72641
rect 13538 72604 13544 72616
rect 13499 72576 13544 72604
rect 13538 72564 13544 72576
rect 13596 72564 13602 72616
rect 78582 72564 78588 72616
rect 78640 72604 78646 72616
rect 83185 72607 83243 72613
rect 83185 72604 83197 72607
rect 78640 72576 83197 72604
rect 78640 72564 78646 72576
rect 83185 72573 83197 72576
rect 83231 72573 83243 72607
rect 83185 72567 83243 72573
rect 50062 72496 50068 72548
rect 50120 72536 50126 72548
rect 50614 72536 50620 72548
rect 50120 72508 50620 72536
rect 50120 72496 50126 72508
rect 50614 72496 50620 72508
rect 50672 72536 50678 72548
rect 59906 72536 59912 72548
rect 50672 72508 59912 72536
rect 50672 72496 50678 72508
rect 59906 72496 59912 72508
rect 59964 72496 59970 72548
rect 82906 72536 82912 72548
rect 74506 72508 82912 72536
rect 74506 72480 74534 72508
rect 82906 72496 82912 72508
rect 82964 72496 82970 72548
rect 13630 72428 13636 72480
rect 13688 72468 13694 72480
rect 14645 72471 14703 72477
rect 14645 72468 14657 72471
rect 13688 72440 14657 72468
rect 13688 72428 13694 72440
rect 14645 72437 14657 72440
rect 14691 72468 14703 72471
rect 74506 72468 74540 72480
rect 14691 72440 74540 72468
rect 14691 72437 14703 72440
rect 14645 72431 14703 72437
rect 74534 72428 74540 72440
rect 74592 72428 74598 72480
rect 79962 72428 79968 72480
rect 80020 72468 80026 72480
rect 84289 72471 84347 72477
rect 84289 72468 84301 72471
rect 80020 72440 84301 72468
rect 80020 72428 80026 72440
rect 84289 72437 84301 72440
rect 84335 72437 84347 72471
rect 84289 72431 84347 72437
rect 1104 72378 98808 72400
rect 1104 72326 19606 72378
rect 19658 72326 19670 72378
rect 19722 72326 19734 72378
rect 19786 72326 19798 72378
rect 19850 72326 50326 72378
rect 50378 72326 50390 72378
rect 50442 72326 50454 72378
rect 50506 72326 50518 72378
rect 50570 72326 81046 72378
rect 81098 72326 81110 72378
rect 81162 72326 81174 72378
rect 81226 72326 81238 72378
rect 81290 72326 98808 72378
rect 1104 72304 98808 72326
rect 1946 72224 1952 72276
rect 2004 72264 2010 72276
rect 30837 72267 30895 72273
rect 30837 72264 30849 72267
rect 2004 72236 30849 72264
rect 2004 72224 2010 72236
rect 30837 72233 30849 72236
rect 30883 72233 30895 72267
rect 30837 72227 30895 72233
rect 9490 72088 9496 72140
rect 9548 72128 9554 72140
rect 9585 72131 9643 72137
rect 9585 72128 9597 72131
rect 9548 72100 9597 72128
rect 9548 72088 9554 72100
rect 9585 72097 9597 72100
rect 9631 72097 9643 72131
rect 30852 72128 30880 72227
rect 50706 72224 50712 72276
rect 50764 72264 50770 72276
rect 79962 72264 79968 72276
rect 50764 72236 60320 72264
rect 50764 72224 50770 72236
rect 48774 72156 48780 72208
rect 48832 72196 48838 72208
rect 48832 72168 59860 72196
rect 48832 72156 48838 72168
rect 31297 72131 31355 72137
rect 31297 72128 31309 72131
rect 30852 72100 31309 72128
rect 9585 72091 9643 72097
rect 31297 72097 31309 72100
rect 31343 72097 31355 72131
rect 31297 72091 31355 72097
rect 55033 72131 55091 72137
rect 55033 72097 55045 72131
rect 55079 72097 55091 72131
rect 55033 72091 55091 72097
rect 55217 72131 55275 72137
rect 55217 72097 55229 72131
rect 55263 72097 55275 72131
rect 55217 72091 55275 72097
rect 30834 72020 30840 72072
rect 30892 72060 30898 72072
rect 31021 72063 31079 72069
rect 31021 72060 31033 72063
rect 30892 72032 31033 72060
rect 30892 72020 30898 72032
rect 31021 72029 31033 72032
rect 31067 72029 31079 72063
rect 31021 72023 31079 72029
rect 23198 71952 23204 72004
rect 23256 71992 23262 72004
rect 23256 71964 27936 71992
rect 23256 71952 23262 71964
rect 9674 71924 9680 71936
rect 9635 71896 9680 71924
rect 9674 71884 9680 71896
rect 9732 71884 9738 71936
rect 25133 71927 25191 71933
rect 25133 71893 25145 71927
rect 25179 71924 25191 71927
rect 25314 71924 25320 71936
rect 25179 71896 25320 71924
rect 25179 71893 25191 71896
rect 25133 71887 25191 71893
rect 25314 71884 25320 71896
rect 25372 71924 25378 71936
rect 25409 71927 25467 71933
rect 25409 71924 25421 71927
rect 25372 71896 25421 71924
rect 25372 71884 25378 71896
rect 25409 71893 25421 71896
rect 25455 71893 25467 71927
rect 27908 71924 27936 71964
rect 32401 71927 32459 71933
rect 32401 71924 32413 71927
rect 27908 71896 32413 71924
rect 25409 71887 25467 71893
rect 32401 71893 32413 71896
rect 32447 71893 32459 71927
rect 54846 71924 54852 71936
rect 54807 71896 54852 71924
rect 32401 71887 32459 71893
rect 54846 71884 54852 71896
rect 54904 71884 54910 71936
rect 55048 71924 55076 72091
rect 55232 72004 55260 72091
rect 55306 72088 55312 72140
rect 55364 72128 55370 72140
rect 59832 72137 59860 72168
rect 59998 72156 60004 72208
rect 60056 72196 60062 72208
rect 60185 72199 60243 72205
rect 60185 72196 60197 72199
rect 60056 72168 60197 72196
rect 60056 72156 60062 72168
rect 60185 72165 60197 72168
rect 60231 72165 60243 72199
rect 60185 72159 60243 72165
rect 59817 72131 59875 72137
rect 55364 72100 55409 72128
rect 55364 72088 55370 72100
rect 59817 72097 59829 72131
rect 59863 72097 59875 72131
rect 59817 72091 59875 72097
rect 59906 72088 59912 72140
rect 59964 72128 59970 72140
rect 60090 72128 60096 72140
rect 59964 72100 60009 72128
rect 60051 72100 60096 72128
rect 59964 72088 59970 72100
rect 60090 72088 60096 72100
rect 60148 72088 60154 72140
rect 60292 72137 60320 72236
rect 64846 72236 79968 72264
rect 60282 72131 60340 72137
rect 60282 72097 60294 72131
rect 60328 72097 60340 72131
rect 60282 72091 60340 72097
rect 60108 72060 60136 72088
rect 64846 72060 64874 72236
rect 79962 72224 79968 72236
rect 80020 72224 80026 72276
rect 78674 72088 78680 72140
rect 78732 72128 78738 72140
rect 79137 72131 79195 72137
rect 79137 72128 79149 72131
rect 78732 72100 79149 72128
rect 78732 72088 78738 72100
rect 79137 72097 79149 72100
rect 79183 72097 79195 72131
rect 79137 72091 79195 72097
rect 78858 72060 78864 72072
rect 60108 72032 64874 72060
rect 78819 72032 78864 72060
rect 78858 72020 78864 72032
rect 78916 72020 78922 72072
rect 55214 71952 55220 72004
rect 55272 71952 55278 72004
rect 59538 71992 59544 72004
rect 55416 71964 59544 71992
rect 55416 71924 55444 71964
rect 59538 71952 59544 71964
rect 59596 71992 59602 72004
rect 63218 71992 63224 72004
rect 59596 71964 63224 71992
rect 59596 71952 59602 71964
rect 63218 71952 63224 71964
rect 63276 71952 63282 72004
rect 93670 71992 93676 72004
rect 84166 71964 93676 71992
rect 55048 71896 55444 71924
rect 60461 71927 60519 71933
rect 60461 71893 60473 71927
rect 60507 71924 60519 71927
rect 78582 71924 78588 71936
rect 60507 71896 78588 71924
rect 60507 71893 60519 71896
rect 60461 71887 60519 71893
rect 78582 71884 78588 71896
rect 78640 71884 78646 71936
rect 78674 71884 78680 71936
rect 78732 71924 78738 71936
rect 80238 71924 80244 71936
rect 78732 71896 78777 71924
rect 80199 71896 80244 71924
rect 78732 71884 78738 71896
rect 80238 71884 80244 71896
rect 80296 71924 80302 71936
rect 84166 71924 84194 71964
rect 93670 71952 93676 71964
rect 93728 71952 93734 72004
rect 89254 71924 89260 71936
rect 80296 71896 84194 71924
rect 89215 71896 89260 71924
rect 80296 71884 80302 71896
rect 89254 71884 89260 71896
rect 89312 71924 89318 71936
rect 89441 71927 89499 71933
rect 89441 71924 89453 71927
rect 89312 71896 89453 71924
rect 89312 71884 89318 71896
rect 89441 71893 89453 71896
rect 89487 71893 89499 71927
rect 89441 71887 89499 71893
rect 1104 71834 98808 71856
rect 1104 71782 4246 71834
rect 4298 71782 4310 71834
rect 4362 71782 4374 71834
rect 4426 71782 4438 71834
rect 4490 71782 34966 71834
rect 35018 71782 35030 71834
rect 35082 71782 35094 71834
rect 35146 71782 35158 71834
rect 35210 71782 65686 71834
rect 65738 71782 65750 71834
rect 65802 71782 65814 71834
rect 65866 71782 65878 71834
rect 65930 71782 96406 71834
rect 96458 71782 96470 71834
rect 96522 71782 96534 71834
rect 96586 71782 96598 71834
rect 96650 71782 98808 71834
rect 1104 71760 98808 71782
rect 71222 71652 71228 71664
rect 71183 71624 71228 71652
rect 71222 71612 71228 71624
rect 71280 71612 71286 71664
rect 65889 71587 65947 71593
rect 65889 71553 65901 71587
rect 65935 71584 65947 71587
rect 66162 71584 66168 71596
rect 65935 71556 66168 71584
rect 65935 71553 65947 71556
rect 65889 71547 65947 71553
rect 66162 71544 66168 71556
rect 66220 71544 66226 71596
rect 85666 71584 85672 71596
rect 70688 71556 85672 71584
rect 70688 71528 70716 71556
rect 85666 71544 85672 71556
rect 85724 71544 85730 71596
rect 22465 71519 22523 71525
rect 22465 71485 22477 71519
rect 22511 71516 22523 71519
rect 22741 71519 22799 71525
rect 22741 71516 22753 71519
rect 22511 71488 22753 71516
rect 22511 71485 22523 71488
rect 22465 71479 22523 71485
rect 22741 71485 22753 71488
rect 22787 71516 22799 71519
rect 27154 71516 27160 71528
rect 22787 71488 27160 71516
rect 22787 71485 22799 71488
rect 22741 71479 22799 71485
rect 27154 71476 27160 71488
rect 27212 71476 27218 71528
rect 54297 71519 54355 71525
rect 54297 71485 54309 71519
rect 54343 71485 54355 71519
rect 54297 71479 54355 71485
rect 65337 71519 65395 71525
rect 65337 71485 65349 71519
rect 65383 71516 65395 71519
rect 65426 71516 65432 71528
rect 65383 71488 65432 71516
rect 65383 71485 65395 71488
rect 65337 71479 65395 71485
rect 54021 71451 54079 71457
rect 54021 71417 54033 71451
rect 54067 71448 54079 71451
rect 54312 71448 54340 71479
rect 65426 71476 65432 71488
rect 65484 71476 65490 71528
rect 66533 71519 66591 71525
rect 66533 71485 66545 71519
rect 66579 71516 66591 71519
rect 66622 71516 66628 71528
rect 66579 71488 66628 71516
rect 66579 71485 66591 71488
rect 66533 71479 66591 71485
rect 66622 71476 66628 71488
rect 66680 71476 66686 71528
rect 70670 71516 70676 71528
rect 70631 71488 70676 71516
rect 70670 71476 70676 71488
rect 70728 71476 70734 71528
rect 70854 71516 70860 71528
rect 70815 71488 70860 71516
rect 70854 71476 70860 71488
rect 70912 71476 70918 71528
rect 71130 71525 71136 71528
rect 71093 71519 71136 71525
rect 71093 71485 71105 71519
rect 71093 71479 71136 71485
rect 71130 71476 71136 71479
rect 71188 71476 71194 71528
rect 70118 71448 70124 71460
rect 54067 71420 54340 71448
rect 54067 71417 54079 71420
rect 54021 71411 54079 71417
rect 24026 71340 24032 71392
rect 24084 71380 24090 71392
rect 26970 71380 26976 71392
rect 24084 71352 26976 71380
rect 24084 71340 24090 71352
rect 26970 71340 26976 71352
rect 27028 71340 27034 71392
rect 54312 71380 54340 71420
rect 64846 71420 70124 71448
rect 64846 71380 64874 71420
rect 70118 71408 70124 71420
rect 70176 71408 70182 71460
rect 70946 71448 70952 71460
rect 70907 71420 70952 71448
rect 70946 71408 70952 71420
rect 71004 71448 71010 71460
rect 75178 71448 75184 71460
rect 71004 71420 75184 71448
rect 71004 71408 71010 71420
rect 75178 71408 75184 71420
rect 75236 71408 75242 71460
rect 54312 71352 64874 71380
rect 65426 71340 65432 71392
rect 65484 71380 65490 71392
rect 66625 71383 66683 71389
rect 66625 71380 66637 71383
rect 65484 71352 66637 71380
rect 65484 71340 65490 71352
rect 66625 71349 66637 71352
rect 66671 71349 66683 71383
rect 66625 71343 66683 71349
rect 1104 71290 98808 71312
rect 1104 71238 19606 71290
rect 19658 71238 19670 71290
rect 19722 71238 19734 71290
rect 19786 71238 19798 71290
rect 19850 71238 50326 71290
rect 50378 71238 50390 71290
rect 50442 71238 50454 71290
rect 50506 71238 50518 71290
rect 50570 71238 81046 71290
rect 81098 71238 81110 71290
rect 81162 71238 81174 71290
rect 81226 71238 81238 71290
rect 81290 71238 98808 71290
rect 1104 71216 98808 71238
rect 16206 71136 16212 71188
rect 16264 71176 16270 71188
rect 26418 71176 26424 71188
rect 16264 71148 26424 71176
rect 16264 71136 16270 71148
rect 26418 71136 26424 71148
rect 26476 71136 26482 71188
rect 26970 71136 26976 71188
rect 27028 71176 27034 71188
rect 27028 71148 35894 71176
rect 27028 71136 27034 71148
rect 2130 71068 2136 71120
rect 2188 71108 2194 71120
rect 24026 71108 24032 71120
rect 2188 71080 24032 71108
rect 2188 71068 2194 71080
rect 24026 71068 24032 71080
rect 24084 71068 24090 71120
rect 26786 71108 26792 71120
rect 26747 71080 26792 71108
rect 26786 71068 26792 71080
rect 26844 71068 26850 71120
rect 35866 71108 35894 71148
rect 36354 71108 36360 71120
rect 35866 71080 36360 71108
rect 36354 71068 36360 71080
rect 36412 71068 36418 71120
rect 53282 71068 53288 71120
rect 53340 71108 53346 71120
rect 63586 71108 63592 71120
rect 53340 71080 63592 71108
rect 53340 71068 53346 71080
rect 63586 71068 63592 71080
rect 63644 71068 63650 71120
rect 26326 71000 26332 71052
rect 26384 71040 26390 71052
rect 26513 71043 26571 71049
rect 26513 71040 26525 71043
rect 26384 71012 26525 71040
rect 26384 71000 26390 71012
rect 26513 71009 26525 71012
rect 26559 71009 26571 71043
rect 26694 71040 26700 71052
rect 26655 71012 26700 71040
rect 26513 71003 26571 71009
rect 26694 71000 26700 71012
rect 26752 71000 26758 71052
rect 26886 71043 26944 71049
rect 26886 71009 26898 71043
rect 26932 71009 26944 71043
rect 26886 71003 26944 71009
rect 6886 70944 25820 70972
rect 2501 70907 2559 70913
rect 2501 70873 2513 70907
rect 2547 70904 2559 70907
rect 2777 70907 2835 70913
rect 2777 70904 2789 70907
rect 2547 70876 2789 70904
rect 2547 70873 2559 70876
rect 2501 70867 2559 70873
rect 2777 70873 2789 70876
rect 2823 70904 2835 70907
rect 6886 70904 6914 70944
rect 2823 70876 6914 70904
rect 2823 70873 2835 70876
rect 2777 70867 2835 70873
rect 25409 70839 25467 70845
rect 25409 70805 25421 70839
rect 25455 70836 25467 70839
rect 25682 70836 25688 70848
rect 25455 70808 25688 70836
rect 25455 70805 25467 70808
rect 25409 70799 25467 70805
rect 25682 70796 25688 70808
rect 25740 70796 25746 70848
rect 25792 70836 25820 70944
rect 26786 70932 26792 70984
rect 26844 70972 26850 70984
rect 26896 70972 26924 71003
rect 53374 71000 53380 71052
rect 53432 71040 53438 71052
rect 68094 71040 68100 71052
rect 53432 71012 68100 71040
rect 53432 71000 53438 71012
rect 68094 71000 68100 71012
rect 68152 71000 68158 71052
rect 26844 70944 26924 70972
rect 26844 70932 26850 70944
rect 27154 70932 27160 70984
rect 27212 70972 27218 70984
rect 95602 70972 95608 70984
rect 27212 70944 95608 70972
rect 27212 70932 27218 70944
rect 95602 70932 95608 70944
rect 95660 70932 95666 70984
rect 27062 70904 27068 70916
rect 27023 70876 27068 70904
rect 27062 70864 27068 70876
rect 27120 70864 27126 70916
rect 94774 70904 94780 70916
rect 35866 70876 94780 70904
rect 35866 70836 35894 70876
rect 94774 70864 94780 70876
rect 94832 70864 94838 70916
rect 25792 70808 35894 70836
rect 83458 70796 83464 70848
rect 83516 70836 83522 70848
rect 83553 70839 83611 70845
rect 83553 70836 83565 70839
rect 83516 70808 83565 70836
rect 83516 70796 83522 70808
rect 83553 70805 83565 70808
rect 83599 70836 83611 70839
rect 83737 70839 83795 70845
rect 83737 70836 83749 70839
rect 83599 70808 83749 70836
rect 83599 70805 83611 70808
rect 83553 70799 83611 70805
rect 83737 70805 83749 70808
rect 83783 70805 83795 70839
rect 83737 70799 83795 70805
rect 1104 70746 98808 70768
rect 1104 70694 4246 70746
rect 4298 70694 4310 70746
rect 4362 70694 4374 70746
rect 4426 70694 4438 70746
rect 4490 70694 34966 70746
rect 35018 70694 35030 70746
rect 35082 70694 35094 70746
rect 35146 70694 35158 70746
rect 35210 70694 65686 70746
rect 65738 70694 65750 70746
rect 65802 70694 65814 70746
rect 65866 70694 65878 70746
rect 65930 70694 96406 70746
rect 96458 70694 96470 70746
rect 96522 70694 96534 70746
rect 96586 70694 96598 70746
rect 96650 70694 98808 70746
rect 1104 70672 98808 70694
rect 25682 70592 25688 70644
rect 25740 70632 25746 70644
rect 70026 70632 70032 70644
rect 25740 70604 70032 70632
rect 25740 70592 25746 70604
rect 70026 70592 70032 70604
rect 70084 70592 70090 70644
rect 52733 70499 52791 70505
rect 52733 70465 52745 70499
rect 52779 70496 52791 70499
rect 53009 70499 53067 70505
rect 53009 70496 53021 70499
rect 52779 70468 53021 70496
rect 52779 70465 52791 70468
rect 52733 70459 52791 70465
rect 53009 70465 53021 70468
rect 53055 70496 53067 70499
rect 64230 70496 64236 70508
rect 53055 70468 64236 70496
rect 53055 70465 53067 70468
rect 53009 70459 53067 70465
rect 64230 70456 64236 70468
rect 64288 70456 64294 70508
rect 84562 70456 84568 70508
rect 84620 70496 84626 70508
rect 87141 70499 87199 70505
rect 87141 70496 87153 70499
rect 84620 70468 87153 70496
rect 84620 70456 84626 70468
rect 87141 70465 87153 70468
rect 87187 70465 87199 70499
rect 87141 70459 87199 70465
rect 57238 70388 57244 70440
rect 57296 70428 57302 70440
rect 59998 70428 60004 70440
rect 57296 70400 60004 70428
rect 57296 70388 57302 70400
rect 59998 70388 60004 70400
rect 60056 70388 60062 70440
rect 85206 70388 85212 70440
rect 85264 70428 85270 70440
rect 85301 70431 85359 70437
rect 85301 70428 85313 70431
rect 85264 70400 85313 70428
rect 85264 70388 85270 70400
rect 85301 70397 85313 70400
rect 85347 70428 85359 70431
rect 86865 70431 86923 70437
rect 86865 70428 86877 70431
rect 85347 70400 86877 70428
rect 85347 70397 85359 70400
rect 85301 70391 85359 70397
rect 86865 70397 86877 70400
rect 86911 70397 86923 70431
rect 86865 70391 86923 70397
rect 55214 70320 55220 70372
rect 55272 70360 55278 70372
rect 77294 70360 77300 70372
rect 55272 70332 77300 70360
rect 55272 70320 55278 70332
rect 77294 70320 77300 70332
rect 77352 70320 77358 70372
rect 85574 70292 85580 70304
rect 85535 70264 85580 70292
rect 85574 70252 85580 70264
rect 85632 70252 85638 70304
rect 1104 70202 98808 70224
rect 1104 70150 19606 70202
rect 19658 70150 19670 70202
rect 19722 70150 19734 70202
rect 19786 70150 19798 70202
rect 19850 70150 50326 70202
rect 50378 70150 50390 70202
rect 50442 70150 50454 70202
rect 50506 70150 50518 70202
rect 50570 70150 81046 70202
rect 81098 70150 81110 70202
rect 81162 70150 81174 70202
rect 81226 70150 81238 70202
rect 81290 70150 98808 70202
rect 1104 70128 98808 70150
rect 15749 69955 15807 69961
rect 15749 69921 15761 69955
rect 15795 69952 15807 69955
rect 43530 69952 43536 69964
rect 15795 69924 43536 69952
rect 15795 69921 15807 69924
rect 15749 69915 15807 69921
rect 43530 69912 43536 69924
rect 43588 69912 43594 69964
rect 50154 69912 50160 69964
rect 50212 69952 50218 69964
rect 78674 69952 78680 69964
rect 50212 69924 78680 69952
rect 50212 69912 50218 69924
rect 78674 69912 78680 69924
rect 78732 69912 78738 69964
rect 11330 69844 11336 69896
rect 11388 69884 11394 69896
rect 55214 69884 55220 69896
rect 11388 69856 55220 69884
rect 11388 69844 11394 69856
rect 55214 69844 55220 69856
rect 55272 69844 55278 69896
rect 61562 69844 61568 69896
rect 61620 69884 61626 69896
rect 93026 69884 93032 69896
rect 61620 69856 93032 69884
rect 61620 69844 61626 69856
rect 93026 69844 93032 69856
rect 93084 69844 93090 69896
rect 15930 69816 15936 69828
rect 15891 69788 15936 69816
rect 15930 69776 15936 69788
rect 15988 69776 15994 69828
rect 37918 69776 37924 69828
rect 37976 69816 37982 69828
rect 89254 69816 89260 69828
rect 37976 69788 89260 69816
rect 37976 69776 37982 69788
rect 89254 69776 89260 69788
rect 89312 69776 89318 69828
rect 23658 69708 23664 69760
rect 23716 69748 23722 69760
rect 77202 69748 77208 69760
rect 23716 69720 77208 69748
rect 23716 69708 23722 69720
rect 77202 69708 77208 69720
rect 77260 69708 77266 69760
rect 1104 69658 98808 69680
rect 1104 69606 4246 69658
rect 4298 69606 4310 69658
rect 4362 69606 4374 69658
rect 4426 69606 4438 69658
rect 4490 69606 34966 69658
rect 35018 69606 35030 69658
rect 35082 69606 35094 69658
rect 35146 69606 35158 69658
rect 35210 69606 65686 69658
rect 65738 69606 65750 69658
rect 65802 69606 65814 69658
rect 65866 69606 65878 69658
rect 65930 69606 96406 69658
rect 96458 69606 96470 69658
rect 96522 69606 96534 69658
rect 96586 69606 96598 69658
rect 96650 69606 98808 69658
rect 1104 69584 98808 69606
rect 2409 69479 2467 69485
rect 2409 69445 2421 69479
rect 2455 69476 2467 69479
rect 5074 69476 5080 69488
rect 2455 69448 5080 69476
rect 2455 69445 2467 69448
rect 2409 69439 2467 69445
rect 5074 69436 5080 69448
rect 5132 69436 5138 69488
rect 61289 69411 61347 69417
rect 61289 69408 61301 69411
rect 41386 69380 61301 69408
rect 26786 69300 26792 69352
rect 26844 69340 26850 69352
rect 28258 69340 28264 69352
rect 26844 69312 28264 69340
rect 26844 69300 26850 69312
rect 28258 69300 28264 69312
rect 28316 69300 28322 69352
rect 33870 69300 33876 69352
rect 33928 69340 33934 69352
rect 41386 69340 41414 69380
rect 61289 69377 61301 69380
rect 61335 69408 61347 69411
rect 61473 69411 61531 69417
rect 61473 69408 61485 69411
rect 61335 69380 61485 69408
rect 61335 69377 61347 69380
rect 61289 69371 61347 69377
rect 61473 69377 61485 69380
rect 61519 69377 61531 69411
rect 61473 69371 61531 69377
rect 33928 69312 41414 69340
rect 52549 69343 52607 69349
rect 33928 69300 33934 69312
rect 52549 69309 52561 69343
rect 52595 69309 52607 69343
rect 52549 69303 52607 69309
rect 88705 69343 88763 69349
rect 88705 69309 88717 69343
rect 88751 69309 88763 69343
rect 88705 69303 88763 69309
rect 2041 69275 2099 69281
rect 2041 69241 2053 69275
rect 2087 69272 2099 69275
rect 2225 69275 2283 69281
rect 2225 69272 2237 69275
rect 2087 69244 2237 69272
rect 2087 69241 2099 69244
rect 2041 69235 2099 69241
rect 2225 69241 2237 69244
rect 2271 69272 2283 69275
rect 5258 69272 5264 69284
rect 2271 69244 5264 69272
rect 2271 69241 2283 69244
rect 2225 69235 2283 69241
rect 5258 69232 5264 69244
rect 5316 69232 5322 69284
rect 47578 69164 47584 69216
rect 47636 69204 47642 69216
rect 52457 69207 52515 69213
rect 52457 69204 52469 69207
rect 47636 69176 52469 69204
rect 47636 69164 47642 69176
rect 52457 69173 52469 69176
rect 52503 69204 52515 69207
rect 52564 69204 52592 69303
rect 88720 69216 88748 69303
rect 52503 69176 52592 69204
rect 88613 69207 88671 69213
rect 52503 69173 52515 69176
rect 52457 69167 52515 69173
rect 88613 69173 88625 69207
rect 88659 69204 88671 69207
rect 88702 69204 88708 69216
rect 88659 69176 88708 69204
rect 88659 69173 88671 69176
rect 88613 69167 88671 69173
rect 88702 69164 88708 69176
rect 88760 69164 88766 69216
rect 1104 69114 98808 69136
rect 1104 69062 19606 69114
rect 19658 69062 19670 69114
rect 19722 69062 19734 69114
rect 19786 69062 19798 69114
rect 19850 69062 50326 69114
rect 50378 69062 50390 69114
rect 50442 69062 50454 69114
rect 50506 69062 50518 69114
rect 50570 69062 81046 69114
rect 81098 69062 81110 69114
rect 81162 69062 81174 69114
rect 81226 69062 81238 69114
rect 81290 69062 98808 69114
rect 1104 69040 98808 69062
rect 5350 68960 5356 69012
rect 5408 69000 5414 69012
rect 77481 69003 77539 69009
rect 77481 69000 77493 69003
rect 5408 68972 77493 69000
rect 5408 68960 5414 68972
rect 77481 68969 77493 68972
rect 77527 69000 77539 69003
rect 77527 68972 78168 69000
rect 77527 68969 77539 68972
rect 77481 68963 77539 68969
rect 70366 68904 78076 68932
rect 15930 68864 15936 68876
rect 15891 68836 15936 68864
rect 15930 68824 15936 68836
rect 15988 68824 15994 68876
rect 61378 68824 61384 68876
rect 61436 68864 61442 68876
rect 70366 68864 70394 68904
rect 78048 68873 78076 68904
rect 78140 68873 78168 68972
rect 78306 68960 78312 69012
rect 78364 69000 78370 69012
rect 78364 68972 85804 69000
rect 78364 68960 78370 68972
rect 85776 68932 85804 68972
rect 85850 68960 85856 69012
rect 85908 69000 85914 69012
rect 85945 69003 86003 69009
rect 85945 69000 85957 69003
rect 85908 68972 85957 69000
rect 85908 68960 85914 68972
rect 85945 68969 85957 68972
rect 85991 68969 86003 69003
rect 92382 69000 92388 69012
rect 85945 68963 86003 68969
rect 86052 68972 92388 69000
rect 86052 68932 86080 68972
rect 92382 68960 92388 68972
rect 92440 68960 92446 69012
rect 85776 68904 86080 68932
rect 61436 68836 70394 68864
rect 77665 68867 77723 68873
rect 61436 68824 61442 68836
rect 77665 68833 77677 68867
rect 77711 68833 77723 68867
rect 77665 68827 77723 68833
rect 78033 68867 78091 68873
rect 78033 68833 78045 68867
rect 78079 68833 78091 68867
rect 78033 68827 78091 68833
rect 78125 68867 78183 68873
rect 78125 68833 78137 68867
rect 78171 68833 78183 68867
rect 78125 68827 78183 68833
rect 16482 68796 16488 68808
rect 16443 68768 16488 68796
rect 16482 68756 16488 68768
rect 16540 68756 16546 68808
rect 61930 68796 61936 68808
rect 61891 68768 61936 68796
rect 61930 68756 61936 68768
rect 61988 68756 61994 68808
rect 62209 68799 62267 68805
rect 62209 68765 62221 68799
rect 62255 68796 62267 68799
rect 62390 68796 62396 68808
rect 62255 68768 62396 68796
rect 62255 68765 62267 68768
rect 62209 68759 62267 68765
rect 62390 68756 62396 68768
rect 62448 68756 62454 68808
rect 77680 68728 77708 68827
rect 78214 68824 78220 68876
rect 78272 68864 78278 68876
rect 78401 68867 78459 68873
rect 78401 68864 78413 68867
rect 78272 68836 78413 68864
rect 78272 68824 78278 68836
rect 78401 68833 78413 68836
rect 78447 68864 78459 68867
rect 78490 68864 78496 68876
rect 78447 68836 78496 68864
rect 78447 68833 78459 68836
rect 78401 68827 78459 68833
rect 78490 68824 78496 68836
rect 78548 68824 78554 68876
rect 83550 68824 83556 68876
rect 83608 68864 83614 68876
rect 90361 68867 90419 68873
rect 90361 68864 90373 68867
rect 83608 68836 90373 68864
rect 83608 68824 83614 68836
rect 90361 68833 90373 68836
rect 90407 68833 90419 68867
rect 90361 68827 90419 68833
rect 92017 68867 92075 68873
rect 92017 68833 92029 68867
rect 92063 68864 92075 68867
rect 92382 68864 92388 68876
rect 92063 68836 92388 68864
rect 92063 68833 92075 68836
rect 92017 68827 92075 68833
rect 92382 68824 92388 68836
rect 92440 68824 92446 68876
rect 78306 68796 78312 68808
rect 78267 68768 78312 68796
rect 78306 68756 78312 68768
rect 78364 68756 78370 68808
rect 80790 68796 80796 68808
rect 78600 68768 80796 68796
rect 78600 68728 78628 68768
rect 80790 68756 80796 68768
rect 80848 68756 80854 68808
rect 84562 68796 84568 68808
rect 84523 68768 84568 68796
rect 84562 68756 84568 68768
rect 84620 68756 84626 68808
rect 84838 68796 84844 68808
rect 84799 68768 84844 68796
rect 84838 68756 84844 68768
rect 84896 68756 84902 68808
rect 91741 68799 91799 68805
rect 91741 68796 91753 68799
rect 90192 68768 91753 68796
rect 78766 68728 78772 68740
rect 77680 68700 78628 68728
rect 78727 68700 78772 68728
rect 78766 68688 78772 68700
rect 78824 68688 78830 68740
rect 90192 68672 90220 68768
rect 91741 68765 91753 68768
rect 91787 68765 91799 68799
rect 91741 68759 91799 68765
rect 63497 68663 63555 68669
rect 63497 68629 63509 68663
rect 63543 68660 63555 68663
rect 63678 68660 63684 68672
rect 63543 68632 63684 68660
rect 63543 68629 63555 68632
rect 63497 68623 63555 68629
rect 63678 68620 63684 68632
rect 63736 68620 63742 68672
rect 90174 68660 90180 68672
rect 90135 68632 90180 68660
rect 90174 68620 90180 68632
rect 90232 68620 90238 68672
rect 1104 68570 98808 68592
rect 1104 68518 4246 68570
rect 4298 68518 4310 68570
rect 4362 68518 4374 68570
rect 4426 68518 4438 68570
rect 4490 68518 34966 68570
rect 35018 68518 35030 68570
rect 35082 68518 35094 68570
rect 35146 68518 35158 68570
rect 35210 68518 65686 68570
rect 65738 68518 65750 68570
rect 65802 68518 65814 68570
rect 65866 68518 65878 68570
rect 65930 68518 96406 68570
rect 96458 68518 96470 68570
rect 96522 68518 96534 68570
rect 96586 68518 96598 68570
rect 96650 68518 98808 68570
rect 1104 68496 98808 68518
rect 46198 68416 46204 68468
rect 46256 68456 46262 68468
rect 46256 68428 46705 68456
rect 46256 68416 46262 68428
rect 45554 68348 45560 68400
rect 45612 68388 45618 68400
rect 46677 68388 46705 68428
rect 91186 68416 91192 68468
rect 91244 68456 91250 68468
rect 92569 68459 92627 68465
rect 92569 68456 92581 68459
rect 91244 68428 92581 68456
rect 91244 68416 91250 68428
rect 92569 68425 92581 68428
rect 92615 68425 92627 68459
rect 92569 68419 92627 68425
rect 90082 68388 90088 68400
rect 45612 68360 46612 68388
rect 45612 68348 45618 68360
rect 10042 68320 10048 68332
rect 10003 68292 10048 68320
rect 10042 68280 10048 68292
rect 10100 68280 10106 68332
rect 15930 68320 15936 68332
rect 10520 68292 15936 68320
rect 6733 68255 6791 68261
rect 6733 68221 6745 68255
rect 6779 68252 6791 68255
rect 7006 68252 7012 68264
rect 6779 68224 7012 68252
rect 6779 68221 6791 68224
rect 6733 68215 6791 68221
rect 7006 68212 7012 68224
rect 7064 68212 7070 68264
rect 9766 68252 9772 68264
rect 9727 68224 9772 68252
rect 9766 68212 9772 68224
rect 9824 68212 9830 68264
rect 10520 68261 10548 68292
rect 15930 68280 15936 68292
rect 15988 68280 15994 68332
rect 31386 68280 31392 68332
rect 31444 68320 31450 68332
rect 31444 68292 46336 68320
rect 31444 68280 31450 68292
rect 10137 68255 10195 68261
rect 10137 68221 10149 68255
rect 10183 68221 10195 68255
rect 10137 68215 10195 68221
rect 10505 68255 10563 68261
rect 10505 68221 10517 68255
rect 10551 68221 10563 68255
rect 10686 68252 10692 68264
rect 10647 68224 10692 68252
rect 10505 68215 10563 68221
rect 10152 68184 10180 68215
rect 10686 68212 10692 68224
rect 10744 68212 10750 68264
rect 26878 68212 26884 68264
rect 26936 68252 26942 68264
rect 46308 68261 46336 68292
rect 46382 68280 46388 68332
rect 46440 68320 46446 68332
rect 46584 68329 46612 68360
rect 46677 68360 90088 68388
rect 46477 68323 46535 68329
rect 46477 68320 46489 68323
rect 46440 68292 46489 68320
rect 46440 68280 46446 68292
rect 46477 68289 46489 68292
rect 46523 68289 46535 68323
rect 46477 68283 46535 68289
rect 46569 68323 46627 68329
rect 46569 68289 46581 68323
rect 46615 68289 46627 68323
rect 46569 68283 46627 68289
rect 46677 68261 46705 68360
rect 90082 68348 90088 68360
rect 90140 68348 90146 68400
rect 91830 68348 91836 68400
rect 91888 68388 91894 68400
rect 91888 68360 92332 68388
rect 91888 68348 91894 68360
rect 80698 68280 80704 68332
rect 80756 68320 80762 68332
rect 91922 68320 91928 68332
rect 80756 68292 91928 68320
rect 80756 68280 80762 68292
rect 91922 68280 91928 68292
rect 91980 68280 91986 68332
rect 92106 68280 92112 68332
rect 92164 68320 92170 68332
rect 92164 68292 92244 68320
rect 92164 68280 92170 68292
rect 46109 68255 46167 68261
rect 46109 68252 46121 68255
rect 26936 68224 46121 68252
rect 26936 68212 26942 68224
rect 46109 68221 46121 68224
rect 46155 68221 46167 68255
rect 46109 68215 46167 68221
rect 46293 68255 46351 68261
rect 46293 68221 46305 68255
rect 46339 68221 46351 68255
rect 46293 68215 46351 68221
rect 46662 68255 46720 68261
rect 46662 68221 46674 68255
rect 46708 68221 46720 68255
rect 46842 68252 46848 68264
rect 46803 68224 46848 68252
rect 46662 68215 46720 68221
rect 46842 68212 46848 68224
rect 46900 68212 46906 68264
rect 91738 68212 91744 68264
rect 91796 68252 91802 68264
rect 92216 68261 92244 68292
rect 92017 68255 92075 68261
rect 92017 68252 92029 68255
rect 91796 68224 92029 68252
rect 91796 68212 91802 68224
rect 92017 68221 92029 68224
rect 92063 68221 92075 68255
rect 92017 68215 92075 68221
rect 92201 68255 92259 68261
rect 92201 68221 92213 68255
rect 92247 68221 92259 68255
rect 92304 68252 92332 68360
rect 92385 68255 92443 68261
rect 92385 68252 92397 68255
rect 92304 68224 92397 68252
rect 92201 68215 92259 68221
rect 92385 68221 92397 68224
rect 92431 68221 92443 68255
rect 92385 68215 92443 68221
rect 16114 68184 16120 68196
rect 10152 68156 16120 68184
rect 16114 68144 16120 68156
rect 16172 68144 16178 68196
rect 38626 68156 46336 68184
rect 10965 68119 11023 68125
rect 10965 68085 10977 68119
rect 11011 68116 11023 68119
rect 38626 68116 38654 68156
rect 11011 68088 38654 68116
rect 11011 68085 11023 68088
rect 10965 68079 11023 68085
rect 39758 68076 39764 68128
rect 39816 68116 39822 68128
rect 45925 68119 45983 68125
rect 45925 68116 45937 68119
rect 39816 68088 45937 68116
rect 39816 68076 39822 68088
rect 45925 68085 45937 68088
rect 45971 68116 45983 68119
rect 46198 68116 46204 68128
rect 45971 68088 46204 68116
rect 45971 68085 45983 68088
rect 45925 68079 45983 68085
rect 46198 68076 46204 68088
rect 46256 68076 46262 68128
rect 46308 68116 46336 68156
rect 75454 68144 75460 68196
rect 75512 68184 75518 68196
rect 92293 68187 92351 68193
rect 75512 68156 92152 68184
rect 75512 68144 75518 68156
rect 84838 68116 84844 68128
rect 46308 68088 84844 68116
rect 84838 68076 84844 68088
rect 84896 68076 84902 68128
rect 92124 68116 92152 68156
rect 92293 68153 92305 68187
rect 92339 68153 92351 68187
rect 92293 68147 92351 68153
rect 92304 68116 92332 68147
rect 92124 68088 92332 68116
rect 1104 68026 98808 68048
rect 1104 67974 19606 68026
rect 19658 67974 19670 68026
rect 19722 67974 19734 68026
rect 19786 67974 19798 68026
rect 19850 67974 50326 68026
rect 50378 67974 50390 68026
rect 50442 67974 50454 68026
rect 50506 67974 50518 68026
rect 50570 67974 81046 68026
rect 81098 67974 81110 68026
rect 81162 67974 81174 68026
rect 81226 67974 81238 68026
rect 81290 67974 98808 68026
rect 1104 67952 98808 67974
rect 16114 67776 16120 67788
rect 16075 67748 16120 67776
rect 16114 67736 16120 67748
rect 16172 67736 16178 67788
rect 43993 67779 44051 67785
rect 43993 67776 44005 67779
rect 16546 67748 44005 67776
rect 4706 67668 4712 67720
rect 4764 67708 4770 67720
rect 5166 67708 5172 67720
rect 4764 67680 5172 67708
rect 4764 67668 4770 67680
rect 5166 67668 5172 67680
rect 5224 67708 5230 67720
rect 16546 67708 16574 67748
rect 43993 67745 44005 67748
rect 44039 67745 44051 67779
rect 43993 67739 44051 67745
rect 16942 67708 16948 67720
rect 5224 67680 16574 67708
rect 16903 67680 16948 67708
rect 5224 67668 5230 67680
rect 16942 67668 16948 67680
rect 17000 67668 17006 67720
rect 44821 67711 44879 67717
rect 44821 67677 44833 67711
rect 44867 67708 44879 67711
rect 44867 67680 60734 67708
rect 44867 67677 44879 67680
rect 44821 67671 44879 67677
rect 60706 67640 60734 67680
rect 73522 67640 73528 67652
rect 60706 67612 73528 67640
rect 73522 67600 73528 67612
rect 73580 67640 73586 67652
rect 74074 67640 74080 67652
rect 73580 67612 74080 67640
rect 73580 67600 73586 67612
rect 74074 67600 74080 67612
rect 74132 67600 74138 67652
rect 90637 67643 90695 67649
rect 90637 67609 90649 67643
rect 90683 67640 90695 67643
rect 90910 67640 90916 67652
rect 90683 67612 90916 67640
rect 90683 67609 90695 67612
rect 90637 67603 90695 67609
rect 90910 67600 90916 67612
rect 90968 67600 90974 67652
rect 4982 67532 4988 67584
rect 5040 67572 5046 67584
rect 5258 67572 5264 67584
rect 5040 67544 5264 67572
rect 5040 67532 5046 67544
rect 5258 67532 5264 67544
rect 5316 67572 5322 67584
rect 23474 67572 23480 67584
rect 5316 67544 23480 67572
rect 5316 67532 5322 67544
rect 23474 67532 23480 67544
rect 23532 67572 23538 67584
rect 23750 67572 23756 67584
rect 23532 67544 23756 67572
rect 23532 67532 23538 67544
rect 23750 67532 23756 67544
rect 23808 67532 23814 67584
rect 29270 67532 29276 67584
rect 29328 67572 29334 67584
rect 29914 67572 29920 67584
rect 29328 67544 29920 67572
rect 29328 67532 29334 67544
rect 29914 67532 29920 67544
rect 29972 67532 29978 67584
rect 1104 67482 98808 67504
rect 1104 67430 4246 67482
rect 4298 67430 4310 67482
rect 4362 67430 4374 67482
rect 4426 67430 4438 67482
rect 4490 67430 34966 67482
rect 35018 67430 35030 67482
rect 35082 67430 35094 67482
rect 35146 67430 35158 67482
rect 35210 67430 65686 67482
rect 65738 67430 65750 67482
rect 65802 67430 65814 67482
rect 65866 67430 65878 67482
rect 65930 67430 96406 67482
rect 96458 67430 96470 67482
rect 96522 67430 96534 67482
rect 96586 67430 96598 67482
rect 96650 67430 98808 67482
rect 1104 67408 98808 67430
rect 3605 67371 3663 67377
rect 3605 67337 3617 67371
rect 3651 67368 3663 67371
rect 4062 67368 4068 67380
rect 3651 67340 4068 67368
rect 3651 67337 3663 67340
rect 3605 67331 3663 67337
rect 4062 67328 4068 67340
rect 4120 67368 4126 67380
rect 73890 67368 73896 67380
rect 4120 67340 73896 67368
rect 4120 67328 4126 67340
rect 73890 67328 73896 67340
rect 73948 67328 73954 67380
rect 4246 67260 4252 67312
rect 4304 67300 4310 67312
rect 4706 67300 4712 67312
rect 4304 67272 4712 67300
rect 4304 67260 4310 67272
rect 4706 67260 4712 67272
rect 4764 67260 4770 67312
rect 16546 67272 26234 67300
rect 4154 67241 4160 67244
rect 4148 67195 4160 67241
rect 4212 67232 4218 67244
rect 4212 67204 4248 67232
rect 4154 67192 4160 67195
rect 4212 67192 4218 67204
rect 5166 67192 5172 67244
rect 5224 67232 5230 67244
rect 13630 67232 13636 67244
rect 5224 67204 13636 67232
rect 5224 67192 5230 67204
rect 13630 67192 13636 67204
rect 13688 67192 13694 67244
rect 3881 67167 3939 67173
rect 3881 67133 3893 67167
rect 3927 67164 3939 67167
rect 3970 67164 3976 67176
rect 3927 67136 3976 67164
rect 3927 67133 3939 67136
rect 3881 67127 3939 67133
rect 3970 67124 3976 67136
rect 4028 67124 4034 67176
rect 4062 67124 4068 67176
rect 4120 67164 4126 67176
rect 4430 67173 4436 67176
rect 4249 67167 4307 67173
rect 4120 67136 4165 67164
rect 4120 67124 4126 67136
rect 4249 67133 4261 67167
rect 4295 67133 4307 67167
rect 4249 67127 4307 67133
rect 4429 67127 4436 67173
rect 4488 67164 4494 67176
rect 4522 67164 4528 67176
rect 4488 67136 4528 67164
rect 3697 67099 3755 67105
rect 3697 67065 3709 67099
rect 3743 67096 3755 67099
rect 4154 67096 4160 67108
rect 3743 67068 4160 67096
rect 3743 67065 3755 67068
rect 3697 67059 3755 67065
rect 4154 67056 4160 67068
rect 4212 67056 4218 67108
rect 4276 67028 4304 67127
rect 4430 67124 4436 67127
rect 4488 67124 4494 67136
rect 4522 67124 4528 67136
rect 4580 67164 4586 67176
rect 4617 67167 4675 67173
rect 4617 67164 4629 67167
rect 4580 67136 4629 67164
rect 4580 67124 4586 67136
rect 4617 67133 4629 67136
rect 4663 67164 4675 67167
rect 16546 67164 16574 67272
rect 19426 67192 19432 67244
rect 19484 67232 19490 67244
rect 19705 67235 19763 67241
rect 19705 67232 19717 67235
rect 19484 67204 19717 67232
rect 19484 67192 19490 67204
rect 19705 67201 19717 67204
rect 19751 67201 19763 67235
rect 20622 67232 20628 67244
rect 20583 67204 20628 67232
rect 19705 67195 19763 67201
rect 20622 67192 20628 67204
rect 20680 67192 20686 67244
rect 26206 67232 26234 67272
rect 30834 67260 30840 67312
rect 30892 67300 30898 67312
rect 33781 67303 33839 67309
rect 33781 67300 33793 67303
rect 30892 67272 33793 67300
rect 30892 67260 30898 67272
rect 33781 67269 33793 67272
rect 33827 67300 33839 67303
rect 33962 67300 33968 67312
rect 33827 67272 33968 67300
rect 33827 67269 33839 67272
rect 33781 67263 33839 67269
rect 33962 67260 33968 67272
rect 34020 67260 34026 67312
rect 52181 67303 52239 67309
rect 52181 67269 52193 67303
rect 52227 67300 52239 67303
rect 89162 67300 89168 67312
rect 52227 67272 89168 67300
rect 52227 67269 52239 67272
rect 52181 67263 52239 67269
rect 89162 67260 89168 67272
rect 89220 67260 89226 67312
rect 35250 67232 35256 67244
rect 26206 67204 35256 67232
rect 35250 67192 35256 67204
rect 35308 67192 35314 67244
rect 76834 67192 76840 67244
rect 76892 67232 76898 67244
rect 76892 67204 89714 67232
rect 76892 67192 76898 67204
rect 4663 67136 16574 67164
rect 19521 67167 19579 67173
rect 4663 67133 4675 67136
rect 4617 67127 4675 67133
rect 19521 67133 19533 67167
rect 19567 67133 19579 67167
rect 19521 67127 19579 67133
rect 19889 67167 19947 67173
rect 19889 67133 19901 67167
rect 19935 67133 19947 67167
rect 20254 67164 20260 67176
rect 20215 67136 20260 67164
rect 19889 67127 19947 67133
rect 4338 67056 4344 67108
rect 4396 67096 4402 67108
rect 13538 67096 13544 67108
rect 4396 67068 13544 67096
rect 4396 67056 4402 67068
rect 13538 67056 13544 67068
rect 13596 67056 13602 67108
rect 10502 67028 10508 67040
rect 4276 67000 10508 67028
rect 10502 66988 10508 67000
rect 10560 66988 10566 67040
rect 19536 67028 19564 67127
rect 19904 67096 19932 67127
rect 20254 67124 20260 67136
rect 20312 67124 20318 67176
rect 20438 67164 20444 67176
rect 20399 67136 20444 67164
rect 20438 67124 20444 67136
rect 20496 67124 20502 67176
rect 27522 67124 27528 67176
rect 27580 67164 27586 67176
rect 33965 67167 34023 67173
rect 33965 67164 33977 67167
rect 27580 67136 33977 67164
rect 27580 67124 27586 67136
rect 33965 67133 33977 67136
rect 34011 67133 34023 67167
rect 52362 67164 52368 67176
rect 52323 67136 52368 67164
rect 33965 67127 34023 67133
rect 52362 67124 52368 67136
rect 52420 67124 52426 67176
rect 63129 67167 63187 67173
rect 63129 67133 63141 67167
rect 63175 67164 63187 67167
rect 63405 67167 63463 67173
rect 63405 67164 63417 67167
rect 63175 67136 63417 67164
rect 63175 67133 63187 67136
rect 63129 67127 63187 67133
rect 63405 67133 63417 67136
rect 63451 67164 63463 67167
rect 63586 67164 63592 67176
rect 63451 67136 63592 67164
rect 63451 67133 63463 67136
rect 63405 67127 63463 67133
rect 63586 67124 63592 67136
rect 63644 67124 63650 67176
rect 72694 67164 72700 67176
rect 72655 67136 72700 67164
rect 72694 67124 72700 67136
rect 72752 67124 72758 67176
rect 86129 67167 86187 67173
rect 86129 67164 86141 67167
rect 73172 67136 86141 67164
rect 29270 67096 29276 67108
rect 19904 67068 29276 67096
rect 29270 67056 29276 67068
rect 29328 67056 29334 67108
rect 52638 67096 52644 67108
rect 52599 67068 52644 67096
rect 52638 67056 52644 67068
rect 52696 67056 52702 67108
rect 70210 67056 70216 67108
rect 70268 67096 70274 67108
rect 73172 67096 73200 67136
rect 86129 67133 86141 67136
rect 86175 67133 86187 67167
rect 89686 67164 89714 67204
rect 90729 67167 90787 67173
rect 90729 67164 90741 67167
rect 89686 67136 90741 67164
rect 86129 67127 86187 67133
rect 90729 67133 90741 67136
rect 90775 67133 90787 67167
rect 90729 67127 90787 67133
rect 70268 67068 73200 67096
rect 73249 67099 73307 67105
rect 70268 67056 70274 67068
rect 73249 67065 73261 67099
rect 73295 67096 73307 67099
rect 76190 67096 76196 67108
rect 73295 67068 76196 67096
rect 73295 67065 73307 67068
rect 73249 67059 73307 67065
rect 76190 67056 76196 67068
rect 76248 67096 76254 67108
rect 76650 67096 76656 67108
rect 76248 67068 76656 67096
rect 76248 67056 76254 67068
rect 76650 67056 76656 67068
rect 76708 67056 76714 67108
rect 86405 67099 86463 67105
rect 86405 67065 86417 67099
rect 86451 67096 86463 67099
rect 86586 67096 86592 67108
rect 86451 67068 86592 67096
rect 86451 67065 86463 67068
rect 86405 67059 86463 67065
rect 86586 67056 86592 67068
rect 86644 67056 86650 67108
rect 91005 67099 91063 67105
rect 91005 67096 91017 67099
rect 89686 67068 91017 67096
rect 20070 67028 20076 67040
rect 19536 67000 20076 67028
rect 20070 66988 20076 67000
rect 20128 66988 20134 67040
rect 52546 67028 52552 67040
rect 52507 67000 52552 67028
rect 52546 66988 52552 67000
rect 52604 66988 52610 67040
rect 56962 66988 56968 67040
rect 57020 67028 57026 67040
rect 57882 67028 57888 67040
rect 57020 67000 57888 67028
rect 57020 66988 57026 67000
rect 57882 66988 57888 67000
rect 57940 66988 57946 67040
rect 79318 66988 79324 67040
rect 79376 67028 79382 67040
rect 79594 67028 79600 67040
rect 79376 67000 79600 67028
rect 79376 66988 79382 67000
rect 79594 66988 79600 67000
rect 79652 67028 79658 67040
rect 89686 67028 89714 67068
rect 91005 67065 91017 67068
rect 91051 67065 91063 67099
rect 91005 67059 91063 67065
rect 79652 67000 89714 67028
rect 79652 66988 79658 67000
rect 1104 66938 98808 66960
rect 1104 66886 19606 66938
rect 19658 66886 19670 66938
rect 19722 66886 19734 66938
rect 19786 66886 19798 66938
rect 19850 66886 50326 66938
rect 50378 66886 50390 66938
rect 50442 66886 50454 66938
rect 50506 66886 50518 66938
rect 50570 66886 81046 66938
rect 81098 66886 81110 66938
rect 81162 66886 81174 66938
rect 81226 66886 81238 66938
rect 81290 66886 98808 66938
rect 1104 66864 98808 66886
rect 27246 66824 27252 66836
rect 20456 66796 27252 66824
rect 20456 66697 20484 66796
rect 27246 66784 27252 66796
rect 27304 66824 27310 66836
rect 27522 66824 27528 66836
rect 27304 66796 27528 66824
rect 27304 66784 27310 66796
rect 27522 66784 27528 66796
rect 27580 66784 27586 66836
rect 34146 66824 34152 66836
rect 34107 66796 34152 66824
rect 34146 66784 34152 66796
rect 34204 66784 34210 66836
rect 63586 66784 63592 66836
rect 63644 66824 63650 66836
rect 89438 66824 89444 66836
rect 63644 66796 89444 66824
rect 63644 66784 63650 66796
rect 89438 66784 89444 66796
rect 89496 66784 89502 66836
rect 20441 66691 20499 66697
rect 20441 66657 20453 66691
rect 20487 66657 20499 66691
rect 20441 66651 20499 66657
rect 23750 66648 23756 66700
rect 23808 66688 23814 66700
rect 77941 66691 77999 66697
rect 77941 66688 77953 66691
rect 23808 66660 77953 66688
rect 23808 66648 23814 66660
rect 77941 66657 77953 66660
rect 77987 66657 77999 66691
rect 77941 66651 77999 66657
rect 4249 66623 4307 66629
rect 4249 66589 4261 66623
rect 4295 66589 4307 66623
rect 4249 66583 4307 66589
rect 4525 66623 4583 66629
rect 4525 66589 4537 66623
rect 4571 66620 4583 66623
rect 6362 66620 6368 66632
rect 4571 66592 6368 66620
rect 4571 66589 4583 66592
rect 4525 66583 4583 66589
rect 4264 66484 4292 66583
rect 6362 66580 6368 66592
rect 6420 66580 6426 66632
rect 32769 66623 32827 66629
rect 32769 66620 32781 66623
rect 26206 66592 32781 66620
rect 5813 66555 5871 66561
rect 5813 66521 5825 66555
rect 5859 66552 5871 66555
rect 17678 66552 17684 66564
rect 5859 66524 17684 66552
rect 5859 66521 5871 66524
rect 5813 66515 5871 66521
rect 17678 66512 17684 66524
rect 17736 66512 17742 66564
rect 9398 66484 9404 66496
rect 4264 66456 9404 66484
rect 9398 66444 9404 66456
rect 9456 66484 9462 66496
rect 13722 66484 13728 66496
rect 9456 66456 13728 66484
rect 9456 66444 9462 66456
rect 13722 66444 13728 66456
rect 13780 66484 13786 66496
rect 20257 66487 20315 66493
rect 20257 66484 20269 66487
rect 13780 66456 20269 66484
rect 13780 66444 13786 66456
rect 20257 66453 20269 66456
rect 20303 66484 20315 66487
rect 26206 66484 26234 66592
rect 32769 66589 32781 66592
rect 32815 66589 32827 66623
rect 32769 66583 32827 66589
rect 33045 66623 33103 66629
rect 33045 66589 33057 66623
rect 33091 66620 33103 66623
rect 46934 66620 46940 66632
rect 33091 66592 46940 66620
rect 33091 66589 33103 66592
rect 33045 66583 33103 66589
rect 46934 66580 46940 66592
rect 46992 66580 46998 66632
rect 20303 66456 26234 66484
rect 20303 66453 20315 66456
rect 20257 66447 20315 66453
rect 53282 66444 53288 66496
rect 53340 66484 53346 66496
rect 64877 66487 64935 66493
rect 64877 66484 64889 66487
rect 53340 66456 64889 66484
rect 53340 66444 53346 66456
rect 64877 66453 64889 66456
rect 64923 66484 64935 66487
rect 65061 66487 65119 66493
rect 65061 66484 65073 66487
rect 64923 66456 65073 66484
rect 64923 66453 64935 66456
rect 64877 66447 64935 66453
rect 65061 66453 65073 66456
rect 65107 66453 65119 66487
rect 77938 66484 77944 66496
rect 77899 66456 77944 66484
rect 65061 66447 65119 66453
rect 77938 66444 77944 66456
rect 77996 66444 78002 66496
rect 1104 66394 98808 66416
rect 1104 66342 4246 66394
rect 4298 66342 4310 66394
rect 4362 66342 4374 66394
rect 4426 66342 4438 66394
rect 4490 66342 34966 66394
rect 35018 66342 35030 66394
rect 35082 66342 35094 66394
rect 35146 66342 35158 66394
rect 35210 66342 65686 66394
rect 65738 66342 65750 66394
rect 65802 66342 65814 66394
rect 65866 66342 65878 66394
rect 65930 66342 96406 66394
rect 96458 66342 96470 66394
rect 96522 66342 96534 66394
rect 96586 66342 96598 66394
rect 96650 66342 98808 66394
rect 1104 66320 98808 66342
rect 80149 66147 80207 66153
rect 80149 66113 80161 66147
rect 80195 66144 80207 66147
rect 91186 66144 91192 66156
rect 80195 66116 80560 66144
rect 80195 66113 80207 66116
rect 80149 66107 80207 66113
rect 80532 66088 80560 66116
rect 82740 66116 91192 66144
rect 49510 66036 49516 66088
rect 49568 66076 49574 66088
rect 49878 66076 49884 66088
rect 49568 66048 49884 66076
rect 49568 66036 49574 66048
rect 49878 66036 49884 66048
rect 49936 66036 49942 66088
rect 78858 66036 78864 66088
rect 78916 66076 78922 66088
rect 80241 66079 80299 66085
rect 80241 66076 80253 66079
rect 78916 66048 80253 66076
rect 78916 66036 78922 66048
rect 80241 66045 80253 66048
rect 80287 66045 80299 66079
rect 80514 66076 80520 66088
rect 80475 66048 80520 66076
rect 80241 66039 80299 66045
rect 80514 66036 80520 66048
rect 80572 66036 80578 66088
rect 81986 66036 81992 66088
rect 82044 66076 82050 66088
rect 82357 66079 82415 66085
rect 82357 66076 82369 66079
rect 82044 66048 82369 66076
rect 82044 66036 82050 66048
rect 82357 66045 82369 66048
rect 82403 66045 82415 66079
rect 82538 66076 82544 66088
rect 82499 66048 82544 66076
rect 82357 66039 82415 66045
rect 82538 66036 82544 66048
rect 82596 66036 82602 66088
rect 82740 66085 82768 66116
rect 91186 66104 91192 66116
rect 91244 66104 91250 66156
rect 82725 66079 82783 66085
rect 82725 66045 82737 66079
rect 82771 66045 82783 66079
rect 83090 66076 83096 66088
rect 83051 66048 83096 66076
rect 82725 66039 82783 66045
rect 83090 66036 83096 66048
rect 83148 66036 83154 66088
rect 83274 66076 83280 66088
rect 83235 66048 83280 66076
rect 83274 66036 83280 66048
rect 83332 66036 83338 66088
rect 77294 65900 77300 65952
rect 77352 65940 77358 65952
rect 81621 65943 81679 65949
rect 81621 65940 81633 65943
rect 77352 65912 81633 65940
rect 77352 65900 77358 65912
rect 81621 65909 81633 65912
rect 81667 65909 81679 65943
rect 83550 65940 83556 65952
rect 83511 65912 83556 65940
rect 81621 65903 81679 65909
rect 83550 65900 83556 65912
rect 83608 65900 83614 65952
rect 1104 65850 98808 65872
rect 1104 65798 19606 65850
rect 19658 65798 19670 65850
rect 19722 65798 19734 65850
rect 19786 65798 19798 65850
rect 19850 65798 50326 65850
rect 50378 65798 50390 65850
rect 50442 65798 50454 65850
rect 50506 65798 50518 65850
rect 50570 65798 81046 65850
rect 81098 65798 81110 65850
rect 81162 65798 81174 65850
rect 81226 65798 81238 65850
rect 81290 65798 98808 65850
rect 1104 65776 98808 65798
rect 36538 65696 36544 65748
rect 36596 65736 36602 65748
rect 83550 65736 83556 65748
rect 36596 65708 83556 65736
rect 36596 65696 36602 65708
rect 83550 65696 83556 65708
rect 83608 65696 83614 65748
rect 2314 65628 2320 65680
rect 2372 65668 2378 65680
rect 27338 65668 27344 65680
rect 2372 65640 27344 65668
rect 2372 65628 2378 65640
rect 27338 65628 27344 65640
rect 27396 65628 27402 65680
rect 38194 65628 38200 65680
rect 38252 65668 38258 65680
rect 46750 65668 46756 65680
rect 38252 65640 46756 65668
rect 38252 65628 38258 65640
rect 46750 65628 46756 65640
rect 46808 65628 46814 65680
rect 6641 65603 6699 65609
rect 6641 65569 6653 65603
rect 6687 65600 6699 65603
rect 7374 65600 7380 65612
rect 6687 65572 7380 65600
rect 6687 65569 6699 65572
rect 6641 65563 6699 65569
rect 7374 65560 7380 65572
rect 7432 65560 7438 65612
rect 21450 65560 21456 65612
rect 21508 65600 21514 65612
rect 52546 65600 52552 65612
rect 21508 65572 52552 65600
rect 21508 65560 21514 65572
rect 52546 65560 52552 65572
rect 52604 65600 52610 65612
rect 53558 65600 53564 65612
rect 52604 65572 53564 65600
rect 52604 65560 52610 65572
rect 53558 65560 53564 65572
rect 53616 65560 53622 65612
rect 74994 65560 75000 65612
rect 75052 65600 75058 65612
rect 81713 65603 81771 65609
rect 81713 65600 81725 65603
rect 75052 65572 81725 65600
rect 75052 65560 75058 65572
rect 81713 65569 81725 65572
rect 81759 65569 81771 65603
rect 81713 65563 81771 65569
rect 7101 65535 7159 65541
rect 7101 65501 7113 65535
rect 7147 65532 7159 65535
rect 25958 65532 25964 65544
rect 7147 65504 25964 65532
rect 7147 65501 7159 65504
rect 7101 65495 7159 65501
rect 25958 65492 25964 65504
rect 26016 65532 26022 65544
rect 33778 65532 33784 65544
rect 26016 65504 33784 65532
rect 26016 65492 26022 65504
rect 33778 65492 33784 65504
rect 33836 65492 33842 65544
rect 35434 65492 35440 65544
rect 35492 65532 35498 65544
rect 72694 65532 72700 65544
rect 35492 65504 72700 65532
rect 35492 65492 35498 65504
rect 72694 65492 72700 65504
rect 72752 65492 72758 65544
rect 81529 65467 81587 65473
rect 81529 65433 81541 65467
rect 81575 65464 81587 65467
rect 84562 65464 84568 65476
rect 81575 65436 84568 65464
rect 81575 65433 81587 65436
rect 81529 65427 81587 65433
rect 84562 65424 84568 65436
rect 84620 65464 84626 65476
rect 85390 65464 85396 65476
rect 84620 65436 85396 65464
rect 84620 65424 84626 65436
rect 85390 65424 85396 65436
rect 85448 65424 85454 65476
rect 44266 65356 44272 65408
rect 44324 65396 44330 65408
rect 45462 65396 45468 65408
rect 44324 65368 45468 65396
rect 44324 65356 44330 65368
rect 45462 65356 45468 65368
rect 45520 65356 45526 65408
rect 1104 65306 98808 65328
rect 1104 65254 4246 65306
rect 4298 65254 4310 65306
rect 4362 65254 4374 65306
rect 4426 65254 4438 65306
rect 4490 65254 34966 65306
rect 35018 65254 35030 65306
rect 35082 65254 35094 65306
rect 35146 65254 35158 65306
rect 35210 65254 65686 65306
rect 65738 65254 65750 65306
rect 65802 65254 65814 65306
rect 65866 65254 65878 65306
rect 65930 65254 96406 65306
rect 96458 65254 96470 65306
rect 96522 65254 96534 65306
rect 96586 65254 96598 65306
rect 96650 65254 98808 65306
rect 1104 65232 98808 65254
rect 80330 65192 80336 65204
rect 59648 65164 80336 65192
rect 46750 65016 46756 65068
rect 46808 65056 46814 65068
rect 59648 65056 59676 65164
rect 80330 65152 80336 65164
rect 80388 65152 80394 65204
rect 90542 65192 90548 65204
rect 90503 65164 90548 65192
rect 90542 65152 90548 65164
rect 90600 65152 90606 65204
rect 91186 65152 91192 65204
rect 91244 65192 91250 65204
rect 91244 65164 92428 65192
rect 91244 65152 91250 65164
rect 80149 65127 80207 65133
rect 46808 65028 59676 65056
rect 46808 65016 46814 65028
rect 27338 64948 27344 65000
rect 27396 64988 27402 65000
rect 27801 64991 27859 64997
rect 27801 64988 27813 64991
rect 27396 64960 27813 64988
rect 27396 64948 27402 64960
rect 27801 64957 27813 64960
rect 27847 64957 27859 64991
rect 27801 64951 27859 64957
rect 58894 64948 58900 65000
rect 58952 64988 58958 65000
rect 59265 64991 59323 64997
rect 59265 64988 59277 64991
rect 58952 64960 59277 64988
rect 58952 64948 58958 64960
rect 59265 64957 59277 64960
rect 59311 64957 59323 64991
rect 59446 64988 59452 65000
rect 59407 64960 59452 64988
rect 59265 64951 59323 64957
rect 59446 64948 59452 64960
rect 59504 64948 59510 65000
rect 59648 64997 59676 65028
rect 60016 65096 60734 65124
rect 60016 64997 60044 65096
rect 60274 65016 60280 65068
rect 60332 65056 60338 65068
rect 60369 65059 60427 65065
rect 60369 65056 60381 65059
rect 60332 65028 60381 65056
rect 60332 65016 60338 65028
rect 60369 65025 60381 65028
rect 60415 65025 60427 65059
rect 60706 65056 60734 65096
rect 80149 65093 80161 65127
rect 80195 65124 80207 65127
rect 80425 65127 80483 65133
rect 80425 65124 80437 65127
rect 80195 65096 80437 65124
rect 80195 65093 80207 65096
rect 80149 65087 80207 65093
rect 80425 65093 80437 65096
rect 80471 65124 80483 65127
rect 88334 65124 88340 65136
rect 80471 65096 88340 65124
rect 80471 65093 80483 65096
rect 80425 65087 80483 65093
rect 88334 65084 88340 65096
rect 88392 65084 88398 65136
rect 80882 65056 80888 65068
rect 60706 65028 80888 65056
rect 60369 65019 60427 65025
rect 80882 65016 80888 65028
rect 80940 65016 80946 65068
rect 90560 65056 90588 65152
rect 92400 65065 92428 65164
rect 92385 65059 92443 65065
rect 90560 65028 91048 65056
rect 59633 64991 59691 64997
rect 59633 64957 59645 64991
rect 59679 64957 59691 64991
rect 59633 64951 59691 64957
rect 60001 64991 60059 64997
rect 60001 64957 60013 64991
rect 60047 64957 60059 64991
rect 60182 64988 60188 65000
rect 60143 64960 60188 64988
rect 60001 64951 60059 64957
rect 9766 64880 9772 64932
rect 9824 64920 9830 64932
rect 11882 64920 11888 64932
rect 9824 64892 11888 64920
rect 9824 64880 9830 64892
rect 11882 64880 11888 64892
rect 11940 64880 11946 64932
rect 28626 64920 28632 64932
rect 28587 64892 28632 64920
rect 28626 64880 28632 64892
rect 28684 64880 28690 64932
rect 45462 64880 45468 64932
rect 45520 64920 45526 64932
rect 60016 64920 60044 64951
rect 60182 64948 60188 64960
rect 60240 64948 60246 65000
rect 90729 64991 90787 64997
rect 90729 64988 90741 64991
rect 60706 64960 80192 64988
rect 45520 64892 60044 64920
rect 45520 64880 45526 64892
rect 60550 64880 60556 64932
rect 60608 64920 60614 64932
rect 60706 64920 60734 64960
rect 60608 64892 60734 64920
rect 80164 64920 80192 64960
rect 84166 64960 90741 64988
rect 84166 64920 84194 64960
rect 90729 64957 90741 64960
rect 90775 64957 90787 64991
rect 91020 64988 91048 65028
rect 92385 65025 92397 65059
rect 92431 65025 92443 65059
rect 92385 65019 92443 65025
rect 92109 64991 92167 64997
rect 92109 64988 92121 64991
rect 91020 64960 92121 64988
rect 90729 64951 90787 64957
rect 92109 64957 92121 64960
rect 92155 64957 92167 64991
rect 92109 64951 92167 64957
rect 80164 64892 84194 64920
rect 60608 64880 60614 64892
rect 85390 64880 85396 64932
rect 85448 64920 85454 64932
rect 86954 64920 86960 64932
rect 85448 64892 86960 64920
rect 85448 64880 85454 64892
rect 86954 64880 86960 64892
rect 87012 64920 87018 64932
rect 91186 64920 91192 64932
rect 87012 64892 91192 64920
rect 87012 64880 87018 64892
rect 91186 64880 91192 64892
rect 91244 64880 91250 64932
rect 39666 64812 39672 64864
rect 39724 64852 39730 64864
rect 81710 64852 81716 64864
rect 39724 64824 81716 64852
rect 39724 64812 39730 64824
rect 81710 64812 81716 64824
rect 81768 64812 81774 64864
rect 1104 64762 98808 64784
rect 1104 64710 19606 64762
rect 19658 64710 19670 64762
rect 19722 64710 19734 64762
rect 19786 64710 19798 64762
rect 19850 64710 50326 64762
rect 50378 64710 50390 64762
rect 50442 64710 50454 64762
rect 50506 64710 50518 64762
rect 50570 64710 81046 64762
rect 81098 64710 81110 64762
rect 81162 64710 81174 64762
rect 81226 64710 81238 64762
rect 81290 64710 98808 64762
rect 1104 64688 98808 64710
rect 27338 64648 27344 64660
rect 27299 64620 27344 64648
rect 27338 64608 27344 64620
rect 27396 64608 27402 64660
rect 49694 64608 49700 64660
rect 49752 64648 49758 64660
rect 50525 64651 50583 64657
rect 50525 64648 50537 64651
rect 49752 64620 50537 64648
rect 49752 64608 49758 64620
rect 50525 64617 50537 64620
rect 50571 64617 50583 64651
rect 50525 64611 50583 64617
rect 50982 64608 50988 64660
rect 51040 64648 51046 64660
rect 51040 64620 95464 64648
rect 51040 64608 51046 64620
rect 16022 64472 16028 64524
rect 16080 64512 16086 64524
rect 27157 64515 27215 64521
rect 27157 64512 27169 64515
rect 16080 64484 27169 64512
rect 16080 64472 16086 64484
rect 27157 64481 27169 64484
rect 27203 64481 27215 64515
rect 49418 64512 49424 64524
rect 49379 64484 49424 64512
rect 27157 64475 27215 64481
rect 49418 64472 49424 64484
rect 49476 64472 49482 64524
rect 49712 64521 49740 64608
rect 50062 64580 50068 64592
rect 49988 64552 50068 64580
rect 49988 64521 50016 64552
rect 50062 64540 50068 64552
rect 50120 64540 50126 64592
rect 50338 64580 50344 64592
rect 50264 64552 50344 64580
rect 50264 64521 50292 64552
rect 50338 64540 50344 64552
rect 50396 64580 50402 64592
rect 80238 64580 80244 64592
rect 50396 64552 80244 64580
rect 50396 64540 50402 64552
rect 80238 64540 80244 64552
rect 80296 64540 80302 64592
rect 91572 64552 92060 64580
rect 49703 64515 49761 64521
rect 49703 64481 49715 64515
rect 49749 64481 49761 64515
rect 49703 64475 49761 64481
rect 49880 64515 49938 64521
rect 49880 64481 49892 64515
rect 49926 64481 49938 64515
rect 49880 64475 49938 64481
rect 49973 64515 50031 64521
rect 49973 64481 49985 64515
rect 50019 64481 50031 64515
rect 49973 64475 50031 64481
rect 50249 64515 50307 64521
rect 50249 64481 50261 64515
rect 50295 64481 50307 64515
rect 50249 64475 50307 64481
rect 49510 64404 49516 64456
rect 49568 64444 49574 64456
rect 49895 64444 49923 64475
rect 55306 64472 55312 64524
rect 55364 64512 55370 64524
rect 56042 64512 56048 64524
rect 55364 64484 56048 64512
rect 55364 64472 55370 64484
rect 56042 64472 56048 64484
rect 56100 64512 56106 64524
rect 91572 64521 91600 64552
rect 91557 64515 91615 64521
rect 91557 64512 91569 64515
rect 56100 64484 91569 64512
rect 56100 64472 56106 64484
rect 91557 64481 91569 64484
rect 91603 64481 91615 64515
rect 91738 64512 91744 64524
rect 91699 64484 91744 64512
rect 91557 64475 91615 64481
rect 91738 64472 91744 64484
rect 91796 64472 91802 64524
rect 91830 64472 91836 64524
rect 91888 64512 91894 64524
rect 92032 64521 92060 64552
rect 92017 64515 92075 64521
rect 91888 64484 91933 64512
rect 91888 64472 91894 64484
rect 92017 64481 92029 64515
rect 92063 64481 92075 64515
rect 95050 64512 95056 64524
rect 95011 64484 95056 64512
rect 92017 64475 92075 64481
rect 95050 64472 95056 64484
rect 95108 64472 95114 64524
rect 95436 64521 95464 64620
rect 95421 64515 95479 64521
rect 95421 64481 95433 64515
rect 95467 64481 95479 64515
rect 95786 64512 95792 64524
rect 95747 64484 95792 64512
rect 95421 64475 95479 64481
rect 95786 64472 95792 64484
rect 95844 64472 95850 64524
rect 49568 64416 49923 64444
rect 50065 64447 50123 64453
rect 49568 64404 49574 64416
rect 50065 64413 50077 64447
rect 50111 64413 50123 64447
rect 50065 64407 50123 64413
rect 29546 64336 29552 64388
rect 29604 64376 29610 64388
rect 49878 64376 49884 64388
rect 29604 64348 49884 64376
rect 29604 64336 29610 64348
rect 49878 64336 49884 64348
rect 49936 64336 49942 64388
rect 26145 64311 26203 64317
rect 26145 64277 26157 64311
rect 26191 64308 26203 64311
rect 26418 64308 26424 64320
rect 26191 64280 26424 64308
rect 26191 64277 26203 64280
rect 26145 64271 26203 64277
rect 26418 64268 26424 64280
rect 26476 64268 26482 64320
rect 49605 64311 49663 64317
rect 49605 64277 49617 64311
rect 49651 64308 49663 64311
rect 49970 64308 49976 64320
rect 49651 64280 49976 64308
rect 49651 64277 49663 64280
rect 49605 64271 49663 64277
rect 49970 64268 49976 64280
rect 50028 64308 50034 64320
rect 50080 64308 50108 64407
rect 75362 64404 75368 64456
rect 75420 64444 75426 64456
rect 75822 64444 75828 64456
rect 75420 64416 75828 64444
rect 75420 64404 75426 64416
rect 75822 64404 75828 64416
rect 75880 64404 75886 64456
rect 87690 64404 87696 64456
rect 87748 64444 87754 64456
rect 92201 64447 92259 64453
rect 92201 64444 92213 64447
rect 87748 64416 92213 64444
rect 87748 64404 87754 64416
rect 92201 64413 92213 64416
rect 92247 64413 92259 64447
rect 95234 64444 95240 64456
rect 95195 64416 95240 64444
rect 92201 64407 92259 64413
rect 95234 64404 95240 64416
rect 95292 64404 95298 64456
rect 95697 64447 95755 64453
rect 95697 64413 95709 64447
rect 95743 64413 95755 64447
rect 95697 64407 95755 64413
rect 50246 64336 50252 64388
rect 50304 64376 50310 64388
rect 50304 64348 91784 64376
rect 50304 64336 50310 64348
rect 50028 64280 50108 64308
rect 50028 64268 50034 64280
rect 50154 64268 50160 64320
rect 50212 64308 50218 64320
rect 50341 64311 50399 64317
rect 50341 64308 50353 64311
rect 50212 64280 50353 64308
rect 50212 64268 50218 64280
rect 50341 64277 50353 64280
rect 50387 64277 50399 64311
rect 50341 64271 50399 64277
rect 50890 64268 50896 64320
rect 50948 64308 50954 64320
rect 51442 64308 51448 64320
rect 50948 64280 51448 64308
rect 50948 64268 50954 64280
rect 51442 64268 51448 64280
rect 51500 64268 51506 64320
rect 67082 64268 67088 64320
rect 67140 64308 67146 64320
rect 67177 64311 67235 64317
rect 67177 64308 67189 64311
rect 67140 64280 67189 64308
rect 67140 64268 67146 64280
rect 67177 64277 67189 64280
rect 67223 64308 67235 64311
rect 67361 64311 67419 64317
rect 67361 64308 67373 64311
rect 67223 64280 67373 64308
rect 67223 64277 67235 64280
rect 67177 64271 67235 64277
rect 67361 64277 67373 64280
rect 67407 64277 67419 64311
rect 91756 64308 91784 64348
rect 92750 64336 92756 64388
rect 92808 64376 92814 64388
rect 95712 64376 95740 64407
rect 92808 64348 95740 64376
rect 92808 64336 92814 64348
rect 96249 64311 96307 64317
rect 96249 64308 96261 64311
rect 91756 64280 96261 64308
rect 67361 64271 67419 64277
rect 96249 64277 96261 64280
rect 96295 64277 96307 64311
rect 96249 64271 96307 64277
rect 1104 64218 98808 64240
rect 1104 64166 4246 64218
rect 4298 64166 4310 64218
rect 4362 64166 4374 64218
rect 4426 64166 4438 64218
rect 4490 64166 34966 64218
rect 35018 64166 35030 64218
rect 35082 64166 35094 64218
rect 35146 64166 35158 64218
rect 35210 64166 65686 64218
rect 65738 64166 65750 64218
rect 65802 64166 65814 64218
rect 65866 64166 65878 64218
rect 65930 64166 96406 64218
rect 96458 64166 96470 64218
rect 96522 64166 96534 64218
rect 96586 64166 96598 64218
rect 96650 64166 98808 64218
rect 1104 64144 98808 64166
rect 8938 64104 8944 64116
rect 8496 64076 8800 64104
rect 8899 64076 8944 64104
rect 8294 63900 8300 63912
rect 8255 63872 8300 63900
rect 8294 63860 8300 63872
rect 8352 63860 8358 63912
rect 8496 63909 8524 64076
rect 8662 63996 8668 64048
rect 8720 63996 8726 64048
rect 8680 63909 8708 63996
rect 8772 63968 8800 64076
rect 8938 64064 8944 64076
rect 8996 64064 9002 64116
rect 34146 64064 34152 64116
rect 34204 64104 34210 64116
rect 34204 64076 49556 64104
rect 34204 64064 34210 64076
rect 14274 63996 14280 64048
rect 14332 64036 14338 64048
rect 49418 64036 49424 64048
rect 14332 64008 49424 64036
rect 14332 63996 14338 64008
rect 49418 63996 49424 64008
rect 49476 63996 49482 64048
rect 49528 64036 49556 64076
rect 49694 64064 49700 64116
rect 49752 64104 49758 64116
rect 50890 64104 50896 64116
rect 49752 64076 50896 64104
rect 49752 64064 49758 64076
rect 50890 64064 50896 64076
rect 50948 64064 50954 64116
rect 61930 64064 61936 64116
rect 61988 64104 61994 64116
rect 66346 64104 66352 64116
rect 61988 64076 66352 64104
rect 61988 64064 61994 64076
rect 66346 64064 66352 64076
rect 66404 64064 66410 64116
rect 68462 64104 68468 64116
rect 66916 64076 68324 64104
rect 68423 64076 68468 64104
rect 49970 64036 49976 64048
rect 49528 64008 49976 64036
rect 49970 63996 49976 64008
rect 50028 64036 50034 64048
rect 52454 64036 52460 64048
rect 50028 64008 52460 64036
rect 50028 63996 50034 64008
rect 52454 63996 52460 64008
rect 52512 64036 52518 64048
rect 53006 64036 53012 64048
rect 52512 64008 53012 64036
rect 52512 63996 52518 64008
rect 53006 63996 53012 64008
rect 53064 63996 53070 64048
rect 8772 63940 16574 63968
rect 8480 63903 8538 63909
rect 8480 63869 8492 63903
rect 8526 63869 8538 63903
rect 8480 63863 8538 63869
rect 8573 63903 8631 63909
rect 8573 63869 8585 63903
rect 8619 63869 8631 63903
rect 8573 63863 8631 63869
rect 8665 63903 8723 63909
rect 8665 63869 8677 63903
rect 8711 63869 8723 63903
rect 8665 63863 8723 63869
rect 8849 63903 8907 63909
rect 8849 63869 8861 63903
rect 8895 63900 8907 63903
rect 16546 63900 16574 63940
rect 40770 63928 40776 63980
rect 40828 63968 40834 63980
rect 62666 63968 62672 63980
rect 40828 63940 62672 63968
rect 40828 63928 40834 63940
rect 62666 63928 62672 63940
rect 62724 63928 62730 63980
rect 54846 63900 54852 63912
rect 8895 63872 12434 63900
rect 16546 63872 54852 63900
rect 8895 63869 8907 63872
rect 8849 63863 8907 63869
rect 8588 63764 8616 63863
rect 12406 63832 12434 63872
rect 54846 63860 54852 63872
rect 54904 63860 54910 63912
rect 66533 63903 66591 63909
rect 66533 63869 66545 63903
rect 66579 63900 66591 63903
rect 66916 63900 66944 64076
rect 66990 63996 66996 64048
rect 67048 64036 67054 64048
rect 68296 64036 68324 64076
rect 68462 64064 68468 64076
rect 68520 64064 68526 64116
rect 74994 64104 75000 64116
rect 70366 64076 75000 64104
rect 70366 64036 70394 64076
rect 74994 64064 75000 64076
rect 75052 64064 75058 64116
rect 67048 64008 67128 64036
rect 68296 64008 70394 64036
rect 67048 63996 67054 64008
rect 67100 63977 67128 64008
rect 75270 63996 75276 64048
rect 75328 64036 75334 64048
rect 82446 64036 82452 64048
rect 75328 64008 82308 64036
rect 82407 64008 82452 64036
rect 75328 63996 75334 64008
rect 67085 63971 67143 63977
rect 67085 63937 67097 63971
rect 67131 63937 67143 63971
rect 67085 63931 67143 63937
rect 67266 63928 67272 63980
rect 67324 63968 67330 63980
rect 67324 63940 82216 63968
rect 67324 63928 67330 63940
rect 67361 63903 67419 63909
rect 67361 63900 67373 63903
rect 66579 63872 66944 63900
rect 67008 63872 67373 63900
rect 66579 63869 66591 63872
rect 66533 63863 66591 63869
rect 24118 63832 24124 63844
rect 12406 63804 24124 63832
rect 24118 63792 24124 63804
rect 24176 63792 24182 63844
rect 33778 63792 33784 63844
rect 33836 63832 33842 63844
rect 49694 63832 49700 63844
rect 33836 63804 49700 63832
rect 33836 63792 33842 63804
rect 49694 63792 49700 63804
rect 49752 63792 49758 63844
rect 45370 63764 45376 63776
rect 8588 63736 45376 63764
rect 45370 63724 45376 63736
rect 45428 63724 45434 63776
rect 47946 63724 47952 63776
rect 48004 63764 48010 63776
rect 66901 63767 66959 63773
rect 66901 63764 66913 63767
rect 48004 63736 66913 63764
rect 48004 63724 48010 63736
rect 66901 63733 66913 63736
rect 66947 63764 66959 63767
rect 67008 63764 67036 63872
rect 67361 63869 67373 63872
rect 67407 63869 67419 63903
rect 67361 63863 67419 63869
rect 75362 63860 75368 63912
rect 75420 63900 75426 63912
rect 82188 63909 82216 63940
rect 82280 63909 82308 64008
rect 82446 63996 82452 64008
rect 82504 63996 82510 64048
rect 81897 63903 81955 63909
rect 81897 63900 81909 63903
rect 75420 63872 81909 63900
rect 75420 63860 75426 63872
rect 81897 63869 81909 63872
rect 81943 63869 81955 63903
rect 81897 63863 81955 63869
rect 82173 63903 82231 63909
rect 82173 63869 82185 63903
rect 82219 63869 82231 63903
rect 82173 63863 82231 63869
rect 82270 63903 82328 63909
rect 82270 63869 82282 63903
rect 82316 63869 82328 63903
rect 82270 63863 82328 63869
rect 93121 63903 93179 63909
rect 93121 63869 93133 63903
rect 93167 63869 93179 63903
rect 93121 63863 93179 63869
rect 71682 63832 71688 63844
rect 70366 63804 71688 63832
rect 66947 63736 67036 63764
rect 66947 63733 66959 63736
rect 66901 63727 66959 63733
rect 67450 63724 67456 63776
rect 67508 63764 67514 63776
rect 70366 63764 70394 63804
rect 71682 63792 71688 63804
rect 71740 63832 71746 63844
rect 78858 63832 78864 63844
rect 71740 63804 78864 63832
rect 71740 63792 71746 63804
rect 78858 63792 78864 63804
rect 78916 63792 78922 63844
rect 81710 63792 81716 63844
rect 81768 63832 81774 63844
rect 82081 63835 82139 63841
rect 82081 63832 82093 63835
rect 81768 63804 82093 63832
rect 81768 63792 81774 63804
rect 82081 63801 82093 63804
rect 82127 63801 82139 63835
rect 82188 63832 82216 63863
rect 92750 63832 92756 63844
rect 82188 63804 92756 63832
rect 82081 63795 82139 63801
rect 92750 63792 92756 63804
rect 92808 63792 92814 63844
rect 92934 63764 92940 63776
rect 67508 63736 70394 63764
rect 92895 63736 92940 63764
rect 67508 63724 67514 63736
rect 92934 63724 92940 63736
rect 92992 63764 92998 63776
rect 93136 63764 93164 63863
rect 92992 63736 93164 63764
rect 92992 63724 92998 63736
rect 1104 63674 98808 63696
rect 1104 63622 19606 63674
rect 19658 63622 19670 63674
rect 19722 63622 19734 63674
rect 19786 63622 19798 63674
rect 19850 63622 50326 63674
rect 50378 63622 50390 63674
rect 50442 63622 50454 63674
rect 50506 63622 50518 63674
rect 50570 63622 81046 63674
rect 81098 63622 81110 63674
rect 81162 63622 81174 63674
rect 81226 63622 81238 63674
rect 81290 63622 98808 63674
rect 1104 63600 98808 63622
rect 28350 63520 28356 63572
rect 28408 63560 28414 63572
rect 34146 63560 34152 63572
rect 28408 63532 34152 63560
rect 28408 63520 28414 63532
rect 34146 63520 34152 63532
rect 34204 63520 34210 63572
rect 45462 63520 45468 63572
rect 45520 63560 45526 63572
rect 50982 63560 50988 63572
rect 45520 63532 50988 63560
rect 45520 63520 45526 63532
rect 50982 63520 50988 63532
rect 51040 63520 51046 63572
rect 48958 63452 48964 63504
rect 49016 63492 49022 63504
rect 49510 63492 49516 63504
rect 49016 63464 49516 63492
rect 49016 63452 49022 63464
rect 49510 63452 49516 63464
rect 49568 63452 49574 63504
rect 8386 63384 8392 63436
rect 8444 63424 8450 63436
rect 18601 63427 18659 63433
rect 18601 63424 18613 63427
rect 8444 63396 18613 63424
rect 8444 63384 8450 63396
rect 18601 63393 18613 63396
rect 18647 63424 18659 63427
rect 19334 63424 19340 63436
rect 18647 63396 19340 63424
rect 18647 63393 18659 63396
rect 18601 63387 18659 63393
rect 19334 63384 19340 63396
rect 19392 63384 19398 63436
rect 27433 63427 27491 63433
rect 27433 63393 27445 63427
rect 27479 63424 27491 63427
rect 28350 63424 28356 63436
rect 27479 63396 28356 63424
rect 27479 63393 27491 63396
rect 27433 63387 27491 63393
rect 28350 63384 28356 63396
rect 28408 63384 28414 63436
rect 57054 63316 57060 63368
rect 57112 63356 57118 63368
rect 57790 63356 57796 63368
rect 57112 63328 57796 63356
rect 57112 63316 57118 63328
rect 57790 63316 57796 63328
rect 57848 63316 57854 63368
rect 15470 63248 15476 63300
rect 15528 63288 15534 63300
rect 27246 63288 27252 63300
rect 15528 63260 26234 63288
rect 27207 63260 27252 63288
rect 15528 63248 15534 63260
rect 9401 63223 9459 63229
rect 9401 63189 9413 63223
rect 9447 63220 9459 63223
rect 9677 63223 9735 63229
rect 9677 63220 9689 63223
rect 9447 63192 9689 63220
rect 9447 63189 9459 63192
rect 9401 63183 9459 63189
rect 9677 63189 9689 63192
rect 9723 63220 9735 63223
rect 11974 63220 11980 63232
rect 9723 63192 11980 63220
rect 9723 63189 9735 63192
rect 9677 63183 9735 63189
rect 11974 63180 11980 63192
rect 12032 63180 12038 63232
rect 18690 63180 18696 63232
rect 18748 63220 18754 63232
rect 18785 63223 18843 63229
rect 18785 63220 18797 63223
rect 18748 63192 18797 63220
rect 18748 63180 18754 63192
rect 18785 63189 18797 63192
rect 18831 63189 18843 63223
rect 26206 63220 26234 63260
rect 27246 63248 27252 63260
rect 27304 63248 27310 63300
rect 34238 63220 34244 63232
rect 26206 63192 34244 63220
rect 18785 63183 18843 63189
rect 34238 63180 34244 63192
rect 34296 63180 34302 63232
rect 44637 63223 44695 63229
rect 44637 63189 44649 63223
rect 44683 63220 44695 63223
rect 44913 63223 44971 63229
rect 44913 63220 44925 63223
rect 44683 63192 44925 63220
rect 44683 63189 44695 63192
rect 44637 63183 44695 63189
rect 44913 63189 44925 63192
rect 44959 63220 44971 63223
rect 53098 63220 53104 63232
rect 44959 63192 53104 63220
rect 44959 63189 44971 63192
rect 44913 63183 44971 63189
rect 53098 63180 53104 63192
rect 53156 63180 53162 63232
rect 79686 63220 79692 63232
rect 79647 63192 79692 63220
rect 79686 63180 79692 63192
rect 79744 63220 79750 63232
rect 79873 63223 79931 63229
rect 79873 63220 79885 63223
rect 79744 63192 79885 63220
rect 79744 63180 79750 63192
rect 79873 63189 79885 63192
rect 79919 63189 79931 63223
rect 79873 63183 79931 63189
rect 1104 63130 98808 63152
rect 1104 63078 4246 63130
rect 4298 63078 4310 63130
rect 4362 63078 4374 63130
rect 4426 63078 4438 63130
rect 4490 63078 34966 63130
rect 35018 63078 35030 63130
rect 35082 63078 35094 63130
rect 35146 63078 35158 63130
rect 35210 63078 65686 63130
rect 65738 63078 65750 63130
rect 65802 63078 65814 63130
rect 65866 63078 65878 63130
rect 65930 63078 96406 63130
rect 96458 63078 96470 63130
rect 96522 63078 96534 63130
rect 96586 63078 96598 63130
rect 96650 63078 98808 63130
rect 1104 63056 98808 63078
rect 22094 63016 22100 63028
rect 16546 62988 22100 63016
rect 13541 62951 13599 62957
rect 13541 62917 13553 62951
rect 13587 62948 13599 62951
rect 14734 62948 14740 62960
rect 13587 62920 14740 62948
rect 13587 62917 13599 62920
rect 13541 62911 13599 62917
rect 14734 62908 14740 62920
rect 14792 62908 14798 62960
rect 14185 62883 14243 62889
rect 14185 62849 14197 62883
rect 14231 62880 14243 62883
rect 15654 62880 15660 62892
rect 14231 62852 15660 62880
rect 14231 62849 14243 62852
rect 14185 62843 14243 62849
rect 15654 62840 15660 62852
rect 15712 62840 15718 62892
rect 13725 62815 13783 62821
rect 13725 62781 13737 62815
rect 13771 62781 13783 62815
rect 13725 62775 13783 62781
rect 14093 62815 14151 62821
rect 14093 62781 14105 62815
rect 14139 62812 14151 62815
rect 16546 62812 16574 62988
rect 22094 62976 22100 62988
rect 22152 63016 22158 63028
rect 37826 63016 37832 63028
rect 22152 62988 37832 63016
rect 22152 62976 22158 62988
rect 37826 62976 37832 62988
rect 37884 62976 37890 63028
rect 20622 62908 20628 62960
rect 20680 62948 20686 62960
rect 57330 62948 57336 62960
rect 20680 62920 57336 62948
rect 20680 62908 20686 62920
rect 57330 62908 57336 62920
rect 57388 62908 57394 62960
rect 20438 62840 20444 62892
rect 20496 62880 20502 62892
rect 60918 62880 60924 62892
rect 20496 62852 60924 62880
rect 20496 62840 20502 62852
rect 60918 62840 60924 62852
rect 60976 62840 60982 62892
rect 33778 62812 33784 62824
rect 14139 62784 16574 62812
rect 33739 62784 33784 62812
rect 14139 62781 14151 62784
rect 14093 62775 14151 62781
rect 12986 62704 12992 62756
rect 13044 62744 13050 62756
rect 13740 62744 13768 62775
rect 33778 62772 33784 62784
rect 33836 62772 33842 62824
rect 33964 62815 34022 62821
rect 33964 62781 33976 62815
rect 34010 62781 34022 62815
rect 33964 62775 34022 62781
rect 34057 62815 34115 62821
rect 34057 62781 34069 62815
rect 34103 62781 34115 62815
rect 34057 62775 34115 62781
rect 15470 62744 15476 62756
rect 13044 62716 15476 62744
rect 13044 62704 13050 62716
rect 15470 62704 15476 62716
rect 15528 62704 15534 62756
rect 33686 62676 33692 62688
rect 33647 62648 33692 62676
rect 33686 62636 33692 62648
rect 33744 62636 33750 62688
rect 33980 62676 34008 62775
rect 34072 62744 34100 62775
rect 34146 62772 34152 62824
rect 34204 62812 34210 62824
rect 34333 62815 34391 62821
rect 34204 62784 34249 62812
rect 34204 62772 34210 62784
rect 34333 62781 34345 62815
rect 34379 62812 34391 62815
rect 34514 62812 34520 62824
rect 34379 62784 34520 62812
rect 34379 62781 34391 62784
rect 34333 62775 34391 62781
rect 34514 62772 34520 62784
rect 34572 62812 34578 62824
rect 35802 62812 35808 62824
rect 34572 62784 35808 62812
rect 34572 62772 34578 62784
rect 35802 62772 35808 62784
rect 35860 62812 35866 62824
rect 93486 62812 93492 62824
rect 35860 62784 93492 62812
rect 35860 62772 35866 62784
rect 93486 62772 93492 62784
rect 93544 62772 93550 62824
rect 34238 62744 34244 62756
rect 34072 62716 34244 62744
rect 34238 62704 34244 62716
rect 34296 62704 34302 62756
rect 34146 62676 34152 62688
rect 33980 62648 34152 62676
rect 34146 62636 34152 62648
rect 34204 62636 34210 62688
rect 34330 62636 34336 62688
rect 34388 62676 34394 62688
rect 34425 62679 34483 62685
rect 34425 62676 34437 62679
rect 34388 62648 34437 62676
rect 34388 62636 34394 62648
rect 34425 62645 34437 62648
rect 34471 62645 34483 62679
rect 34425 62639 34483 62645
rect 1104 62586 98808 62608
rect 1104 62534 19606 62586
rect 19658 62534 19670 62586
rect 19722 62534 19734 62586
rect 19786 62534 19798 62586
rect 19850 62534 50326 62586
rect 50378 62534 50390 62586
rect 50442 62534 50454 62586
rect 50506 62534 50518 62586
rect 50570 62534 81046 62586
rect 81098 62534 81110 62586
rect 81162 62534 81174 62586
rect 81226 62534 81238 62586
rect 81290 62534 98808 62586
rect 1104 62512 98808 62534
rect 33686 62432 33692 62484
rect 33744 62472 33750 62484
rect 34514 62472 34520 62484
rect 33744 62444 34520 62472
rect 33744 62432 33750 62444
rect 34514 62432 34520 62444
rect 34572 62432 34578 62484
rect 60706 62444 74948 62472
rect 32398 62404 32404 62416
rect 13188 62376 32404 62404
rect 13188 62348 13216 62376
rect 32398 62364 32404 62376
rect 32456 62364 32462 62416
rect 34146 62364 34152 62416
rect 34204 62404 34210 62416
rect 34790 62404 34796 62416
rect 34204 62376 34796 62404
rect 34204 62364 34210 62376
rect 34790 62364 34796 62376
rect 34848 62364 34854 62416
rect 53558 62364 53564 62416
rect 53616 62404 53622 62416
rect 60706 62404 60734 62444
rect 53616 62376 60734 62404
rect 53616 62364 53622 62376
rect 65702 62364 65708 62416
rect 65760 62404 65766 62416
rect 72418 62404 72424 62416
rect 65760 62376 72424 62404
rect 65760 62364 65766 62376
rect 72418 62364 72424 62376
rect 72476 62364 72482 62416
rect 74092 62376 74764 62404
rect 12986 62336 12992 62348
rect 12947 62308 12992 62336
rect 12986 62296 12992 62308
rect 13044 62296 13050 62348
rect 13170 62336 13176 62348
rect 13131 62308 13176 62336
rect 13170 62296 13176 62308
rect 13228 62296 13234 62348
rect 13265 62339 13323 62345
rect 13265 62305 13277 62339
rect 13311 62336 13323 62339
rect 15838 62336 15844 62348
rect 13311 62308 15844 62336
rect 13311 62305 13323 62308
rect 13265 62299 13323 62305
rect 6454 62228 6460 62280
rect 6512 62268 6518 62280
rect 13280 62268 13308 62299
rect 15838 62296 15844 62308
rect 15896 62296 15902 62348
rect 49602 62296 49608 62348
rect 49660 62336 49666 62348
rect 65610 62336 65616 62348
rect 49660 62308 65616 62336
rect 49660 62296 49666 62308
rect 65610 62296 65616 62308
rect 65668 62296 65674 62348
rect 65794 62296 65800 62348
rect 65852 62336 65858 62348
rect 73982 62336 73988 62348
rect 65852 62308 73988 62336
rect 65852 62296 65858 62308
rect 73982 62296 73988 62308
rect 74040 62296 74046 62348
rect 6512 62240 13308 62268
rect 6512 62228 6518 62240
rect 49510 62228 49516 62280
rect 49568 62268 49574 62280
rect 65702 62268 65708 62280
rect 49568 62240 65708 62268
rect 49568 62228 49574 62240
rect 65702 62228 65708 62240
rect 65760 62228 65766 62280
rect 70302 62228 70308 62280
rect 70360 62268 70366 62280
rect 74092 62268 74120 62376
rect 74353 62339 74411 62345
rect 74353 62305 74365 62339
rect 74399 62336 74411 62339
rect 74442 62336 74448 62348
rect 74399 62308 74448 62336
rect 74399 62305 74411 62308
rect 74353 62299 74411 62305
rect 74442 62296 74448 62308
rect 74500 62296 74506 62348
rect 74736 62345 74764 62376
rect 74920 62345 74948 62444
rect 74721 62339 74779 62345
rect 74721 62305 74733 62339
rect 74767 62305 74779 62339
rect 74721 62299 74779 62305
rect 74905 62339 74963 62345
rect 74905 62305 74917 62339
rect 74951 62305 74963 62339
rect 83458 62336 83464 62348
rect 83419 62308 83464 62336
rect 74905 62299 74963 62305
rect 83458 62296 83464 62308
rect 83516 62296 83522 62348
rect 74258 62268 74264 62280
rect 70360 62240 74120 62268
rect 74219 62240 74264 62268
rect 70360 62228 70366 62240
rect 74258 62228 74264 62240
rect 74316 62228 74322 62280
rect 83737 62271 83795 62277
rect 83737 62268 83749 62271
rect 80026 62240 83749 62268
rect 39942 62160 39948 62212
rect 40000 62200 40006 62212
rect 75089 62203 75147 62209
rect 75089 62200 75101 62203
rect 40000 62172 75101 62200
rect 40000 62160 40006 62172
rect 75089 62169 75101 62172
rect 75135 62169 75147 62203
rect 75089 62163 75147 62169
rect 12805 62135 12863 62141
rect 12805 62101 12817 62135
rect 12851 62132 12863 62135
rect 15102 62132 15108 62144
rect 12851 62104 15108 62132
rect 12851 62101 12863 62104
rect 12805 62095 12863 62101
rect 15102 62092 15108 62104
rect 15160 62092 15166 62144
rect 36630 62092 36636 62144
rect 36688 62132 36694 62144
rect 45462 62132 45468 62144
rect 36688 62104 45468 62132
rect 36688 62092 36694 62104
rect 45462 62092 45468 62104
rect 45520 62092 45526 62144
rect 72418 62092 72424 62144
rect 72476 62132 72482 62144
rect 80026 62132 80054 62240
rect 83737 62237 83749 62240
rect 83783 62237 83795 62271
rect 83737 62231 83795 62237
rect 72476 62104 80054 62132
rect 72476 62092 72482 62104
rect 1104 62042 98808 62064
rect 1104 61990 4246 62042
rect 4298 61990 4310 62042
rect 4362 61990 4374 62042
rect 4426 61990 4438 62042
rect 4490 61990 34966 62042
rect 35018 61990 35030 62042
rect 35082 61990 35094 62042
rect 35146 61990 35158 62042
rect 35210 61990 65686 62042
rect 65738 61990 65750 62042
rect 65802 61990 65814 62042
rect 65866 61990 65878 62042
rect 65930 61990 96406 62042
rect 96458 61990 96470 62042
rect 96522 61990 96534 62042
rect 96586 61990 96598 62042
rect 96650 61990 98808 62042
rect 1104 61968 98808 61990
rect 57514 61928 57520 61940
rect 41386 61900 57520 61928
rect 30650 61792 30656 61804
rect 30611 61764 30656 61792
rect 30650 61752 30656 61764
rect 30708 61752 30714 61804
rect 41386 61792 41414 61900
rect 57514 61888 57520 61900
rect 57572 61888 57578 61940
rect 58618 61888 58624 61940
rect 58676 61928 58682 61940
rect 74994 61928 75000 61940
rect 58676 61900 60734 61928
rect 74955 61900 75000 61928
rect 58676 61888 58682 61900
rect 60706 61860 60734 61900
rect 74994 61888 75000 61900
rect 75052 61888 75058 61940
rect 77938 61860 77944 61872
rect 60706 61832 77944 61860
rect 77938 61820 77944 61832
rect 77996 61860 78002 61872
rect 77996 61832 80054 61860
rect 77996 61820 78002 61832
rect 31220 61764 41414 61792
rect 50709 61795 50767 61801
rect 30469 61727 30527 61733
rect 30469 61693 30481 61727
rect 30515 61693 30527 61727
rect 30834 61724 30840 61736
rect 30795 61696 30840 61724
rect 30469 61687 30527 61693
rect 30484 61656 30512 61687
rect 30834 61684 30840 61696
rect 30892 61684 30898 61736
rect 31220 61733 31248 61764
rect 50709 61761 50721 61795
rect 50755 61792 50767 61795
rect 54202 61792 54208 61804
rect 50755 61764 54208 61792
rect 50755 61761 50767 61764
rect 50709 61755 50767 61761
rect 54202 61752 54208 61764
rect 54260 61792 54266 61804
rect 57422 61792 57428 61804
rect 54260 61764 57428 61792
rect 54260 61752 54266 61764
rect 57422 61752 57428 61764
rect 57480 61752 57486 61804
rect 31205 61727 31263 61733
rect 31205 61693 31217 61727
rect 31251 61693 31263 61727
rect 31386 61724 31392 61736
rect 31347 61696 31392 61724
rect 31205 61687 31263 61693
rect 31386 61684 31392 61696
rect 31444 61684 31450 61736
rect 48774 61724 48780 61736
rect 48735 61696 48780 61724
rect 48774 61684 48780 61696
rect 48832 61684 48838 61736
rect 50982 61724 50988 61736
rect 50943 61696 50988 61724
rect 50982 61684 50988 61696
rect 51040 61684 51046 61736
rect 71314 61684 71320 61736
rect 71372 61724 71378 61736
rect 75181 61727 75239 61733
rect 75181 61724 75193 61727
rect 71372 61696 75193 61724
rect 71372 61684 71378 61696
rect 75181 61693 75193 61696
rect 75227 61693 75239 61727
rect 80026 61724 80054 61832
rect 83277 61727 83335 61733
rect 83277 61724 83289 61727
rect 80026 61696 83289 61724
rect 75181 61687 75239 61693
rect 83277 61693 83289 61696
rect 83323 61693 83335 61727
rect 83277 61687 83335 61693
rect 90818 61684 90824 61736
rect 90876 61724 90882 61736
rect 93213 61727 93271 61733
rect 93213 61724 93225 61727
rect 90876 61696 93225 61724
rect 90876 61684 90882 61696
rect 93213 61693 93225 61696
rect 93259 61693 93271 61727
rect 93213 61687 93271 61693
rect 44542 61656 44548 61668
rect 30484 61628 44548 61656
rect 44542 61616 44548 61628
rect 44600 61616 44606 61668
rect 49602 61656 49608 61668
rect 49563 61628 49608 61656
rect 49602 61616 49608 61628
rect 49660 61616 49666 61668
rect 83458 61616 83464 61668
rect 83516 61656 83522 61668
rect 83645 61659 83703 61665
rect 83645 61656 83657 61659
rect 83516 61628 83657 61656
rect 83516 61616 83522 61628
rect 83645 61625 83657 61628
rect 83691 61656 83703 61659
rect 84930 61656 84936 61668
rect 83691 61628 84936 61656
rect 83691 61625 83703 61628
rect 83645 61619 83703 61625
rect 84930 61616 84936 61628
rect 84988 61616 84994 61668
rect 31662 61588 31668 61600
rect 31623 61560 31668 61588
rect 31662 61548 31668 61560
rect 31720 61548 31726 61600
rect 42702 61548 42708 61600
rect 42760 61588 42766 61600
rect 52089 61591 52147 61597
rect 52089 61588 52101 61591
rect 42760 61560 52101 61588
rect 42760 61548 42766 61560
rect 52089 61557 52101 61560
rect 52135 61557 52147 61591
rect 52089 61551 52147 61557
rect 57422 61548 57428 61600
rect 57480 61588 57486 61600
rect 61930 61588 61936 61600
rect 57480 61560 61936 61588
rect 57480 61548 57486 61560
rect 61930 61548 61936 61560
rect 61988 61548 61994 61600
rect 93394 61588 93400 61600
rect 93355 61560 93400 61588
rect 93394 61548 93400 61560
rect 93452 61548 93458 61600
rect 1104 61498 98808 61520
rect 1104 61446 19606 61498
rect 19658 61446 19670 61498
rect 19722 61446 19734 61498
rect 19786 61446 19798 61498
rect 19850 61446 50326 61498
rect 50378 61446 50390 61498
rect 50442 61446 50454 61498
rect 50506 61446 50518 61498
rect 50570 61446 81046 61498
rect 81098 61446 81110 61498
rect 81162 61446 81174 61498
rect 81226 61446 81238 61498
rect 81290 61446 98808 61498
rect 1104 61424 98808 61446
rect 23106 61344 23112 61396
rect 23164 61384 23170 61396
rect 41598 61384 41604 61396
rect 23164 61356 41604 61384
rect 23164 61344 23170 61356
rect 41598 61344 41604 61356
rect 41656 61384 41662 61396
rect 42702 61384 42708 61396
rect 41656 61356 42708 61384
rect 41656 61344 41662 61356
rect 42702 61344 42708 61356
rect 42760 61344 42766 61396
rect 52914 61384 52920 61396
rect 43088 61356 52920 61384
rect 30834 61276 30840 61328
rect 30892 61316 30898 61328
rect 43088 61316 43116 61356
rect 52914 61344 52920 61356
rect 52972 61344 52978 61396
rect 73614 61384 73620 61396
rect 53024 61356 73620 61384
rect 30892 61288 43116 61316
rect 30892 61276 30898 61288
rect 44542 61276 44548 61328
rect 44600 61316 44606 61328
rect 53024 61316 53052 61356
rect 73614 61344 73620 61356
rect 73672 61344 73678 61396
rect 74810 61344 74816 61396
rect 74868 61384 74874 61396
rect 93394 61384 93400 61396
rect 74868 61356 93400 61384
rect 74868 61344 74874 61356
rect 93394 61344 93400 61356
rect 93452 61344 93458 61396
rect 82446 61316 82452 61328
rect 44600 61288 53052 61316
rect 53208 61288 57744 61316
rect 44600 61276 44606 61288
rect 9398 61208 9404 61260
rect 9456 61248 9462 61260
rect 9493 61251 9551 61257
rect 9493 61248 9505 61251
rect 9456 61220 9505 61248
rect 9456 61208 9462 61220
rect 9493 61217 9505 61220
rect 9539 61217 9551 61251
rect 9493 61211 9551 61217
rect 9769 61251 9827 61257
rect 9769 61217 9781 61251
rect 9815 61248 9827 61251
rect 10134 61248 10140 61260
rect 9815 61220 10140 61248
rect 9815 61217 9827 61220
rect 9769 61211 9827 61217
rect 9508 61180 9536 61211
rect 10134 61208 10140 61220
rect 10192 61208 10198 61260
rect 41138 61248 41144 61260
rect 41099 61220 41144 61248
rect 41138 61208 41144 61220
rect 41196 61208 41202 61260
rect 41414 61208 41420 61260
rect 41472 61248 41478 61260
rect 41690 61248 41696 61260
rect 41472 61220 41517 61248
rect 41651 61220 41696 61248
rect 41472 61208 41478 61220
rect 41690 61208 41696 61220
rect 41748 61208 41754 61260
rect 41785 61251 41843 61257
rect 41785 61217 41797 61251
rect 41831 61217 41843 61251
rect 41785 61211 41843 61217
rect 14734 61180 14740 61192
rect 9508 61152 14740 61180
rect 14734 61140 14740 61152
rect 14792 61140 14798 61192
rect 35434 61140 35440 61192
rect 35492 61180 35498 61192
rect 41800 61180 41828 61211
rect 42886 61208 42892 61260
rect 42944 61248 42950 61260
rect 52546 61248 52552 61260
rect 42944 61220 52552 61248
rect 42944 61208 42950 61220
rect 52546 61208 52552 61220
rect 52604 61208 52610 61260
rect 52914 61208 52920 61260
rect 52972 61248 52978 61260
rect 53208 61248 53236 61288
rect 52972 61220 53236 61248
rect 52972 61208 52978 61220
rect 57422 61208 57428 61260
rect 57480 61248 57486 61260
rect 57609 61251 57667 61257
rect 57609 61248 57621 61251
rect 57480 61220 57621 61248
rect 57480 61208 57486 61220
rect 57609 61217 57621 61220
rect 57655 61217 57667 61251
rect 57716 61248 57744 61288
rect 60706 61288 82452 61316
rect 60706 61248 60734 61288
rect 82446 61276 82452 61288
rect 82504 61276 82510 61328
rect 57716 61220 60734 61248
rect 57609 61211 57667 61217
rect 91922 61208 91928 61260
rect 91980 61248 91986 61260
rect 92017 61251 92075 61257
rect 92017 61248 92029 61251
rect 91980 61220 92029 61248
rect 91980 61208 91986 61220
rect 92017 61217 92029 61220
rect 92063 61217 92075 61251
rect 92017 61211 92075 61217
rect 35492 61152 41828 61180
rect 35492 61140 35498 61152
rect 41874 61140 41880 61192
rect 41932 61180 41938 61192
rect 57928 61189 57934 61192
rect 41969 61183 42027 61189
rect 41969 61180 41981 61183
rect 41932 61152 41981 61180
rect 41932 61140 41938 61152
rect 41969 61149 41981 61152
rect 42015 61149 42027 61183
rect 41969 61143 42027 61149
rect 57885 61183 57934 61189
rect 57885 61149 57897 61183
rect 57931 61149 57934 61183
rect 57885 61143 57934 61149
rect 57928 61140 57934 61143
rect 57986 61140 57992 61192
rect 92201 61183 92259 61189
rect 92201 61180 92213 61183
rect 92032 61152 92213 61180
rect 92032 61124 92060 61152
rect 92201 61149 92213 61152
rect 92247 61149 92259 61183
rect 92201 61143 92259 61149
rect 75454 61112 75460 61124
rect 58544 61084 75460 61112
rect 4157 61047 4215 61053
rect 4157 61013 4169 61047
rect 4203 61044 4215 61047
rect 4433 61047 4491 61053
rect 4433 61044 4445 61047
rect 4203 61016 4445 61044
rect 4203 61013 4215 61016
rect 4157 61007 4215 61013
rect 4433 61013 4445 61016
rect 4479 61044 4491 61047
rect 9030 61044 9036 61056
rect 4479 61016 9036 61044
rect 4479 61013 4491 61016
rect 4433 61007 4491 61013
rect 9030 61004 9036 61016
rect 9088 61004 9094 61056
rect 11057 61047 11115 61053
rect 11057 61013 11069 61047
rect 11103 61044 11115 61047
rect 58544 61044 58572 61084
rect 75454 61072 75460 61084
rect 75512 61072 75518 61124
rect 76650 61072 76656 61124
rect 76708 61112 76714 61124
rect 83734 61112 83740 61124
rect 76708 61084 83740 61112
rect 76708 61072 76714 61084
rect 83734 61072 83740 61084
rect 83792 61072 83798 61124
rect 92014 61072 92020 61124
rect 92072 61072 92078 61124
rect 58986 61044 58992 61056
rect 11103 61016 58572 61044
rect 58947 61016 58992 61044
rect 11103 61013 11115 61016
rect 11057 61007 11115 61013
rect 58986 61004 58992 61016
rect 59044 61004 59050 61056
rect 74997 61047 75055 61053
rect 74997 61013 75009 61047
rect 75043 61044 75055 61047
rect 75273 61047 75331 61053
rect 75273 61044 75285 61047
rect 75043 61016 75285 61044
rect 75043 61013 75055 61016
rect 74997 61007 75055 61013
rect 75273 61013 75285 61016
rect 75319 61044 75331 61047
rect 79318 61044 79324 61056
rect 75319 61016 79324 61044
rect 75319 61013 75331 61016
rect 75273 61007 75331 61013
rect 79318 61004 79324 61016
rect 79376 61004 79382 61056
rect 89070 61004 89076 61056
rect 89128 61044 89134 61056
rect 96985 61047 97043 61053
rect 96985 61044 96997 61047
rect 89128 61016 96997 61044
rect 89128 61004 89134 61016
rect 96985 61013 96997 61016
rect 97031 61044 97043 61047
rect 97169 61047 97227 61053
rect 97169 61044 97181 61047
rect 97031 61016 97181 61044
rect 97031 61013 97043 61016
rect 96985 61007 97043 61013
rect 97169 61013 97181 61016
rect 97215 61013 97227 61047
rect 97169 61007 97227 61013
rect 1104 60954 98808 60976
rect 1104 60902 4246 60954
rect 4298 60902 4310 60954
rect 4362 60902 4374 60954
rect 4426 60902 4438 60954
rect 4490 60902 34966 60954
rect 35018 60902 35030 60954
rect 35082 60902 35094 60954
rect 35146 60902 35158 60954
rect 35210 60902 65686 60954
rect 65738 60902 65750 60954
rect 65802 60902 65814 60954
rect 65866 60902 65878 60954
rect 65930 60902 96406 60954
rect 96458 60902 96470 60954
rect 96522 60902 96534 60954
rect 96586 60902 96598 60954
rect 96650 60902 98808 60954
rect 1104 60880 98808 60902
rect 52546 60800 52552 60852
rect 52604 60840 52610 60852
rect 58986 60840 58992 60852
rect 52604 60812 58992 60840
rect 52604 60800 52610 60812
rect 58986 60800 58992 60812
rect 59044 60800 59050 60852
rect 68094 60840 68100 60852
rect 60706 60812 67860 60840
rect 68055 60812 68100 60840
rect 7374 60732 7380 60784
rect 7432 60772 7438 60784
rect 60706 60772 60734 60812
rect 7432 60744 60734 60772
rect 67832 60772 67860 60812
rect 68094 60800 68100 60812
rect 68152 60800 68158 60852
rect 70366 60812 83596 60840
rect 70366 60772 70394 60812
rect 83568 60772 83596 60812
rect 83734 60800 83740 60852
rect 83792 60840 83798 60852
rect 89898 60840 89904 60852
rect 83792 60812 89904 60840
rect 83792 60800 83798 60812
rect 89898 60800 89904 60812
rect 89956 60840 89962 60852
rect 90818 60840 90824 60852
rect 89956 60812 90824 60840
rect 89956 60800 89962 60812
rect 90818 60800 90824 60812
rect 90876 60800 90882 60852
rect 67832 60744 70394 60772
rect 82832 60744 83504 60772
rect 83568 60744 91140 60772
rect 7432 60732 7438 60744
rect 75365 60707 75423 60713
rect 75365 60704 75377 60707
rect 57946 60676 67772 60704
rect 4985 60639 5043 60645
rect 4985 60605 4997 60639
rect 5031 60636 5043 60639
rect 5261 60639 5319 60645
rect 5261 60636 5273 60639
rect 5031 60608 5273 60636
rect 5031 60605 5043 60608
rect 4985 60599 5043 60605
rect 5261 60605 5273 60608
rect 5307 60636 5319 60639
rect 31754 60636 31760 60648
rect 5307 60608 31760 60636
rect 5307 60605 5319 60608
rect 5261 60599 5319 60605
rect 31754 60596 31760 60608
rect 31812 60596 31818 60648
rect 52730 60596 52736 60648
rect 52788 60636 52794 60648
rect 57946 60636 57974 60676
rect 67542 60636 67548 60648
rect 52788 60608 57974 60636
rect 67503 60608 67548 60636
rect 52788 60596 52794 60608
rect 67542 60596 67548 60608
rect 67600 60596 67606 60648
rect 67744 60645 67772 60676
rect 68204 60676 75377 60704
rect 67729 60639 67787 60645
rect 67729 60605 67741 60639
rect 67775 60605 67787 60639
rect 67729 60599 67787 60605
rect 67818 60596 67824 60648
rect 67876 60636 67882 60648
rect 68002 60645 68008 60648
rect 67959 60639 68008 60645
rect 67876 60608 67921 60636
rect 67876 60596 67882 60608
rect 67959 60605 67971 60639
rect 68005 60605 68008 60639
rect 67959 60599 68008 60605
rect 68002 60596 68008 60599
rect 68060 60596 68066 60648
rect 54846 60528 54852 60580
rect 54904 60568 54910 60580
rect 57054 60568 57060 60580
rect 54904 60540 57060 60568
rect 54904 60528 54910 60540
rect 57054 60528 57060 60540
rect 57112 60568 57118 60580
rect 68204 60568 68232 60676
rect 75365 60673 75377 60676
rect 75411 60673 75423 60707
rect 75365 60667 75423 60673
rect 80146 60664 80152 60716
rect 80204 60704 80210 60716
rect 82832 60704 82860 60744
rect 83476 60704 83504 60744
rect 89990 60704 89996 60716
rect 80204 60676 83044 60704
rect 83476 60676 89996 60704
rect 80204 60664 80210 60676
rect 75089 60639 75147 60645
rect 75089 60605 75101 60639
rect 75135 60636 75147 60639
rect 75914 60636 75920 60648
rect 75135 60608 75920 60636
rect 75135 60605 75147 60608
rect 75089 60599 75147 60605
rect 75914 60596 75920 60608
rect 75972 60636 75978 60648
rect 76926 60636 76932 60648
rect 75972 60608 76932 60636
rect 75972 60596 75978 60608
rect 76926 60596 76932 60608
rect 76984 60596 76990 60648
rect 83016 60645 83044 60676
rect 89990 60664 89996 60676
rect 90048 60664 90054 60716
rect 91112 60704 91140 60744
rect 91112 60676 91876 60704
rect 83001 60639 83059 60645
rect 83001 60605 83013 60639
rect 83047 60605 83059 60639
rect 83182 60636 83188 60648
rect 83143 60608 83188 60636
rect 83001 60599 83059 60605
rect 83182 60596 83188 60608
rect 83240 60596 83246 60648
rect 83366 60636 83372 60648
rect 83327 60608 83372 60636
rect 83366 60596 83372 60608
rect 83424 60596 83430 60648
rect 83642 60636 83648 60648
rect 83603 60608 83648 60636
rect 83642 60596 83648 60608
rect 83700 60596 83706 60648
rect 83737 60639 83795 60645
rect 83737 60605 83749 60639
rect 83783 60605 83795 60639
rect 83737 60599 83795 60605
rect 57112 60540 68232 60568
rect 70366 60540 74534 60568
rect 57112 60528 57118 60540
rect 29730 60460 29736 60512
rect 29788 60500 29794 60512
rect 70366 60500 70394 60540
rect 29788 60472 70394 60500
rect 74506 60500 74534 60540
rect 80882 60528 80888 60580
rect 80940 60568 80946 60580
rect 83752 60568 83780 60599
rect 84838 60596 84844 60648
rect 84896 60636 84902 60648
rect 91741 60639 91799 60645
rect 91741 60636 91753 60639
rect 84896 60608 91753 60636
rect 84896 60596 84902 60608
rect 91741 60605 91753 60608
rect 91787 60605 91799 60639
rect 91848 60636 91876 60676
rect 91922 60636 91928 60648
rect 91835 60608 91928 60636
rect 91741 60599 91799 60605
rect 91922 60596 91928 60608
rect 91980 60636 91986 60648
rect 92017 60639 92075 60645
rect 92017 60636 92029 60639
rect 91980 60608 92029 60636
rect 91980 60596 91986 60608
rect 92017 60605 92029 60608
rect 92063 60605 92075 60639
rect 92017 60599 92075 60605
rect 80940 60540 83780 60568
rect 80940 60528 80946 60540
rect 84197 60503 84255 60509
rect 84197 60500 84209 60503
rect 74506 60472 84209 60500
rect 29788 60460 29794 60472
rect 84197 60469 84209 60472
rect 84243 60469 84255 60503
rect 84197 60463 84255 60469
rect 1104 60410 98808 60432
rect 1104 60358 19606 60410
rect 19658 60358 19670 60410
rect 19722 60358 19734 60410
rect 19786 60358 19798 60410
rect 19850 60358 50326 60410
rect 50378 60358 50390 60410
rect 50442 60358 50454 60410
rect 50506 60358 50518 60410
rect 50570 60358 81046 60410
rect 81098 60358 81110 60410
rect 81162 60358 81174 60410
rect 81226 60358 81238 60410
rect 81290 60358 98808 60410
rect 1104 60336 98808 60358
rect 44266 60296 44272 60308
rect 36004 60268 44272 60296
rect 33962 60188 33968 60240
rect 34020 60228 34026 60240
rect 35894 60228 35900 60240
rect 34020 60200 35900 60228
rect 34020 60188 34026 60200
rect 35894 60188 35900 60200
rect 35952 60188 35958 60240
rect 5074 60120 5080 60172
rect 5132 60160 5138 60172
rect 5169 60163 5227 60169
rect 5169 60160 5181 60163
rect 5132 60132 5181 60160
rect 5132 60120 5138 60132
rect 5169 60129 5181 60132
rect 5215 60129 5227 60163
rect 5169 60123 5227 60129
rect 27706 60120 27712 60172
rect 27764 60160 27770 60172
rect 36004 60160 36032 60268
rect 44266 60256 44272 60268
rect 44324 60256 44330 60308
rect 54386 60256 54392 60308
rect 54444 60296 54450 60308
rect 54754 60296 54760 60308
rect 54444 60268 54760 60296
rect 54444 60256 54450 60268
rect 54754 60256 54760 60268
rect 54812 60296 54818 60308
rect 54812 60268 60734 60296
rect 54812 60256 54818 60268
rect 60706 60228 60734 60268
rect 62022 60256 62028 60308
rect 62080 60296 62086 60308
rect 68002 60296 68008 60308
rect 62080 60268 68008 60296
rect 62080 60256 62086 60268
rect 68002 60256 68008 60268
rect 68060 60256 68066 60308
rect 75730 60256 75736 60308
rect 75788 60296 75794 60308
rect 83642 60296 83648 60308
rect 75788 60268 83648 60296
rect 75788 60256 75794 60268
rect 83642 60256 83648 60268
rect 83700 60256 83706 60308
rect 67634 60228 67640 60240
rect 60706 60200 67640 60228
rect 67634 60188 67640 60200
rect 67692 60188 67698 60240
rect 72694 60188 72700 60240
rect 72752 60228 72758 60240
rect 84838 60228 84844 60240
rect 72752 60200 84844 60228
rect 72752 60188 72758 60200
rect 84838 60188 84844 60200
rect 84896 60188 84902 60240
rect 36541 60163 36599 60169
rect 36541 60160 36553 60163
rect 27764 60132 36032 60160
rect 36188 60132 36553 60160
rect 27764 60120 27770 60132
rect 5994 60092 6000 60104
rect 5955 60064 6000 60092
rect 5994 60052 6000 60064
rect 6052 60052 6058 60104
rect 34146 60052 34152 60104
rect 34204 60092 34210 60104
rect 36188 60092 36216 60132
rect 36541 60129 36553 60132
rect 36587 60129 36599 60163
rect 74810 60160 74816 60172
rect 74771 60132 74816 60160
rect 36541 60123 36599 60129
rect 74810 60120 74816 60132
rect 74868 60120 74874 60172
rect 80422 60120 80428 60172
rect 80480 60160 80486 60172
rect 83366 60160 83372 60172
rect 80480 60132 83372 60160
rect 80480 60120 80486 60132
rect 83366 60120 83372 60132
rect 83424 60120 83430 60172
rect 89809 60163 89867 60169
rect 89809 60129 89821 60163
rect 89855 60160 89867 60163
rect 89898 60160 89904 60172
rect 89855 60132 89904 60160
rect 89855 60129 89867 60132
rect 89809 60123 89867 60129
rect 89898 60120 89904 60132
rect 89956 60120 89962 60172
rect 34204 60064 36216 60092
rect 36265 60095 36323 60101
rect 34204 60052 34210 60064
rect 36265 60061 36277 60095
rect 36311 60061 36323 60095
rect 36265 60055 36323 60061
rect 34514 59984 34520 60036
rect 34572 60024 34578 60036
rect 35250 60024 35256 60036
rect 34572 59996 35256 60024
rect 34572 59984 34578 59996
rect 35250 59984 35256 59996
rect 35308 59984 35314 60036
rect 35894 59984 35900 60036
rect 35952 60024 35958 60036
rect 36280 60024 36308 60055
rect 54478 60052 54484 60104
rect 54536 60092 54542 60104
rect 56962 60092 56968 60104
rect 54536 60064 56968 60092
rect 54536 60052 54542 60064
rect 56962 60052 56968 60064
rect 57020 60092 57026 60104
rect 74997 60095 75055 60101
rect 74997 60092 75009 60095
rect 57020 60064 75009 60092
rect 57020 60052 57026 60064
rect 74997 60061 75009 60064
rect 75043 60061 75055 60095
rect 89990 60092 89996 60104
rect 89951 60064 89996 60092
rect 74997 60055 75055 60061
rect 89990 60052 89996 60064
rect 90048 60052 90054 60104
rect 72326 60024 72332 60036
rect 35952 59996 36308 60024
rect 45526 59996 72332 60024
rect 35952 59984 35958 59996
rect 33778 59916 33784 59968
rect 33836 59956 33842 59968
rect 37829 59959 37887 59965
rect 37829 59956 37841 59959
rect 33836 59928 37841 59956
rect 33836 59916 33842 59928
rect 37829 59925 37841 59928
rect 37875 59956 37887 59959
rect 45526 59956 45554 59996
rect 72326 59984 72332 59996
rect 72384 59984 72390 60036
rect 67174 59956 67180 59968
rect 37875 59928 45554 59956
rect 67135 59928 67180 59956
rect 37875 59925 37887 59928
rect 37829 59919 37887 59925
rect 67174 59916 67180 59928
rect 67232 59956 67238 59968
rect 67361 59959 67419 59965
rect 67361 59956 67373 59959
rect 67232 59928 67373 59956
rect 67232 59916 67238 59928
rect 67361 59925 67373 59928
rect 67407 59925 67419 59959
rect 67361 59919 67419 59925
rect 1104 59866 98808 59888
rect 1104 59814 4246 59866
rect 4298 59814 4310 59866
rect 4362 59814 4374 59866
rect 4426 59814 4438 59866
rect 4490 59814 34966 59866
rect 35018 59814 35030 59866
rect 35082 59814 35094 59866
rect 35146 59814 35158 59866
rect 35210 59814 65686 59866
rect 65738 59814 65750 59866
rect 65802 59814 65814 59866
rect 65866 59814 65878 59866
rect 65930 59814 96406 59866
rect 96458 59814 96470 59866
rect 96522 59814 96534 59866
rect 96586 59814 96598 59866
rect 96650 59814 98808 59866
rect 1104 59792 98808 59814
rect 29454 59712 29460 59764
rect 29512 59752 29518 59764
rect 30282 59752 30288 59764
rect 29512 59724 30288 59752
rect 29512 59712 29518 59724
rect 30282 59712 30288 59724
rect 30340 59752 30346 59764
rect 38105 59755 38163 59761
rect 38105 59752 38117 59755
rect 30340 59724 38117 59752
rect 30340 59712 30346 59724
rect 38105 59721 38117 59724
rect 38151 59721 38163 59755
rect 38105 59715 38163 59721
rect 38120 59616 38148 59715
rect 38286 59644 38292 59696
rect 38344 59684 38350 59696
rect 42981 59687 43039 59693
rect 42981 59684 42993 59687
rect 38344 59656 42993 59684
rect 38344 59644 38350 59656
rect 42981 59653 42993 59656
rect 43027 59653 43039 59687
rect 42981 59647 43039 59653
rect 64874 59644 64880 59696
rect 64932 59684 64938 59696
rect 65426 59684 65432 59696
rect 64932 59656 65432 59684
rect 64932 59644 64938 59656
rect 65426 59644 65432 59656
rect 65484 59644 65490 59696
rect 38565 59619 38623 59625
rect 6886 59588 22094 59616
rect 38120 59588 38516 59616
rect 6454 59508 6460 59560
rect 6512 59548 6518 59560
rect 6886 59548 6914 59588
rect 6512 59520 6914 59548
rect 18049 59551 18107 59557
rect 6512 59508 6518 59520
rect 18049 59517 18061 59551
rect 18095 59548 18107 59551
rect 18138 59548 18144 59560
rect 18095 59520 18144 59548
rect 18095 59517 18107 59520
rect 18049 59511 18107 59517
rect 18138 59508 18144 59520
rect 18196 59508 18202 59560
rect 22066 59480 22094 59588
rect 38286 59548 38292 59560
rect 38247 59520 38292 59548
rect 38286 59508 38292 59520
rect 38344 59508 38350 59560
rect 38488 59557 38516 59588
rect 38565 59585 38577 59619
rect 38611 59616 38623 59619
rect 54846 59616 54852 59628
rect 38611 59588 54852 59616
rect 38611 59585 38623 59588
rect 38565 59579 38623 59585
rect 38472 59551 38530 59557
rect 38472 59517 38484 59551
rect 38518 59517 38530 59551
rect 38472 59511 38530 59517
rect 38580 59480 38608 59579
rect 54846 59576 54852 59588
rect 54904 59576 54910 59628
rect 57146 59576 57152 59628
rect 57204 59616 57210 59628
rect 57790 59616 57796 59628
rect 57204 59588 57796 59616
rect 57204 59576 57210 59588
rect 57790 59576 57796 59588
rect 57848 59576 57854 59628
rect 38657 59551 38715 59557
rect 38657 59517 38669 59551
rect 38703 59517 38715 59551
rect 38838 59548 38844 59560
rect 38799 59520 38844 59548
rect 38657 59511 38715 59517
rect 22066 59452 38608 59480
rect 18233 59415 18291 59421
rect 18233 59381 18245 59415
rect 18279 59412 18291 59415
rect 18598 59412 18604 59424
rect 18279 59384 18604 59412
rect 18279 59381 18291 59384
rect 18233 59375 18291 59381
rect 18598 59372 18604 59384
rect 18656 59372 18662 59424
rect 37734 59372 37740 59424
rect 37792 59412 37798 59424
rect 38672 59412 38700 59511
rect 38838 59508 38844 59520
rect 38896 59508 38902 59560
rect 58158 59548 58164 59560
rect 39224 59520 58164 59548
rect 39022 59480 39028 59492
rect 38983 59452 39028 59480
rect 39022 59440 39028 59452
rect 39080 59440 39086 59492
rect 39224 59412 39252 59520
rect 58158 59508 58164 59520
rect 58216 59548 58222 59560
rect 58710 59548 58716 59560
rect 58216 59520 58716 59548
rect 58216 59508 58222 59520
rect 58710 59508 58716 59520
rect 58768 59508 58774 59560
rect 60737 59551 60795 59557
rect 60737 59517 60749 59551
rect 60783 59517 60795 59551
rect 60737 59511 60795 59517
rect 61013 59551 61071 59557
rect 61013 59517 61025 59551
rect 61059 59548 61071 59551
rect 64874 59548 64880 59560
rect 61059 59520 64880 59548
rect 61059 59517 61071 59520
rect 61013 59511 61071 59517
rect 42981 59483 43039 59489
rect 42981 59449 42993 59483
rect 43027 59480 43039 59483
rect 54478 59480 54484 59492
rect 43027 59452 54484 59480
rect 43027 59449 43039 59452
rect 42981 59443 43039 59449
rect 54478 59440 54484 59452
rect 54536 59440 54542 59492
rect 60752 59480 60780 59511
rect 64874 59508 64880 59520
rect 64932 59508 64938 59560
rect 60752 59452 65380 59480
rect 65352 59424 65380 59452
rect 37792 59384 39252 59412
rect 37792 59372 37798 59384
rect 55766 59372 55772 59424
rect 55824 59412 55830 59424
rect 60553 59415 60611 59421
rect 60553 59412 60565 59415
rect 55824 59384 60565 59412
rect 55824 59372 55830 59384
rect 60553 59381 60565 59384
rect 60599 59381 60611 59415
rect 60553 59375 60611 59381
rect 60921 59415 60979 59421
rect 60921 59381 60933 59415
rect 60967 59412 60979 59415
rect 63678 59412 63684 59424
rect 60967 59384 63684 59412
rect 60967 59381 60979 59384
rect 60921 59375 60979 59381
rect 63678 59372 63684 59384
rect 63736 59412 63742 59424
rect 63954 59412 63960 59424
rect 63736 59384 63960 59412
rect 63736 59372 63742 59384
rect 63954 59372 63960 59384
rect 64012 59372 64018 59424
rect 65334 59372 65340 59424
rect 65392 59412 65398 59424
rect 66070 59412 66076 59424
rect 65392 59384 66076 59412
rect 65392 59372 65398 59384
rect 66070 59372 66076 59384
rect 66128 59372 66134 59424
rect 1104 59322 98808 59344
rect 1104 59270 19606 59322
rect 19658 59270 19670 59322
rect 19722 59270 19734 59322
rect 19786 59270 19798 59322
rect 19850 59270 50326 59322
rect 50378 59270 50390 59322
rect 50442 59270 50454 59322
rect 50506 59270 50518 59322
rect 50570 59270 81046 59322
rect 81098 59270 81110 59322
rect 81162 59270 81174 59322
rect 81226 59270 81238 59322
rect 81290 59270 98808 59322
rect 1104 59248 98808 59270
rect 34790 59168 34796 59220
rect 34848 59208 34854 59220
rect 37645 59211 37703 59217
rect 37645 59208 37657 59211
rect 34848 59180 37657 59208
rect 34848 59168 34854 59180
rect 37645 59177 37657 59180
rect 37691 59177 37703 59211
rect 37645 59171 37703 59177
rect 38013 59211 38071 59217
rect 38013 59177 38025 59211
rect 38059 59208 38071 59211
rect 38059 59180 38976 59208
rect 38059 59177 38071 59180
rect 38013 59171 38071 59177
rect 15654 59100 15660 59152
rect 15712 59140 15718 59152
rect 15712 59112 38148 59140
rect 15712 59100 15718 59112
rect 20990 59032 20996 59084
rect 21048 59072 21054 59084
rect 21269 59075 21327 59081
rect 21269 59072 21281 59075
rect 21048 59044 21281 59072
rect 21048 59032 21054 59044
rect 21269 59041 21281 59044
rect 21315 59041 21327 59075
rect 37734 59072 37740 59084
rect 21269 59035 21327 59041
rect 35866 59044 37740 59072
rect 21821 59007 21879 59013
rect 21821 58973 21833 59007
rect 21867 59004 21879 59007
rect 27706 59004 27712 59016
rect 21867 58976 27712 59004
rect 21867 58973 21879 58976
rect 21821 58967 21879 58973
rect 27706 58964 27712 58976
rect 27764 59004 27770 59016
rect 28166 59004 28172 59016
rect 27764 58976 28172 59004
rect 27764 58964 27770 58976
rect 28166 58964 28172 58976
rect 28224 58964 28230 59016
rect 6546 58896 6552 58948
rect 6604 58936 6610 58948
rect 35866 58936 35894 59044
rect 37734 59032 37740 59044
rect 37792 59032 37798 59084
rect 38120 59081 38148 59112
rect 37829 59075 37887 59081
rect 37829 59041 37841 59075
rect 37875 59041 37887 59075
rect 37829 59035 37887 59041
rect 38105 59075 38163 59081
rect 38105 59041 38117 59075
rect 38151 59041 38163 59075
rect 38948 59072 38976 59180
rect 39022 59168 39028 59220
rect 39080 59208 39086 59220
rect 93213 59211 93271 59217
rect 93213 59208 93225 59211
rect 39080 59180 93225 59208
rect 39080 59168 39086 59180
rect 93213 59177 93225 59180
rect 93259 59208 93271 59211
rect 93670 59208 93676 59220
rect 93259 59180 93676 59208
rect 93259 59177 93271 59180
rect 93213 59171 93271 59177
rect 93670 59168 93676 59180
rect 93728 59168 93734 59220
rect 58894 59100 58900 59152
rect 58952 59140 58958 59152
rect 80146 59140 80152 59152
rect 58952 59112 80152 59140
rect 58952 59100 58958 59112
rect 80146 59100 80152 59112
rect 80204 59100 80210 59152
rect 43070 59072 43076 59084
rect 38948 59044 43076 59072
rect 38105 59035 38163 59041
rect 6604 58908 35894 58936
rect 37844 59004 37872 59035
rect 43070 59032 43076 59044
rect 43128 59072 43134 59084
rect 53558 59072 53564 59084
rect 43128 59044 53564 59072
rect 43128 59032 43134 59044
rect 53558 59032 53564 59044
rect 53616 59032 53622 59084
rect 76558 59032 76564 59084
rect 76616 59072 76622 59084
rect 76616 59044 93854 59072
rect 76616 59032 76622 59044
rect 37844 58976 45554 59004
rect 6604 58896 6610 58908
rect 15470 58828 15476 58880
rect 15528 58868 15534 58880
rect 37553 58871 37611 58877
rect 37553 58868 37565 58871
rect 15528 58840 37565 58868
rect 15528 58828 15534 58840
rect 37553 58837 37565 58840
rect 37599 58868 37611 58871
rect 37844 58868 37872 58976
rect 37599 58840 37872 58868
rect 45526 58868 45554 58976
rect 86862 58964 86868 59016
rect 86920 59004 86926 59016
rect 93397 59007 93455 59013
rect 93397 59004 93409 59007
rect 86920 58976 93409 59004
rect 86920 58964 86926 58976
rect 93397 58973 93409 58976
rect 93443 58973 93455 59007
rect 93670 59004 93676 59016
rect 93631 58976 93676 59004
rect 93397 58967 93455 58973
rect 93670 58964 93676 58976
rect 93728 58964 93734 59016
rect 93826 59004 93854 59044
rect 94777 59007 94835 59013
rect 94777 59004 94789 59007
rect 93826 58976 94789 59004
rect 94777 58973 94789 58976
rect 94823 58973 94835 59007
rect 94777 58967 94835 58973
rect 51442 58896 51448 58948
rect 51500 58936 51506 58948
rect 78582 58936 78588 58948
rect 51500 58908 78588 58936
rect 51500 58896 51506 58908
rect 78582 58896 78588 58908
rect 78640 58896 78646 58948
rect 83918 58868 83924 58880
rect 45526 58840 83924 58868
rect 37599 58837 37611 58840
rect 37553 58831 37611 58837
rect 83918 58828 83924 58840
rect 83976 58828 83982 58880
rect 1104 58778 98808 58800
rect 1104 58726 4246 58778
rect 4298 58726 4310 58778
rect 4362 58726 4374 58778
rect 4426 58726 4438 58778
rect 4490 58726 34966 58778
rect 35018 58726 35030 58778
rect 35082 58726 35094 58778
rect 35146 58726 35158 58778
rect 35210 58726 65686 58778
rect 65738 58726 65750 58778
rect 65802 58726 65814 58778
rect 65866 58726 65878 58778
rect 65930 58726 96406 58778
rect 96458 58726 96470 58778
rect 96522 58726 96534 58778
rect 96586 58726 96598 58778
rect 96650 58726 98808 58778
rect 1104 58704 98808 58726
rect 19334 58624 19340 58676
rect 19392 58664 19398 58676
rect 86218 58664 86224 58676
rect 19392 58636 86224 58664
rect 19392 58624 19398 58636
rect 86218 58624 86224 58636
rect 86276 58624 86282 58676
rect 57054 58488 57060 58540
rect 57112 58528 57118 58540
rect 57422 58528 57428 58540
rect 57112 58500 57428 58528
rect 57112 58488 57118 58500
rect 57422 58488 57428 58500
rect 57480 58528 57486 58540
rect 57609 58531 57667 58537
rect 57609 58528 57621 58531
rect 57480 58500 57621 58528
rect 57480 58488 57486 58500
rect 57609 58497 57621 58500
rect 57655 58497 57667 58531
rect 57609 58491 57667 58497
rect 57333 58463 57391 58469
rect 57333 58429 57345 58463
rect 57379 58460 57391 58463
rect 58158 58460 58164 58472
rect 57379 58432 58164 58460
rect 57379 58429 57391 58432
rect 57333 58423 57391 58429
rect 58158 58420 58164 58432
rect 58216 58460 58222 58472
rect 58618 58460 58624 58472
rect 58216 58432 58624 58460
rect 58216 58420 58222 58432
rect 58618 58420 58624 58432
rect 58676 58420 58682 58472
rect 81161 58463 81219 58469
rect 81161 58429 81173 58463
rect 81207 58429 81219 58463
rect 81161 58423 81219 58429
rect 81069 58327 81127 58333
rect 81069 58293 81081 58327
rect 81115 58324 81127 58327
rect 81176 58324 81204 58423
rect 81342 58324 81348 58336
rect 81115 58296 81348 58324
rect 81115 58293 81127 58296
rect 81069 58287 81127 58293
rect 81342 58284 81348 58296
rect 81400 58284 81406 58336
rect 1104 58234 98808 58256
rect 1104 58182 19606 58234
rect 19658 58182 19670 58234
rect 19722 58182 19734 58234
rect 19786 58182 19798 58234
rect 19850 58182 50326 58234
rect 50378 58182 50390 58234
rect 50442 58182 50454 58234
rect 50506 58182 50518 58234
rect 50570 58182 81046 58234
rect 81098 58182 81110 58234
rect 81162 58182 81174 58234
rect 81226 58182 81238 58234
rect 81290 58182 98808 58234
rect 1104 58160 98808 58182
rect 55858 57876 55864 57928
rect 55916 57916 55922 57928
rect 56502 57916 56508 57928
rect 55916 57888 56508 57916
rect 55916 57876 55922 57888
rect 56502 57876 56508 57888
rect 56560 57876 56566 57928
rect 53929 57783 53987 57789
rect 53929 57749 53941 57783
rect 53975 57780 53987 57783
rect 54205 57783 54263 57789
rect 54205 57780 54217 57783
rect 53975 57752 54217 57780
rect 53975 57749 53987 57752
rect 53929 57743 53987 57749
rect 54205 57749 54217 57752
rect 54251 57780 54263 57783
rect 93670 57780 93676 57792
rect 54251 57752 93676 57780
rect 54251 57749 54263 57752
rect 54205 57743 54263 57749
rect 93670 57740 93676 57752
rect 93728 57740 93734 57792
rect 1104 57690 98808 57712
rect 1104 57638 4246 57690
rect 4298 57638 4310 57690
rect 4362 57638 4374 57690
rect 4426 57638 4438 57690
rect 4490 57638 34966 57690
rect 35018 57638 35030 57690
rect 35082 57638 35094 57690
rect 35146 57638 35158 57690
rect 35210 57638 65686 57690
rect 65738 57638 65750 57690
rect 65802 57638 65814 57690
rect 65866 57638 65878 57690
rect 65930 57638 96406 57690
rect 96458 57638 96470 57690
rect 96522 57638 96534 57690
rect 96586 57638 96598 57690
rect 96650 57638 98808 57690
rect 1104 57616 98808 57638
rect 9214 57536 9220 57588
rect 9272 57576 9278 57588
rect 10321 57579 10379 57585
rect 10321 57576 10333 57579
rect 9272 57548 10333 57576
rect 9272 57536 9278 57548
rect 10321 57545 10333 57548
rect 10367 57545 10379 57579
rect 10321 57539 10379 57545
rect 18782 57468 18788 57520
rect 18840 57508 18846 57520
rect 64046 57508 64052 57520
rect 18840 57480 64052 57508
rect 18840 57468 18846 57480
rect 64046 57468 64052 57480
rect 64104 57468 64110 57520
rect 5350 57400 5356 57452
rect 5408 57440 5414 57452
rect 10413 57443 10471 57449
rect 10413 57440 10425 57443
rect 5408 57412 10425 57440
rect 5408 57400 5414 57412
rect 10413 57409 10425 57412
rect 10459 57409 10471 57443
rect 10413 57403 10471 57409
rect 22738 57400 22744 57452
rect 22796 57440 22802 57452
rect 37550 57440 37556 57452
rect 22796 57412 37556 57440
rect 22796 57400 22802 57412
rect 37550 57400 37556 57412
rect 37608 57400 37614 57452
rect 84197 57443 84255 57449
rect 84197 57409 84209 57443
rect 84243 57440 84255 57443
rect 85942 57440 85948 57452
rect 84243 57412 85948 57440
rect 84243 57409 84255 57412
rect 84197 57403 84255 57409
rect 85942 57400 85948 57412
rect 86000 57440 86006 57452
rect 86862 57440 86868 57452
rect 86000 57412 86868 57440
rect 86000 57400 86006 57412
rect 86862 57400 86868 57412
rect 86920 57400 86926 57452
rect 7190 57332 7196 57384
rect 7248 57372 7254 57384
rect 10192 57375 10250 57381
rect 10192 57372 10204 57375
rect 7248 57344 10204 57372
rect 7248 57332 7254 57344
rect 10192 57341 10204 57344
rect 10238 57341 10250 57375
rect 10192 57335 10250 57341
rect 13725 57375 13783 57381
rect 13725 57341 13737 57375
rect 13771 57372 13783 57375
rect 13998 57372 14004 57384
rect 13771 57344 14004 57372
rect 13771 57341 13783 57344
rect 13725 57335 13783 57341
rect 13998 57332 14004 57344
rect 14056 57332 14062 57384
rect 20717 57375 20775 57381
rect 20717 57341 20729 57375
rect 20763 57372 20775 57375
rect 20993 57375 21051 57381
rect 20993 57372 21005 57375
rect 20763 57344 21005 57372
rect 20763 57341 20775 57344
rect 20717 57335 20775 57341
rect 20993 57341 21005 57344
rect 21039 57372 21051 57375
rect 46934 57372 46940 57384
rect 21039 57344 46940 57372
rect 21039 57341 21051 57344
rect 20993 57335 21051 57341
rect 46934 57332 46940 57344
rect 46992 57332 46998 57384
rect 83921 57375 83979 57381
rect 83921 57372 83933 57375
rect 82924 57344 83933 57372
rect 8478 57264 8484 57316
rect 8536 57304 8542 57316
rect 10045 57307 10103 57313
rect 10045 57304 10057 57307
rect 8536 57276 10057 57304
rect 8536 57264 8542 57276
rect 10045 57273 10057 57276
rect 10091 57273 10103 57307
rect 10045 57267 10103 57273
rect 15010 57264 15016 57316
rect 15068 57304 15074 57316
rect 51902 57304 51908 57316
rect 15068 57276 51908 57304
rect 15068 57264 15074 57276
rect 51902 57264 51908 57276
rect 51960 57304 51966 57316
rect 51960 57276 55214 57304
rect 51960 57264 51966 57276
rect 10686 57236 10692 57248
rect 10647 57208 10692 57236
rect 10686 57196 10692 57208
rect 10744 57196 10750 57248
rect 55186 57236 55214 57276
rect 56502 57264 56508 57316
rect 56560 57304 56566 57316
rect 64506 57304 64512 57316
rect 56560 57276 64512 57304
rect 56560 57264 56566 57276
rect 64506 57264 64512 57276
rect 64564 57264 64570 57316
rect 82541 57307 82599 57313
rect 82541 57304 82553 57307
rect 70366 57276 82553 57304
rect 70366 57236 70394 57276
rect 82541 57273 82553 57276
rect 82587 57273 82599 57307
rect 82541 57267 82599 57273
rect 82354 57236 82360 57248
rect 55186 57208 70394 57236
rect 82315 57208 82360 57236
rect 82354 57196 82360 57208
rect 82412 57236 82418 57248
rect 82924 57236 82952 57344
rect 83921 57341 83933 57344
rect 83967 57341 83979 57375
rect 83921 57335 83979 57341
rect 85393 57375 85451 57381
rect 85393 57341 85405 57375
rect 85439 57372 85451 57375
rect 85669 57375 85727 57381
rect 85669 57372 85681 57375
rect 85439 57344 85681 57372
rect 85439 57341 85451 57344
rect 85393 57335 85451 57341
rect 85669 57341 85681 57344
rect 85715 57372 85727 57375
rect 94314 57372 94320 57384
rect 85715 57344 94320 57372
rect 85715 57341 85727 57344
rect 85669 57335 85727 57341
rect 94314 57332 94320 57344
rect 94372 57332 94378 57384
rect 82412 57208 82952 57236
rect 82412 57196 82418 57208
rect 1104 57146 98808 57168
rect 1104 57094 19606 57146
rect 19658 57094 19670 57146
rect 19722 57094 19734 57146
rect 19786 57094 19798 57146
rect 19850 57094 50326 57146
rect 50378 57094 50390 57146
rect 50442 57094 50454 57146
rect 50506 57094 50518 57146
rect 50570 57094 81046 57146
rect 81098 57094 81110 57146
rect 81162 57094 81174 57146
rect 81226 57094 81238 57146
rect 81290 57094 98808 57146
rect 1104 57072 98808 57094
rect 10686 56992 10692 57044
rect 10744 57032 10750 57044
rect 35434 57032 35440 57044
rect 10744 57004 35440 57032
rect 10744 56992 10750 57004
rect 35434 56992 35440 57004
rect 35492 56992 35498 57044
rect 59262 56992 59268 57044
rect 59320 57032 59326 57044
rect 64785 57035 64843 57041
rect 64785 57032 64797 57035
rect 59320 57004 64797 57032
rect 59320 56992 59326 57004
rect 64785 57001 64797 57004
rect 64831 57001 64843 57035
rect 64785 56995 64843 57001
rect 64046 56964 64052 56976
rect 64007 56936 64052 56964
rect 64046 56924 64052 56936
rect 64104 56964 64110 56976
rect 64506 56964 64512 56976
rect 64104 56936 64368 56964
rect 64467 56936 64512 56964
rect 64104 56924 64110 56936
rect 37458 56896 37464 56908
rect 37419 56868 37464 56896
rect 37458 56856 37464 56868
rect 37516 56856 37522 56908
rect 60642 56856 60648 56908
rect 60700 56896 60706 56908
rect 64233 56899 64291 56905
rect 64233 56896 64245 56899
rect 60700 56868 64245 56896
rect 60700 56856 60706 56868
rect 64233 56865 64245 56868
rect 64279 56865 64291 56899
rect 64340 56896 64368 56936
rect 64506 56924 64512 56936
rect 64564 56924 64570 56976
rect 94038 56924 94044 56976
rect 94096 56964 94102 56976
rect 94096 56936 97396 56964
rect 94096 56924 94102 56936
rect 64417 56899 64475 56905
rect 64417 56896 64429 56899
rect 64340 56868 64429 56896
rect 64233 56859 64291 56865
rect 64417 56865 64429 56868
rect 64463 56865 64475 56899
rect 64598 56896 64604 56908
rect 64559 56868 64604 56896
rect 64417 56859 64475 56865
rect 64598 56856 64604 56868
rect 64656 56856 64662 56908
rect 68738 56896 68744 56908
rect 68699 56868 68744 56896
rect 68738 56856 68744 56868
rect 68796 56856 68802 56908
rect 68848 56868 74534 56896
rect 38013 56831 38071 56837
rect 38013 56797 38025 56831
rect 38059 56828 38071 56831
rect 50430 56828 50436 56840
rect 38059 56800 50436 56828
rect 38059 56797 38071 56800
rect 38013 56791 38071 56797
rect 50430 56788 50436 56800
rect 50488 56788 50494 56840
rect 53742 56788 53748 56840
rect 53800 56828 53806 56840
rect 68848 56828 68876 56868
rect 53800 56800 68876 56828
rect 68925 56831 68983 56837
rect 53800 56788 53806 56800
rect 68925 56797 68937 56831
rect 68971 56797 68983 56831
rect 74506 56828 74534 56868
rect 96062 56856 96068 56908
rect 96120 56896 96126 56908
rect 96709 56899 96767 56905
rect 96709 56896 96721 56899
rect 96120 56868 96721 56896
rect 96120 56856 96126 56868
rect 96709 56865 96721 56868
rect 96755 56865 96767 56899
rect 97166 56896 97172 56908
rect 97127 56868 97172 56896
rect 96709 56859 96767 56865
rect 97166 56856 97172 56868
rect 97224 56856 97230 56908
rect 97368 56905 97396 56936
rect 97353 56899 97411 56905
rect 97353 56865 97365 56899
rect 97399 56865 97411 56899
rect 97353 56859 97411 56865
rect 97537 56899 97595 56905
rect 97537 56865 97549 56899
rect 97583 56865 97595 56899
rect 97537 56859 97595 56865
rect 97552 56828 97580 56859
rect 74506 56800 97580 56828
rect 68925 56791 68983 56797
rect 45554 56720 45560 56772
rect 45612 56760 45618 56772
rect 46842 56760 46848 56772
rect 45612 56732 46848 56760
rect 45612 56720 45618 56732
rect 46842 56720 46848 56732
rect 46900 56760 46906 56772
rect 68940 56760 68968 56791
rect 46900 56732 68968 56760
rect 46900 56720 46906 56732
rect 59265 56695 59323 56701
rect 59265 56661 59277 56695
rect 59311 56692 59323 56695
rect 59541 56695 59599 56701
rect 59541 56692 59553 56695
rect 59311 56664 59553 56692
rect 59311 56661 59323 56664
rect 59265 56655 59323 56661
rect 59541 56661 59553 56664
rect 59587 56692 59599 56695
rect 94958 56692 94964 56704
rect 59587 56664 94964 56692
rect 59587 56661 59599 56664
rect 59541 56655 59599 56661
rect 94958 56652 94964 56664
rect 95016 56652 95022 56704
rect 1104 56602 98808 56624
rect 1104 56550 4246 56602
rect 4298 56550 4310 56602
rect 4362 56550 4374 56602
rect 4426 56550 4438 56602
rect 4490 56550 34966 56602
rect 35018 56550 35030 56602
rect 35082 56550 35094 56602
rect 35146 56550 35158 56602
rect 35210 56550 65686 56602
rect 65738 56550 65750 56602
rect 65802 56550 65814 56602
rect 65866 56550 65878 56602
rect 65930 56550 96406 56602
rect 96458 56550 96470 56602
rect 96522 56550 96534 56602
rect 96586 56550 96598 56602
rect 96650 56550 98808 56602
rect 1104 56528 98808 56550
rect 31754 56448 31760 56500
rect 31812 56488 31818 56500
rect 96246 56488 96252 56500
rect 31812 56460 96252 56488
rect 31812 56448 31818 56460
rect 96246 56448 96252 56460
rect 96304 56448 96310 56500
rect 45738 56380 45744 56432
rect 45796 56420 45802 56432
rect 47578 56420 47584 56432
rect 45796 56392 47584 56420
rect 45796 56380 45802 56392
rect 47578 56380 47584 56392
rect 47636 56380 47642 56432
rect 22066 56324 35894 56352
rect 3237 56287 3295 56293
rect 3237 56253 3249 56287
rect 3283 56284 3295 56287
rect 9490 56284 9496 56296
rect 3283 56256 9496 56284
rect 3283 56253 3295 56256
rect 3237 56247 3295 56253
rect 9490 56244 9496 56256
rect 9548 56284 9554 56296
rect 10873 56287 10931 56293
rect 10873 56284 10885 56287
rect 9548 56256 10885 56284
rect 9548 56244 9554 56256
rect 10873 56253 10885 56256
rect 10919 56284 10931 56287
rect 22066 56284 22094 56324
rect 27154 56284 27160 56296
rect 10919 56256 22094 56284
rect 26528 56256 27160 56284
rect 10919 56253 10931 56256
rect 10873 56247 10931 56253
rect 3789 56219 3847 56225
rect 3789 56185 3801 56219
rect 3835 56216 3847 56219
rect 26326 56216 26332 56228
rect 3835 56188 26332 56216
rect 3835 56185 3847 56188
rect 3789 56179 3847 56185
rect 26326 56176 26332 56188
rect 26384 56216 26390 56228
rect 26528 56216 26556 56256
rect 27154 56244 27160 56256
rect 27212 56244 27218 56296
rect 33962 56284 33968 56296
rect 33923 56256 33968 56284
rect 33962 56244 33968 56256
rect 34020 56244 34026 56296
rect 34241 56287 34299 56293
rect 34241 56284 34253 56287
rect 34072 56256 34253 56284
rect 26384 56188 26556 56216
rect 26384 56176 26390 56188
rect 26602 56176 26608 56228
rect 26660 56216 26666 56228
rect 34072 56216 34100 56256
rect 34241 56253 34253 56256
rect 34287 56253 34299 56287
rect 35866 56284 35894 56324
rect 37458 56312 37464 56364
rect 37516 56352 37522 56364
rect 38102 56352 38108 56364
rect 37516 56324 38108 56352
rect 37516 56312 37522 56324
rect 38102 56312 38108 56324
rect 38160 56352 38166 56364
rect 69842 56352 69848 56364
rect 38160 56324 69848 56352
rect 38160 56312 38166 56324
rect 69842 56312 69848 56324
rect 69900 56352 69906 56364
rect 69900 56324 74534 56352
rect 69900 56312 69906 56324
rect 42245 56287 42303 56293
rect 42245 56284 42257 56287
rect 35866 56256 42257 56284
rect 34241 56247 34299 56253
rect 42245 56253 42257 56256
rect 42291 56253 42303 56287
rect 42245 56247 42303 56253
rect 49970 56244 49976 56296
rect 50028 56284 50034 56296
rect 50430 56284 50436 56296
rect 50028 56256 50436 56284
rect 50028 56244 50034 56256
rect 50430 56244 50436 56256
rect 50488 56244 50494 56296
rect 50706 56284 50712 56296
rect 50667 56256 50712 56284
rect 50706 56244 50712 56256
rect 50764 56244 50770 56296
rect 54202 56284 54208 56296
rect 54163 56256 54208 56284
rect 54202 56244 54208 56256
rect 54260 56244 54266 56296
rect 54478 56284 54484 56296
rect 54439 56256 54484 56284
rect 54478 56244 54484 56256
rect 54536 56244 54542 56296
rect 74506 56284 74534 56324
rect 82906 56284 82912 56296
rect 74506 56256 82912 56284
rect 82906 56244 82912 56256
rect 82964 56244 82970 56296
rect 41874 56216 41880 56228
rect 26660 56188 34100 56216
rect 41835 56188 41880 56216
rect 26660 56176 26666 56188
rect 41874 56176 41880 56188
rect 41932 56216 41938 56228
rect 44634 56216 44640 56228
rect 41932 56188 44640 56216
rect 41932 56176 41938 56188
rect 44634 56176 44640 56188
rect 44692 56176 44698 56228
rect 48774 56176 48780 56228
rect 48832 56216 48838 56228
rect 53374 56216 53380 56228
rect 48832 56188 53380 56216
rect 48832 56176 48838 56188
rect 53374 56176 53380 56188
rect 53432 56176 53438 56228
rect 75822 56176 75828 56228
rect 75880 56216 75886 56228
rect 92658 56216 92664 56228
rect 75880 56188 92664 56216
rect 75880 56176 75886 56188
rect 92658 56176 92664 56188
rect 92716 56176 92722 56228
rect 11057 56151 11115 56157
rect 11057 56117 11069 56151
rect 11103 56148 11115 56151
rect 11146 56148 11152 56160
rect 11103 56120 11152 56148
rect 11103 56117 11115 56120
rect 11057 56111 11115 56117
rect 11146 56108 11152 56120
rect 11204 56108 11210 56160
rect 26510 56108 26516 56160
rect 26568 56148 26574 56160
rect 26970 56148 26976 56160
rect 26568 56120 26976 56148
rect 26568 56108 26574 56120
rect 26970 56108 26976 56120
rect 27028 56148 27034 56160
rect 35345 56151 35403 56157
rect 35345 56148 35357 56151
rect 27028 56120 35357 56148
rect 27028 56108 27034 56120
rect 35345 56117 35357 56120
rect 35391 56117 35403 56151
rect 35345 56111 35403 56117
rect 47762 56108 47768 56160
rect 47820 56148 47826 56160
rect 50062 56148 50068 56160
rect 47820 56120 50068 56148
rect 47820 56108 47826 56120
rect 50062 56108 50068 56120
rect 50120 56108 50126 56160
rect 55490 56108 55496 56160
rect 55548 56148 55554 56160
rect 55769 56151 55827 56157
rect 55769 56148 55781 56151
rect 55548 56120 55781 56148
rect 55548 56108 55554 56120
rect 55769 56117 55781 56120
rect 55815 56148 55827 56151
rect 85482 56148 85488 56160
rect 55815 56120 85488 56148
rect 55815 56117 55827 56120
rect 55769 56111 55827 56117
rect 85482 56108 85488 56120
rect 85540 56108 85546 56160
rect 1104 56058 98808 56080
rect 1104 56006 19606 56058
rect 19658 56006 19670 56058
rect 19722 56006 19734 56058
rect 19786 56006 19798 56058
rect 19850 56006 50326 56058
rect 50378 56006 50390 56058
rect 50442 56006 50454 56058
rect 50506 56006 50518 56058
rect 50570 56006 81046 56058
rect 81098 56006 81110 56058
rect 81162 56006 81174 56058
rect 81226 56006 81238 56058
rect 81290 56006 98808 56058
rect 1104 55984 98808 56006
rect 11606 55904 11612 55956
rect 11664 55944 11670 55956
rect 80514 55944 80520 55956
rect 11664 55916 80520 55944
rect 11664 55904 11670 55916
rect 80514 55904 80520 55916
rect 80572 55904 80578 55956
rect 7006 55836 7012 55888
rect 7064 55876 7070 55888
rect 77478 55876 77484 55888
rect 7064 55848 77484 55876
rect 7064 55836 7070 55848
rect 77478 55836 77484 55848
rect 77536 55836 77542 55888
rect 83734 55836 83740 55888
rect 83792 55876 83798 55888
rect 85666 55876 85672 55888
rect 83792 55848 85672 55876
rect 83792 55836 83798 55848
rect 85666 55836 85672 55848
rect 85724 55836 85730 55888
rect 95050 55876 95056 55888
rect 89686 55848 95056 55876
rect 35250 55768 35256 55820
rect 35308 55808 35314 55820
rect 49053 55811 49111 55817
rect 35308 55780 49004 55808
rect 35308 55768 35314 55780
rect 11054 55632 11060 55684
rect 11112 55672 11118 55684
rect 48774 55672 48780 55684
rect 11112 55644 48780 55672
rect 11112 55632 11118 55644
rect 48774 55632 48780 55644
rect 48832 55632 48838 55684
rect 34330 55564 34336 55616
rect 34388 55604 34394 55616
rect 47762 55604 47768 55616
rect 34388 55576 47768 55604
rect 34388 55564 34394 55576
rect 47762 55564 47768 55576
rect 47820 55564 47826 55616
rect 48976 55604 49004 55780
rect 49053 55777 49065 55811
rect 49099 55777 49111 55811
rect 49053 55771 49111 55777
rect 49068 55684 49096 55771
rect 49142 55768 49148 55820
rect 49200 55817 49206 55820
rect 49510 55817 49516 55820
rect 49200 55811 49259 55817
rect 49200 55777 49213 55811
rect 49247 55777 49259 55811
rect 49200 55771 49259 55777
rect 49467 55811 49516 55817
rect 49467 55777 49479 55811
rect 49513 55777 49516 55811
rect 49467 55771 49516 55777
rect 49200 55768 49206 55771
rect 49510 55768 49516 55771
rect 49568 55768 49574 55820
rect 49605 55811 49663 55817
rect 49605 55777 49617 55811
rect 49651 55808 49663 55811
rect 49694 55808 49700 55820
rect 49651 55780 49700 55808
rect 49651 55777 49663 55780
rect 49605 55771 49663 55777
rect 49694 55768 49700 55780
rect 49752 55768 49758 55820
rect 49789 55811 49847 55817
rect 49789 55777 49801 55811
rect 49835 55808 49847 55811
rect 64046 55808 64052 55820
rect 49835 55780 64052 55808
rect 49835 55777 49847 55780
rect 49789 55771 49847 55777
rect 64046 55768 64052 55780
rect 64104 55768 64110 55820
rect 68557 55811 68615 55817
rect 68557 55777 68569 55811
rect 68603 55808 68615 55811
rect 76650 55808 76656 55820
rect 68603 55780 76656 55808
rect 68603 55777 68615 55780
rect 68557 55771 68615 55777
rect 76650 55768 76656 55780
rect 76708 55768 76714 55820
rect 49329 55743 49387 55749
rect 49329 55740 49341 55743
rect 49252 55712 49341 55740
rect 49050 55632 49056 55684
rect 49108 55632 49114 55684
rect 49252 55672 49280 55712
rect 49329 55709 49341 55712
rect 49375 55709 49387 55743
rect 59262 55740 59268 55752
rect 49329 55703 49387 55709
rect 55186 55712 59268 55740
rect 55186 55672 55214 55712
rect 59262 55700 59268 55712
rect 59320 55700 59326 55752
rect 68738 55700 68744 55752
rect 68796 55740 68802 55752
rect 68833 55743 68891 55749
rect 68833 55740 68845 55743
rect 68796 55712 68845 55740
rect 68796 55700 68802 55712
rect 68833 55709 68845 55712
rect 68879 55740 68891 55743
rect 80606 55740 80612 55752
rect 68879 55712 80612 55740
rect 68879 55709 68891 55712
rect 68833 55703 68891 55709
rect 80606 55700 80612 55712
rect 80664 55740 80670 55752
rect 89686 55740 89714 55848
rect 95050 55836 95056 55848
rect 95108 55836 95114 55888
rect 80664 55712 89714 55740
rect 80664 55700 80670 55712
rect 49252 55644 55214 55672
rect 49694 55604 49700 55616
rect 48976 55576 49700 55604
rect 49694 55564 49700 55576
rect 49752 55564 49758 55616
rect 1104 55514 98808 55536
rect 1104 55462 4246 55514
rect 4298 55462 4310 55514
rect 4362 55462 4374 55514
rect 4426 55462 4438 55514
rect 4490 55462 34966 55514
rect 35018 55462 35030 55514
rect 35082 55462 35094 55514
rect 35146 55462 35158 55514
rect 35210 55462 65686 55514
rect 65738 55462 65750 55514
rect 65802 55462 65814 55514
rect 65866 55462 65878 55514
rect 65930 55462 96406 55514
rect 96458 55462 96470 55514
rect 96522 55462 96534 55514
rect 96586 55462 96598 55514
rect 96650 55462 98808 55514
rect 1104 55440 98808 55462
rect 15102 55360 15108 55412
rect 15160 55400 15166 55412
rect 56594 55400 56600 55412
rect 15160 55372 56600 55400
rect 15160 55360 15166 55372
rect 56594 55360 56600 55372
rect 56652 55360 56658 55412
rect 42702 55292 42708 55344
rect 42760 55332 42766 55344
rect 62022 55332 62028 55344
rect 42760 55304 62028 55332
rect 42760 55292 42766 55304
rect 62022 55292 62028 55304
rect 62080 55292 62086 55344
rect 44266 55264 44272 55276
rect 44227 55236 44272 55264
rect 44266 55224 44272 55236
rect 44324 55224 44330 55276
rect 49694 55224 49700 55276
rect 49752 55264 49758 55276
rect 74810 55264 74816 55276
rect 49752 55236 74816 55264
rect 49752 55224 49758 55236
rect 74810 55224 74816 55236
rect 74868 55264 74874 55276
rect 75822 55264 75828 55276
rect 74868 55236 75828 55264
rect 74868 55224 74874 55236
rect 75822 55224 75828 55236
rect 75880 55224 75886 55276
rect 43622 55196 43628 55208
rect 43583 55168 43628 55196
rect 43622 55156 43628 55168
rect 43680 55156 43686 55208
rect 44174 55196 44180 55208
rect 44135 55168 44180 55196
rect 44174 55156 44180 55168
rect 44232 55156 44238 55208
rect 44450 55196 44456 55208
rect 44411 55168 44456 55196
rect 44450 55156 44456 55168
rect 44508 55156 44514 55208
rect 61013 55199 61071 55205
rect 61013 55196 61025 55199
rect 45526 55168 61025 55196
rect 43530 55088 43536 55140
rect 43588 55128 43594 55140
rect 45526 55128 45554 55168
rect 61013 55165 61025 55168
rect 61059 55165 61071 55199
rect 61013 55159 61071 55165
rect 84102 55156 84108 55208
rect 84160 55196 84166 55208
rect 91738 55196 91744 55208
rect 84160 55168 91744 55196
rect 84160 55156 84166 55168
rect 91738 55156 91744 55168
rect 91796 55156 91802 55208
rect 91922 55196 91928 55208
rect 91883 55168 91928 55196
rect 91922 55156 91928 55168
rect 91980 55156 91986 55208
rect 61286 55128 61292 55140
rect 43588 55100 45554 55128
rect 61247 55100 61292 55128
rect 43588 55088 43594 55100
rect 61286 55088 61292 55100
rect 61344 55088 61350 55140
rect 66346 55088 66352 55140
rect 66404 55128 66410 55140
rect 66622 55128 66628 55140
rect 66404 55100 66628 55128
rect 66404 55088 66410 55100
rect 66622 55088 66628 55100
rect 66680 55128 66686 55140
rect 92753 55131 92811 55137
rect 92753 55128 92765 55131
rect 66680 55100 92765 55128
rect 66680 55088 66686 55100
rect 92753 55097 92765 55100
rect 92799 55128 92811 55131
rect 94038 55128 94044 55140
rect 92799 55100 94044 55128
rect 92799 55097 92811 55100
rect 92753 55091 92811 55097
rect 94038 55088 94044 55100
rect 94096 55088 94102 55140
rect 14826 55020 14832 55072
rect 14884 55060 14890 55072
rect 60458 55060 60464 55072
rect 14884 55032 60464 55060
rect 14884 55020 14890 55032
rect 60458 55020 60464 55032
rect 60516 55020 60522 55072
rect 1104 54970 98808 54992
rect 1104 54918 19606 54970
rect 19658 54918 19670 54970
rect 19722 54918 19734 54970
rect 19786 54918 19798 54970
rect 19850 54918 50326 54970
rect 50378 54918 50390 54970
rect 50442 54918 50454 54970
rect 50506 54918 50518 54970
rect 50570 54918 81046 54970
rect 81098 54918 81110 54970
rect 81162 54918 81174 54970
rect 81226 54918 81238 54970
rect 81290 54918 98808 54970
rect 1104 54896 98808 54918
rect 1762 54816 1768 54868
rect 1820 54856 1826 54868
rect 44450 54856 44456 54868
rect 1820 54828 44456 54856
rect 1820 54816 1826 54828
rect 44450 54816 44456 54828
rect 44508 54816 44514 54868
rect 46934 54816 46940 54868
rect 46992 54856 46998 54868
rect 95418 54856 95424 54868
rect 46992 54828 95424 54856
rect 46992 54816 46998 54828
rect 95418 54816 95424 54828
rect 95476 54816 95482 54868
rect 84102 54788 84108 54800
rect 80026 54760 84108 54788
rect 36538 54720 36544 54732
rect 36499 54692 36544 54720
rect 36538 54680 36544 54692
rect 36596 54680 36602 54732
rect 79686 54720 79692 54732
rect 37844 54692 79692 54720
rect 33962 54612 33968 54664
rect 34020 54652 34026 54664
rect 34422 54652 34428 54664
rect 34020 54624 34428 54652
rect 34020 54612 34026 54624
rect 34422 54612 34428 54624
rect 34480 54652 34486 54664
rect 36265 54655 36323 54661
rect 36265 54652 36277 54655
rect 34480 54624 36277 54652
rect 34480 54612 34486 54624
rect 36265 54621 36277 54624
rect 36311 54621 36323 54655
rect 36265 54615 36323 54621
rect 37844 54584 37872 54692
rect 79686 54680 79692 54692
rect 79744 54680 79750 54732
rect 43438 54612 43444 54664
rect 43496 54652 43502 54664
rect 53834 54652 53840 54664
rect 43496 54624 53840 54652
rect 43496 54612 43502 54624
rect 53834 54612 53840 54624
rect 53892 54612 53898 54664
rect 58250 54612 58256 54664
rect 58308 54652 58314 54664
rect 76742 54652 76748 54664
rect 58308 54624 76748 54652
rect 58308 54612 58314 54624
rect 76742 54612 76748 54624
rect 76800 54612 76806 54664
rect 78122 54612 78128 54664
rect 78180 54652 78186 54664
rect 80026 54652 80054 54760
rect 84102 54748 84108 54760
rect 84160 54748 84166 54800
rect 83642 54720 83648 54732
rect 83555 54692 83648 54720
rect 83642 54680 83648 54692
rect 83700 54720 83706 54732
rect 88610 54720 88616 54732
rect 83700 54692 88616 54720
rect 83700 54680 83706 54692
rect 88610 54680 88616 54692
rect 88668 54680 88674 54732
rect 86129 54655 86187 54661
rect 86129 54652 86141 54655
rect 78180 54624 80054 54652
rect 84580 54624 86141 54652
rect 78180 54612 78186 54624
rect 37568 54556 37872 54584
rect 32582 54476 32588 54528
rect 32640 54516 32646 54528
rect 37568 54516 37596 54556
rect 53006 54544 53012 54596
rect 53064 54584 53070 54596
rect 78950 54584 78956 54596
rect 53064 54556 78956 54584
rect 53064 54544 53070 54556
rect 78950 54544 78956 54556
rect 79008 54544 79014 54596
rect 84580 54528 84608 54624
rect 86129 54621 86141 54624
rect 86175 54621 86187 54655
rect 86129 54615 86187 54621
rect 86405 54655 86463 54661
rect 86405 54621 86417 54655
rect 86451 54621 86463 54655
rect 86405 54615 86463 54621
rect 37826 54516 37832 54528
rect 32640 54488 37596 54516
rect 37787 54488 37832 54516
rect 32640 54476 32646 54488
rect 37826 54476 37832 54488
rect 37884 54476 37890 54528
rect 47765 54519 47823 54525
rect 47765 54485 47777 54519
rect 47811 54516 47823 54519
rect 48041 54519 48099 54525
rect 48041 54516 48053 54519
rect 47811 54488 48053 54516
rect 47811 54485 47823 54488
rect 47765 54479 47823 54485
rect 48041 54485 48053 54488
rect 48087 54516 48099 54519
rect 69934 54516 69940 54528
rect 48087 54488 69940 54516
rect 48087 54485 48099 54488
rect 48041 54479 48099 54485
rect 69934 54476 69940 54488
rect 69992 54476 69998 54528
rect 84562 54516 84568 54528
rect 84523 54488 84568 54516
rect 84562 54476 84568 54488
rect 84620 54476 84626 54528
rect 84838 54516 84844 54528
rect 84799 54488 84844 54516
rect 84838 54476 84844 54488
rect 84896 54476 84902 54528
rect 85942 54476 85948 54528
rect 86000 54516 86006 54528
rect 86420 54516 86448 54615
rect 86000 54488 86448 54516
rect 86000 54476 86006 54488
rect 1104 54426 98808 54448
rect 1104 54374 4246 54426
rect 4298 54374 4310 54426
rect 4362 54374 4374 54426
rect 4426 54374 4438 54426
rect 4490 54374 34966 54426
rect 35018 54374 35030 54426
rect 35082 54374 35094 54426
rect 35146 54374 35158 54426
rect 35210 54374 65686 54426
rect 65738 54374 65750 54426
rect 65802 54374 65814 54426
rect 65866 54374 65878 54426
rect 65930 54374 96406 54426
rect 96458 54374 96470 54426
rect 96522 54374 96534 54426
rect 96586 54374 96598 54426
rect 96650 54374 98808 54426
rect 1104 54352 98808 54374
rect 6886 54284 25452 54312
rect 1578 54136 1584 54188
rect 1636 54176 1642 54188
rect 6886 54176 6914 54284
rect 15930 54204 15936 54256
rect 15988 54244 15994 54256
rect 15988 54216 24440 54244
rect 15988 54204 15994 54216
rect 1636 54148 6914 54176
rect 1636 54136 1642 54148
rect 6178 54068 6184 54120
rect 6236 54108 6242 54120
rect 8938 54108 8944 54120
rect 6236 54080 8944 54108
rect 6236 54068 6242 54080
rect 8938 54068 8944 54080
rect 8996 54068 9002 54120
rect 24305 54111 24363 54117
rect 24305 54077 24317 54111
rect 24351 54077 24363 54111
rect 24305 54071 24363 54077
rect 24029 53975 24087 53981
rect 24029 53941 24041 53975
rect 24075 53972 24087 53975
rect 24320 53972 24348 54071
rect 24412 54040 24440 54216
rect 25424 54185 25452 54284
rect 25409 54179 25467 54185
rect 25409 54145 25421 54179
rect 25455 54145 25467 54179
rect 25409 54139 25467 54145
rect 25590 54108 25596 54120
rect 25551 54080 25596 54108
rect 25590 54068 25596 54080
rect 25648 54068 25654 54120
rect 25777 54043 25835 54049
rect 25777 54040 25789 54043
rect 24412 54012 25789 54040
rect 25777 54009 25789 54012
rect 25823 54009 25835 54043
rect 25777 54003 25835 54009
rect 44910 54000 44916 54052
rect 44968 54040 44974 54052
rect 46750 54040 46756 54052
rect 44968 54012 46756 54040
rect 44968 54000 44974 54012
rect 46750 54000 46756 54012
rect 46808 54000 46814 54052
rect 32398 53972 32404 53984
rect 24075 53944 32404 53972
rect 24075 53941 24087 53944
rect 24029 53935 24087 53941
rect 32398 53932 32404 53944
rect 32456 53932 32462 53984
rect 45186 53932 45192 53984
rect 45244 53972 45250 53984
rect 46842 53972 46848 53984
rect 45244 53944 46848 53972
rect 45244 53932 45250 53944
rect 46842 53932 46848 53944
rect 46900 53932 46906 53984
rect 1104 53882 98808 53904
rect 1104 53830 19606 53882
rect 19658 53830 19670 53882
rect 19722 53830 19734 53882
rect 19786 53830 19798 53882
rect 19850 53830 50326 53882
rect 50378 53830 50390 53882
rect 50442 53830 50454 53882
rect 50506 53830 50518 53882
rect 50570 53830 81046 53882
rect 81098 53830 81110 53882
rect 81162 53830 81174 53882
rect 81226 53830 81238 53882
rect 81290 53830 98808 53882
rect 1104 53808 98808 53830
rect 62850 53768 62856 53780
rect 21008 53740 62856 53768
rect 14734 53632 14740 53644
rect 14695 53604 14740 53632
rect 14734 53592 14740 53604
rect 14792 53592 14798 53644
rect 21008 53641 21036 53740
rect 62850 53728 62856 53740
rect 62908 53728 62914 53780
rect 23934 53700 23940 53712
rect 21100 53672 23940 53700
rect 20993 53635 21051 53641
rect 20993 53601 21005 53635
rect 21039 53601 21051 53635
rect 20993 53595 21051 53601
rect 15010 53564 15016 53576
rect 14971 53536 15016 53564
rect 15010 53524 15016 53536
rect 15068 53524 15074 53576
rect 21100 53564 21128 53672
rect 23934 53660 23940 53672
rect 23992 53700 23998 53712
rect 24210 53700 24216 53712
rect 23992 53672 24216 53700
rect 23992 53660 23998 53672
rect 24210 53660 24216 53672
rect 24268 53660 24274 53712
rect 27706 53660 27712 53712
rect 27764 53700 27770 53712
rect 28258 53700 28264 53712
rect 27764 53672 28264 53700
rect 27764 53660 27770 53672
rect 28258 53660 28264 53672
rect 28316 53660 28322 53712
rect 53374 53700 53380 53712
rect 53335 53672 53380 53700
rect 53374 53660 53380 53672
rect 53432 53700 53438 53712
rect 53745 53703 53803 53709
rect 53745 53700 53757 53703
rect 53432 53672 53757 53700
rect 53432 53660 53438 53672
rect 53745 53669 53757 53672
rect 53791 53669 53803 53703
rect 53745 53663 53803 53669
rect 53834 53660 53840 53712
rect 53892 53700 53898 53712
rect 53892 53672 53937 53700
rect 53892 53660 53898 53672
rect 58710 53660 58716 53712
rect 58768 53700 58774 53712
rect 58768 53672 70394 53700
rect 58768 53660 58774 53672
rect 21174 53592 21180 53644
rect 21232 53632 21238 53644
rect 21542 53632 21548 53644
rect 21232 53604 21276 53632
rect 21503 53604 21548 53632
rect 21232 53592 21238 53604
rect 21542 53592 21548 53604
rect 21600 53592 21606 53644
rect 54018 53641 54024 53644
rect 53561 53635 53619 53641
rect 53561 53601 53573 53635
rect 53607 53601 53619 53635
rect 53561 53595 53619 53601
rect 53981 53635 54024 53641
rect 53981 53601 53993 53635
rect 53981 53595 54024 53601
rect 21269 53567 21327 53573
rect 21269 53564 21281 53567
rect 21100 53536 21281 53564
rect 21269 53533 21281 53536
rect 21315 53533 21327 53567
rect 21269 53527 21327 53533
rect 21358 53524 21364 53576
rect 21416 53564 21422 53576
rect 21416 53536 21461 53564
rect 21416 53524 21422 53536
rect 27154 53524 27160 53576
rect 27212 53564 27218 53576
rect 53576 53564 53604 53595
rect 54018 53592 54024 53595
rect 54076 53592 54082 53644
rect 60642 53632 60648 53644
rect 55186 53604 60648 53632
rect 55186 53564 55214 53604
rect 60642 53592 60648 53604
rect 60700 53592 60706 53644
rect 63034 53592 63040 53644
rect 63092 53632 63098 53644
rect 63129 53635 63187 53641
rect 63129 53632 63141 53635
rect 63092 53604 63141 53632
rect 63092 53592 63098 53604
rect 63129 53601 63141 53604
rect 63175 53601 63187 53635
rect 63129 53595 63187 53601
rect 27212 53536 55214 53564
rect 27212 53524 27218 53536
rect 62850 53524 62856 53576
rect 62908 53564 62914 53576
rect 63497 53567 63555 53573
rect 63497 53564 63509 53567
rect 62908 53536 63509 53564
rect 62908 53524 62914 53536
rect 63497 53533 63509 53536
rect 63543 53533 63555 53567
rect 70366 53564 70394 53672
rect 75457 53635 75515 53641
rect 75457 53601 75469 53635
rect 75503 53632 75515 53635
rect 76098 53632 76104 53644
rect 75503 53604 76104 53632
rect 75503 53601 75515 53604
rect 75457 53595 75515 53601
rect 76098 53592 76104 53604
rect 76156 53632 76162 53644
rect 76156 53604 77248 53632
rect 76156 53592 76162 53604
rect 75733 53567 75791 53573
rect 75733 53564 75745 53567
rect 70366 53536 75745 53564
rect 63497 53527 63555 53533
rect 75733 53533 75745 53536
rect 75779 53533 75791 53567
rect 77220 53564 77248 53604
rect 79962 53592 79968 53644
rect 80020 53632 80026 53644
rect 84933 53635 84991 53641
rect 84933 53632 84945 53635
rect 80020 53604 84945 53632
rect 80020 53592 80026 53604
rect 84933 53601 84945 53604
rect 84979 53601 84991 53635
rect 84933 53595 84991 53601
rect 85209 53567 85267 53573
rect 85209 53564 85221 53567
rect 77220 53536 85221 53564
rect 75733 53527 75791 53533
rect 85209 53533 85221 53536
rect 85255 53533 85267 53567
rect 85209 53527 85267 53533
rect 16301 53499 16359 53505
rect 16301 53465 16313 53499
rect 16347 53496 16359 53499
rect 25682 53496 25688 53508
rect 16347 53468 25688 53496
rect 16347 53465 16359 53468
rect 16301 53459 16359 53465
rect 25682 53456 25688 53468
rect 25740 53456 25746 53508
rect 54018 53456 54024 53508
rect 54076 53496 54082 53508
rect 54297 53499 54355 53505
rect 54297 53496 54309 53499
rect 54076 53468 54309 53496
rect 54076 53456 54082 53468
rect 54297 53465 54309 53468
rect 54343 53465 54355 53499
rect 54297 53459 54355 53465
rect 21082 53388 21088 53440
rect 21140 53428 21146 53440
rect 21358 53428 21364 53440
rect 21140 53400 21364 53428
rect 21140 53388 21146 53400
rect 21358 53388 21364 53400
rect 21416 53388 21422 53440
rect 21634 53428 21640 53440
rect 21595 53400 21640 53428
rect 21634 53388 21640 53400
rect 21692 53388 21698 53440
rect 54113 53431 54171 53437
rect 54113 53397 54125 53431
rect 54159 53428 54171 53431
rect 54202 53428 54208 53440
rect 54159 53400 54208 53428
rect 54159 53397 54171 53400
rect 54113 53391 54171 53397
rect 54202 53388 54208 53400
rect 54260 53388 54266 53440
rect 54312 53428 54340 53459
rect 54386 53456 54392 53508
rect 54444 53496 54450 53508
rect 81066 53496 81072 53508
rect 54444 53468 81072 53496
rect 54444 53456 54450 53468
rect 81066 53456 81072 53468
rect 81124 53456 81130 53508
rect 61010 53428 61016 53440
rect 54312 53400 61016 53428
rect 61010 53388 61016 53400
rect 61068 53388 61074 53440
rect 1104 53338 98808 53360
rect 1104 53286 4246 53338
rect 4298 53286 4310 53338
rect 4362 53286 4374 53338
rect 4426 53286 4438 53338
rect 4490 53286 34966 53338
rect 35018 53286 35030 53338
rect 35082 53286 35094 53338
rect 35146 53286 35158 53338
rect 35210 53286 65686 53338
rect 65738 53286 65750 53338
rect 65802 53286 65814 53338
rect 65866 53286 65878 53338
rect 65930 53286 96406 53338
rect 96458 53286 96470 53338
rect 96522 53286 96534 53338
rect 96586 53286 96598 53338
rect 96650 53286 98808 53338
rect 1104 53264 98808 53286
rect 7834 53184 7840 53236
rect 7892 53224 7898 53236
rect 7892 53196 70394 53224
rect 7892 53184 7898 53196
rect 4430 53116 4436 53168
rect 4488 53156 4494 53168
rect 6178 53156 6184 53168
rect 4488 53128 6184 53156
rect 4488 53116 4494 53128
rect 6178 53116 6184 53128
rect 6236 53156 6242 53168
rect 23014 53156 23020 53168
rect 6236 53128 23020 53156
rect 6236 53116 6242 53128
rect 23014 53116 23020 53128
rect 23072 53116 23078 53168
rect 28258 53116 28264 53168
rect 28316 53156 28322 53168
rect 54018 53156 54024 53168
rect 28316 53128 54024 53156
rect 28316 53116 28322 53128
rect 54018 53116 54024 53128
rect 54076 53116 54082 53168
rect 58161 53159 58219 53165
rect 58161 53125 58173 53159
rect 58207 53156 58219 53159
rect 58250 53156 58256 53168
rect 58207 53128 58256 53156
rect 58207 53125 58219 53128
rect 58161 53119 58219 53125
rect 58250 53116 58256 53128
rect 58308 53116 58314 53168
rect 60458 53156 60464 53168
rect 60419 53128 60464 53156
rect 60458 53116 60464 53128
rect 60516 53156 60522 53168
rect 61197 53159 61255 53165
rect 60516 53128 60734 53156
rect 60516 53116 60522 53128
rect 38286 53088 38292 53100
rect 12406 53060 38292 53088
rect 5810 52912 5816 52964
rect 5868 52952 5874 52964
rect 7558 52952 7564 52964
rect 5868 52924 7564 52952
rect 5868 52912 5874 52924
rect 7558 52912 7564 52924
rect 7616 52912 7622 52964
rect 3970 52844 3976 52896
rect 4028 52884 4034 52896
rect 4982 52884 4988 52896
rect 4028 52856 4988 52884
rect 4028 52844 4034 52856
rect 4982 52844 4988 52856
rect 5040 52884 5046 52896
rect 11422 52884 11428 52896
rect 5040 52856 11428 52884
rect 5040 52844 5046 52856
rect 11422 52844 11428 52856
rect 11480 52884 11486 52896
rect 12406 52884 12434 53060
rect 38286 53048 38292 53060
rect 38344 53048 38350 53100
rect 60706 53088 60734 53128
rect 61197 53125 61209 53159
rect 61243 53156 61255 53159
rect 61378 53156 61384 53168
rect 61243 53128 61384 53156
rect 61243 53125 61255 53128
rect 61197 53119 61255 53125
rect 61378 53116 61384 53128
rect 61436 53116 61442 53168
rect 61473 53159 61531 53165
rect 61473 53125 61485 53159
rect 61519 53156 61531 53159
rect 64598 53156 64604 53168
rect 61519 53128 64604 53156
rect 61519 53125 61531 53128
rect 61473 53119 61531 53125
rect 60706 53060 60780 53088
rect 18690 52980 18696 53032
rect 18748 53020 18754 53032
rect 18785 53023 18843 53029
rect 18785 53020 18797 53023
rect 18748 52992 18797 53020
rect 18748 52980 18754 52992
rect 18785 52989 18797 52992
rect 18831 52989 18843 53023
rect 18785 52983 18843 52989
rect 46290 52980 46296 53032
rect 46348 53020 46354 53032
rect 46842 53020 46848 53032
rect 46348 52992 46848 53020
rect 46348 52980 46354 52992
rect 46842 52980 46848 52992
rect 46900 53020 46906 53032
rect 57425 53023 57483 53029
rect 57425 53020 57437 53023
rect 46900 52992 57437 53020
rect 46900 52980 46906 52992
rect 57425 52989 57437 52992
rect 57471 52989 57483 53023
rect 57425 52983 57483 52989
rect 57514 52980 57520 53032
rect 57572 53029 57578 53032
rect 57572 53023 57631 53029
rect 57572 52989 57585 53023
rect 57619 52989 57631 53023
rect 57698 53020 57704 53032
rect 57659 52992 57704 53020
rect 57572 52983 57631 52989
rect 57572 52980 57578 52983
rect 57698 52980 57704 52992
rect 57756 52980 57762 53032
rect 57793 53023 57851 53029
rect 57793 52989 57805 53023
rect 57839 52989 57851 53023
rect 57974 53020 57980 53032
rect 57935 52992 57980 53020
rect 57793 52983 57851 52989
rect 19613 52955 19671 52961
rect 19613 52921 19625 52955
rect 19659 52952 19671 52955
rect 19886 52952 19892 52964
rect 19659 52924 19892 52952
rect 19659 52921 19671 52924
rect 19613 52915 19671 52921
rect 19886 52912 19892 52924
rect 19944 52912 19950 52964
rect 46750 52912 46756 52964
rect 46808 52952 46814 52964
rect 57808 52952 57836 52983
rect 57974 52980 57980 52992
rect 58032 52980 58038 53032
rect 60642 53020 60648 53032
rect 60603 52992 60648 53020
rect 60642 52980 60648 52992
rect 60700 52980 60706 53032
rect 46808 52924 57836 52952
rect 60752 52952 60780 53060
rect 60918 53020 60924 53032
rect 60879 52992 60924 53020
rect 60918 52980 60924 52992
rect 60976 52980 60982 53032
rect 61010 52980 61016 53032
rect 61068 53029 61074 53032
rect 61068 53023 61123 53029
rect 61068 52989 61077 53023
rect 61111 53020 61123 53023
rect 61488 53020 61516 53119
rect 64598 53116 64604 53128
rect 64656 53116 64662 53168
rect 66898 53116 66904 53168
rect 66956 53156 66962 53168
rect 66993 53159 67051 53165
rect 66993 53156 67005 53159
rect 66956 53128 67005 53156
rect 66956 53116 66962 53128
rect 66993 53125 67005 53128
rect 67039 53125 67051 53159
rect 70366 53156 70394 53196
rect 71240 53196 74534 53224
rect 71130 53156 71136 53168
rect 70366 53128 71136 53156
rect 66993 53119 67051 53125
rect 71130 53116 71136 53128
rect 71188 53116 71194 53168
rect 71240 53088 71268 53196
rect 74506 53156 74534 53196
rect 85758 53156 85764 53168
rect 74506 53128 85764 53156
rect 85758 53116 85764 53128
rect 85816 53116 85822 53168
rect 66916 53060 71268 53088
rect 61111 52992 61516 53020
rect 61111 52989 61123 52992
rect 61068 52983 61123 52989
rect 61068 52980 61074 52983
rect 66070 52980 66076 53032
rect 66128 53020 66134 53032
rect 66916 53029 66944 53060
rect 71682 53048 71688 53100
rect 71740 53088 71746 53100
rect 73617 53091 73675 53097
rect 73617 53088 73629 53091
rect 71740 53060 73629 53088
rect 71740 53048 71746 53060
rect 73617 53057 73629 53060
rect 73663 53057 73675 53091
rect 81066 53088 81072 53100
rect 81027 53060 81072 53088
rect 73617 53051 73675 53057
rect 81066 53048 81072 53060
rect 81124 53048 81130 53100
rect 66901 53023 66959 53029
rect 66901 53020 66913 53023
rect 66128 52992 66913 53020
rect 66128 52980 66134 52992
rect 66901 52989 66913 52992
rect 66947 52989 66959 53023
rect 66901 52983 66959 52989
rect 66990 52980 66996 53032
rect 67048 53020 67054 53032
rect 67177 53023 67235 53029
rect 67177 53020 67189 53023
rect 67048 52992 67189 53020
rect 67048 52980 67054 52992
rect 67177 52989 67189 52992
rect 67223 52989 67235 53023
rect 73341 53023 73399 53029
rect 73341 53020 73353 53023
rect 67177 52983 67235 52989
rect 72068 52992 73353 53020
rect 60829 52955 60887 52961
rect 60829 52952 60841 52955
rect 60752 52924 60841 52952
rect 46808 52912 46814 52924
rect 60829 52921 60841 52924
rect 60875 52921 60887 52955
rect 60829 52915 60887 52921
rect 62022 52912 62028 52964
rect 62080 52952 62086 52964
rect 63678 52952 63684 52964
rect 62080 52924 63684 52952
rect 62080 52912 62086 52924
rect 63678 52912 63684 52924
rect 63736 52952 63742 52964
rect 71961 52955 72019 52961
rect 71961 52952 71973 52955
rect 63736 52924 71973 52952
rect 63736 52912 63742 52924
rect 71961 52921 71973 52924
rect 72007 52921 72019 52955
rect 71961 52915 72019 52921
rect 67358 52884 67364 52896
rect 11480 52856 12434 52884
rect 67319 52856 67364 52884
rect 11480 52844 11486 52856
rect 67358 52844 67364 52856
rect 67416 52844 67422 52896
rect 71774 52884 71780 52896
rect 71735 52856 71780 52884
rect 71774 52844 71780 52856
rect 71832 52884 71838 52896
rect 72068 52884 72096 52992
rect 73341 52989 73353 52992
rect 73387 52989 73399 53023
rect 73341 52983 73399 52989
rect 80698 52980 80704 53032
rect 80756 53020 80762 53032
rect 80793 53023 80851 53029
rect 80793 53020 80805 53023
rect 80756 52992 80805 53020
rect 80756 52980 80762 52992
rect 80793 52989 80805 52992
rect 80839 53020 80851 53023
rect 95786 53020 95792 53032
rect 80839 52992 95792 53020
rect 80839 52989 80851 52992
rect 80793 52983 80851 52989
rect 95786 52980 95792 52992
rect 95844 52980 95850 53032
rect 71832 52856 72096 52884
rect 71832 52844 71838 52856
rect 1104 52794 98808 52816
rect 1104 52742 19606 52794
rect 19658 52742 19670 52794
rect 19722 52742 19734 52794
rect 19786 52742 19798 52794
rect 19850 52742 50326 52794
rect 50378 52742 50390 52794
rect 50442 52742 50454 52794
rect 50506 52742 50518 52794
rect 50570 52742 81046 52794
rect 81098 52742 81110 52794
rect 81162 52742 81174 52794
rect 81226 52742 81238 52794
rect 81290 52742 98808 52794
rect 1104 52720 98808 52742
rect 3970 52680 3976 52692
rect 3931 52652 3976 52680
rect 3970 52640 3976 52652
rect 4028 52640 4034 52692
rect 4249 52683 4307 52689
rect 4249 52649 4261 52683
rect 4295 52680 4307 52683
rect 5074 52680 5080 52692
rect 4295 52652 5080 52680
rect 4295 52649 4307 52652
rect 4249 52643 4307 52649
rect 5074 52640 5080 52652
rect 5132 52640 5138 52692
rect 5169 52683 5227 52689
rect 5169 52649 5181 52683
rect 5215 52680 5227 52683
rect 5534 52680 5540 52692
rect 5215 52652 5540 52680
rect 5215 52649 5227 52652
rect 5169 52643 5227 52649
rect 5534 52640 5540 52652
rect 5592 52680 5598 52692
rect 6454 52680 6460 52692
rect 5592 52652 6460 52680
rect 5592 52640 5598 52652
rect 6454 52640 6460 52652
rect 6512 52640 6518 52692
rect 7377 52683 7435 52689
rect 7377 52649 7389 52683
rect 7423 52680 7435 52683
rect 7834 52680 7840 52692
rect 7423 52652 7840 52680
rect 7423 52649 7435 52652
rect 7377 52643 7435 52649
rect 7834 52640 7840 52652
rect 7892 52640 7898 52692
rect 8021 52683 8079 52689
rect 8021 52649 8033 52683
rect 8067 52680 8079 52683
rect 17862 52680 17868 52692
rect 8067 52652 17868 52680
rect 8067 52649 8079 52652
rect 8021 52643 8079 52649
rect 17862 52640 17868 52652
rect 17920 52640 17926 52692
rect 45554 52680 45560 52692
rect 36280 52652 45560 52680
rect 5810 52612 5816 52624
rect 4724 52584 5816 52612
rect 4430 52544 4436 52556
rect 4391 52516 4436 52544
rect 4430 52504 4436 52516
rect 4488 52504 4494 52556
rect 4724 52544 4752 52584
rect 5810 52572 5816 52584
rect 5868 52572 5874 52624
rect 7650 52612 7656 52624
rect 7611 52584 7656 52612
rect 7650 52572 7656 52584
rect 7708 52572 7714 52624
rect 7745 52615 7803 52621
rect 7745 52581 7757 52615
rect 7791 52612 7803 52615
rect 7791 52584 12434 52612
rect 7791 52581 7803 52584
rect 7745 52575 7803 52581
rect 4797 52547 4855 52553
rect 4797 52544 4809 52547
rect 4724 52516 4809 52544
rect 4797 52513 4809 52516
rect 4843 52513 4855 52547
rect 4982 52544 4988 52556
rect 4943 52516 4988 52544
rect 4797 52507 4855 52513
rect 4982 52504 4988 52516
rect 5040 52504 5046 52556
rect 7469 52547 7527 52553
rect 7469 52513 7481 52547
rect 7515 52513 7527 52547
rect 7834 52544 7840 52556
rect 7795 52516 7840 52544
rect 7469 52507 7527 52513
rect 4157 52479 4215 52485
rect 4157 52445 4169 52479
rect 4203 52476 4215 52479
rect 4617 52479 4675 52485
rect 4617 52476 4629 52479
rect 4203 52448 4629 52476
rect 4203 52445 4215 52448
rect 4157 52439 4215 52445
rect 4617 52445 4629 52448
rect 4663 52445 4675 52479
rect 4617 52439 4675 52445
rect 4709 52479 4767 52485
rect 4709 52445 4721 52479
rect 4755 52476 4767 52479
rect 5534 52476 5540 52488
rect 4755 52448 5540 52476
rect 4755 52445 4767 52448
rect 4709 52439 4767 52445
rect 4632 52408 4660 52439
rect 5534 52436 5540 52448
rect 5592 52436 5598 52488
rect 6546 52476 6552 52488
rect 5644 52448 6552 52476
rect 5644 52408 5672 52448
rect 6546 52436 6552 52448
rect 6604 52436 6610 52488
rect 7484 52476 7512 52507
rect 7834 52504 7840 52516
rect 7892 52504 7898 52556
rect 8110 52476 8116 52488
rect 7484 52448 8116 52476
rect 8110 52436 8116 52448
rect 8168 52436 8174 52488
rect 12406 52476 12434 52584
rect 36280 52556 36308 52652
rect 45554 52640 45560 52652
rect 45612 52640 45618 52692
rect 53650 52640 53656 52692
rect 53708 52680 53714 52692
rect 57974 52680 57980 52692
rect 53708 52652 57980 52680
rect 53708 52640 53714 52652
rect 57974 52640 57980 52652
rect 58032 52640 58038 52692
rect 67358 52640 67364 52692
rect 67416 52680 67422 52692
rect 67416 52652 80744 52680
rect 67416 52640 67422 52652
rect 42702 52612 42708 52624
rect 37016 52584 42288 52612
rect 42663 52584 42708 52612
rect 37016 52556 37044 52584
rect 36262 52544 36268 52556
rect 36175 52516 36268 52544
rect 36262 52504 36268 52516
rect 36320 52504 36326 52556
rect 36630 52544 36636 52556
rect 36591 52516 36636 52544
rect 36630 52504 36636 52516
rect 36688 52504 36694 52556
rect 36998 52544 37004 52556
rect 36911 52516 37004 52544
rect 36998 52504 37004 52516
rect 37056 52504 37062 52556
rect 37185 52547 37243 52553
rect 37185 52513 37197 52547
rect 37231 52544 37243 52547
rect 38010 52544 38016 52556
rect 37231 52516 38016 52544
rect 37231 52513 37243 52516
rect 37185 52507 37243 52513
rect 38010 52504 38016 52516
rect 38068 52504 38074 52556
rect 42150 52544 42156 52556
rect 42111 52516 42156 52544
rect 42150 52504 42156 52516
rect 42208 52504 42214 52556
rect 42260 52544 42288 52584
rect 42702 52572 42708 52584
rect 42760 52572 42766 52624
rect 57514 52572 57520 52624
rect 57572 52612 57578 52624
rect 80716 52612 80744 52652
rect 57572 52584 80376 52612
rect 80716 52584 89668 52612
rect 57572 52572 57578 52584
rect 46474 52544 46480 52556
rect 42260 52516 46480 52544
rect 46474 52504 46480 52516
rect 46532 52544 46538 52556
rect 54386 52544 54392 52556
rect 46532 52516 54392 52544
rect 46532 52504 46538 52516
rect 54386 52504 54392 52516
rect 54444 52504 54450 52556
rect 71130 52504 71136 52556
rect 71188 52544 71194 52556
rect 74442 52544 74448 52556
rect 71188 52516 74448 52544
rect 71188 52504 71194 52516
rect 74442 52504 74448 52516
rect 74500 52504 74506 52556
rect 80146 52544 80152 52556
rect 80107 52516 80152 52544
rect 80146 52504 80152 52516
rect 80204 52504 80210 52556
rect 80348 52553 80376 52584
rect 80333 52547 80391 52553
rect 80333 52513 80345 52547
rect 80379 52513 80391 52547
rect 80333 52507 80391 52513
rect 80514 52504 80520 52556
rect 80572 52544 80578 52556
rect 80882 52544 80888 52556
rect 80572 52516 80617 52544
rect 80843 52516 80888 52544
rect 80572 52504 80578 52516
rect 80882 52504 80888 52516
rect 80940 52504 80946 52556
rect 89640 52553 89668 52584
rect 89625 52547 89683 52553
rect 89625 52513 89637 52547
rect 89671 52513 89683 52547
rect 89625 52507 89683 52513
rect 33778 52476 33784 52488
rect 12406 52448 33784 52476
rect 33778 52436 33784 52448
rect 33836 52476 33842 52488
rect 33962 52476 33968 52488
rect 33836 52448 33968 52476
rect 33836 52436 33842 52448
rect 33962 52436 33968 52448
rect 34020 52436 34026 52488
rect 36446 52476 36452 52488
rect 36407 52448 36452 52476
rect 36446 52436 36452 52448
rect 36504 52436 36510 52488
rect 4632 52380 5672 52408
rect 30190 52368 30196 52420
rect 30248 52408 30254 52420
rect 36648 52408 36676 52504
rect 37366 52476 37372 52488
rect 37327 52448 37372 52476
rect 37366 52436 37372 52448
rect 37424 52436 37430 52488
rect 51718 52436 51724 52488
rect 51776 52476 51782 52488
rect 52270 52476 52276 52488
rect 51776 52448 52276 52476
rect 51776 52436 51782 52448
rect 52270 52436 52276 52448
rect 52328 52476 52334 52488
rect 80793 52479 80851 52485
rect 80793 52476 80805 52479
rect 52328 52448 80805 52476
rect 52328 52436 52334 52448
rect 80793 52445 80805 52448
rect 80839 52445 80851 52479
rect 80793 52439 80851 52445
rect 80974 52436 80980 52488
rect 81032 52476 81038 52488
rect 81253 52479 81311 52485
rect 81253 52476 81265 52479
rect 81032 52448 81265 52476
rect 81032 52436 81038 52448
rect 81253 52445 81265 52448
rect 81299 52445 81311 52479
rect 81253 52439 81311 52445
rect 82906 52436 82912 52488
rect 82964 52476 82970 52488
rect 89533 52479 89591 52485
rect 89533 52476 89545 52479
rect 82964 52448 89545 52476
rect 82964 52436 82970 52448
rect 89533 52445 89545 52448
rect 89579 52445 89591 52479
rect 89533 52439 89591 52445
rect 30248 52380 36676 52408
rect 30248 52368 30254 52380
rect 37826 52368 37832 52420
rect 37884 52408 37890 52420
rect 83274 52408 83280 52420
rect 37884 52380 83280 52408
rect 37884 52368 37890 52380
rect 83274 52368 83280 52380
rect 83332 52368 83338 52420
rect 13541 52343 13599 52349
rect 13541 52309 13553 52343
rect 13587 52340 13599 52343
rect 13817 52343 13875 52349
rect 13817 52340 13829 52343
rect 13587 52312 13829 52340
rect 13587 52309 13599 52312
rect 13541 52303 13599 52309
rect 13817 52309 13829 52312
rect 13863 52340 13875 52343
rect 39298 52340 39304 52352
rect 13863 52312 39304 52340
rect 13863 52309 13875 52312
rect 13817 52303 13875 52309
rect 39298 52300 39304 52312
rect 39356 52300 39362 52352
rect 64414 52300 64420 52352
rect 64472 52340 64478 52352
rect 67358 52340 67364 52352
rect 64472 52312 67364 52340
rect 64472 52300 64478 52312
rect 67358 52300 67364 52312
rect 67416 52300 67422 52352
rect 71038 52300 71044 52352
rect 71096 52340 71102 52352
rect 82817 52343 82875 52349
rect 82817 52340 82829 52343
rect 71096 52312 82829 52340
rect 71096 52300 71102 52312
rect 82817 52309 82829 52312
rect 82863 52340 82875 52343
rect 82909 52343 82967 52349
rect 82909 52340 82921 52343
rect 82863 52312 82921 52340
rect 82863 52309 82875 52312
rect 82817 52303 82875 52309
rect 82909 52309 82921 52312
rect 82955 52309 82967 52343
rect 82909 52303 82967 52309
rect 1104 52250 98808 52272
rect 1104 52198 4246 52250
rect 4298 52198 4310 52250
rect 4362 52198 4374 52250
rect 4426 52198 4438 52250
rect 4490 52198 34966 52250
rect 35018 52198 35030 52250
rect 35082 52198 35094 52250
rect 35146 52198 35158 52250
rect 35210 52198 65686 52250
rect 65738 52198 65750 52250
rect 65802 52198 65814 52250
rect 65866 52198 65878 52250
rect 65930 52198 96406 52250
rect 96458 52198 96470 52250
rect 96522 52198 96534 52250
rect 96586 52198 96598 52250
rect 96650 52198 98808 52250
rect 1104 52176 98808 52198
rect 54570 52096 54576 52148
rect 54628 52136 54634 52148
rect 59449 52139 59507 52145
rect 59449 52136 59461 52139
rect 54628 52108 59461 52136
rect 54628 52096 54634 52108
rect 59449 52105 59461 52108
rect 59495 52105 59507 52139
rect 59449 52099 59507 52105
rect 10594 52028 10600 52080
rect 10652 52068 10658 52080
rect 52638 52068 52644 52080
rect 10652 52040 52644 52068
rect 10652 52028 10658 52040
rect 52638 52028 52644 52040
rect 52696 52068 52702 52080
rect 58802 52068 58808 52080
rect 52696 52040 58808 52068
rect 52696 52028 52702 52040
rect 58802 52028 58808 52040
rect 58860 52028 58866 52080
rect 21358 51960 21364 52012
rect 21416 52000 21422 52012
rect 29546 52000 29552 52012
rect 21416 51972 29552 52000
rect 21416 51960 21422 51972
rect 29546 51960 29552 51972
rect 29604 51960 29610 52012
rect 9769 51935 9827 51941
rect 9769 51901 9781 51935
rect 9815 51932 9827 51935
rect 9858 51932 9864 51944
rect 9815 51904 9864 51932
rect 9815 51901 9827 51904
rect 9769 51895 9827 51901
rect 9858 51892 9864 51904
rect 9916 51892 9922 51944
rect 24210 51892 24216 51944
rect 24268 51932 24274 51944
rect 36998 51932 37004 51944
rect 24268 51904 37004 51932
rect 24268 51892 24274 51904
rect 36998 51892 37004 51904
rect 37056 51892 37062 51944
rect 41785 51935 41843 51941
rect 41785 51901 41797 51935
rect 41831 51932 41843 51935
rect 41874 51932 41880 51944
rect 41831 51904 41880 51932
rect 41831 51901 41843 51904
rect 41785 51895 41843 51901
rect 41874 51892 41880 51904
rect 41932 51892 41938 51944
rect 54570 51932 54576 51944
rect 54531 51904 54576 51932
rect 54570 51892 54576 51904
rect 54628 51892 54634 51944
rect 59262 51932 59268 51944
rect 59223 51904 59268 51932
rect 59262 51892 59268 51904
rect 59320 51932 59326 51944
rect 66346 51932 66352 51944
rect 59320 51904 66352 51932
rect 59320 51892 59326 51904
rect 66346 51892 66352 51904
rect 66404 51892 66410 51944
rect 10413 51867 10471 51873
rect 10413 51833 10425 51867
rect 10459 51864 10471 51867
rect 10594 51864 10600 51876
rect 10459 51836 10600 51864
rect 10459 51833 10471 51836
rect 10413 51827 10471 51833
rect 10594 51824 10600 51836
rect 10652 51824 10658 51876
rect 36630 51824 36636 51876
rect 36688 51864 36694 51876
rect 42061 51867 42119 51873
rect 42061 51864 42073 51867
rect 36688 51836 42073 51864
rect 36688 51824 36694 51836
rect 42061 51833 42073 51836
rect 42107 51864 42119 51867
rect 42150 51864 42156 51876
rect 42107 51836 42156 51864
rect 42107 51833 42119 51836
rect 42061 51827 42119 51833
rect 42150 51824 42156 51836
rect 42208 51824 42214 51876
rect 55122 51864 55128 51876
rect 55083 51836 55128 51864
rect 55122 51824 55128 51836
rect 55180 51824 55186 51876
rect 80514 51824 80520 51876
rect 80572 51864 80578 51876
rect 80974 51864 80980 51876
rect 80572 51836 80980 51864
rect 80572 51824 80578 51836
rect 80974 51824 80980 51836
rect 81032 51824 81038 51876
rect 12158 51756 12164 51808
rect 12216 51796 12222 51808
rect 21634 51796 21640 51808
rect 12216 51768 21640 51796
rect 12216 51756 12222 51768
rect 21634 51756 21640 51768
rect 21692 51756 21698 51808
rect 23106 51756 23112 51808
rect 23164 51796 23170 51808
rect 37826 51796 37832 51808
rect 23164 51768 37832 51796
rect 23164 51756 23170 51768
rect 37826 51756 37832 51768
rect 37884 51756 37890 51808
rect 43070 51756 43076 51808
rect 43128 51796 43134 51808
rect 62022 51796 62028 51808
rect 43128 51768 62028 51796
rect 43128 51756 43134 51768
rect 62022 51756 62028 51768
rect 62080 51756 62086 51808
rect 1104 51706 98808 51728
rect 1104 51654 19606 51706
rect 19658 51654 19670 51706
rect 19722 51654 19734 51706
rect 19786 51654 19798 51706
rect 19850 51654 50326 51706
rect 50378 51654 50390 51706
rect 50442 51654 50454 51706
rect 50506 51654 50518 51706
rect 50570 51654 81046 51706
rect 81098 51654 81110 51706
rect 81162 51654 81174 51706
rect 81226 51654 81238 51706
rect 81290 51654 98808 51706
rect 1104 51632 98808 51654
rect 83274 51552 83280 51604
rect 83332 51592 83338 51604
rect 83734 51592 83740 51604
rect 83332 51564 83740 51592
rect 83332 51552 83338 51564
rect 83734 51552 83740 51564
rect 83792 51552 83798 51604
rect 41141 51459 41199 51465
rect 41141 51425 41153 51459
rect 41187 51456 41199 51459
rect 41417 51459 41475 51465
rect 41417 51456 41429 51459
rect 41187 51428 41429 51456
rect 41187 51425 41199 51428
rect 41141 51419 41199 51425
rect 41417 51425 41429 51428
rect 41463 51425 41475 51459
rect 41417 51419 41475 51425
rect 41601 51459 41659 51465
rect 41601 51425 41613 51459
rect 41647 51425 41659 51459
rect 41601 51419 41659 51425
rect 29914 51348 29920 51400
rect 29972 51388 29978 51400
rect 41616 51388 41644 51419
rect 42061 51391 42119 51397
rect 42061 51388 42073 51391
rect 29972 51360 42073 51388
rect 29972 51348 29978 51360
rect 42061 51357 42073 51360
rect 42107 51357 42119 51391
rect 42061 51351 42119 51357
rect 39666 51212 39672 51264
rect 39724 51252 39730 51264
rect 41141 51255 41199 51261
rect 41141 51252 41153 51255
rect 39724 51224 41153 51252
rect 39724 51212 39730 51224
rect 41141 51221 41153 51224
rect 41187 51252 41199 51255
rect 41233 51255 41291 51261
rect 41233 51252 41245 51255
rect 41187 51224 41245 51252
rect 41187 51221 41199 51224
rect 41141 51215 41199 51221
rect 41233 51221 41245 51224
rect 41279 51221 41291 51255
rect 41690 51252 41696 51264
rect 41651 51224 41696 51252
rect 41233 51215 41291 51221
rect 41690 51212 41696 51224
rect 41748 51212 41754 51264
rect 61378 51212 61384 51264
rect 61436 51252 61442 51264
rect 77481 51255 77539 51261
rect 77481 51252 77493 51255
rect 61436 51224 77493 51252
rect 61436 51212 61442 51224
rect 77481 51221 77493 51224
rect 77527 51252 77539 51255
rect 77665 51255 77723 51261
rect 77665 51252 77677 51255
rect 77527 51224 77677 51252
rect 77527 51221 77539 51224
rect 77481 51215 77539 51221
rect 77665 51221 77677 51224
rect 77711 51221 77723 51255
rect 77665 51215 77723 51221
rect 1104 51162 98808 51184
rect 1104 51110 4246 51162
rect 4298 51110 4310 51162
rect 4362 51110 4374 51162
rect 4426 51110 4438 51162
rect 4490 51110 34966 51162
rect 35018 51110 35030 51162
rect 35082 51110 35094 51162
rect 35146 51110 35158 51162
rect 35210 51110 65686 51162
rect 65738 51110 65750 51162
rect 65802 51110 65814 51162
rect 65866 51110 65878 51162
rect 65930 51110 96406 51162
rect 96458 51110 96470 51162
rect 96522 51110 96534 51162
rect 96586 51110 96598 51162
rect 96650 51110 98808 51162
rect 1104 51088 98808 51110
rect 14918 51008 14924 51060
rect 14976 51048 14982 51060
rect 18966 51048 18972 51060
rect 14976 51020 18972 51048
rect 14976 51008 14982 51020
rect 18966 51008 18972 51020
rect 19024 51048 19030 51060
rect 49510 51048 49516 51060
rect 19024 51020 49516 51048
rect 19024 51008 19030 51020
rect 49510 51008 49516 51020
rect 49568 51008 49574 51060
rect 22462 50940 22468 50992
rect 22520 50980 22526 50992
rect 56042 50980 56048 50992
rect 22520 50952 56048 50980
rect 22520 50940 22526 50952
rect 56042 50940 56048 50952
rect 56100 50940 56106 50992
rect 1118 50872 1124 50924
rect 1176 50912 1182 50924
rect 48038 50912 48044 50924
rect 1176 50884 48044 50912
rect 1176 50872 1182 50884
rect 48038 50872 48044 50884
rect 48096 50872 48102 50924
rect 47578 50844 47584 50856
rect 47539 50816 47584 50844
rect 47578 50804 47584 50816
rect 47636 50804 47642 50856
rect 13446 50736 13452 50788
rect 13504 50776 13510 50788
rect 85206 50776 85212 50788
rect 13504 50748 85212 50776
rect 13504 50736 13510 50748
rect 85206 50736 85212 50748
rect 85264 50736 85270 50788
rect 8662 50668 8668 50720
rect 8720 50708 8726 50720
rect 23290 50708 23296 50720
rect 8720 50680 23296 50708
rect 8720 50668 8726 50680
rect 23290 50668 23296 50680
rect 23348 50668 23354 50720
rect 28350 50668 28356 50720
rect 28408 50708 28414 50720
rect 32950 50708 32956 50720
rect 28408 50680 32956 50708
rect 28408 50668 28414 50680
rect 32950 50668 32956 50680
rect 33008 50668 33014 50720
rect 33594 50668 33600 50720
rect 33652 50708 33658 50720
rect 34422 50708 34428 50720
rect 33652 50680 34428 50708
rect 33652 50668 33658 50680
rect 34422 50668 34428 50680
rect 34480 50708 34486 50720
rect 42334 50708 42340 50720
rect 34480 50680 42340 50708
rect 34480 50668 34486 50680
rect 42334 50668 42340 50680
rect 42392 50668 42398 50720
rect 47489 50711 47547 50717
rect 47489 50677 47501 50711
rect 47535 50708 47547 50711
rect 47578 50708 47584 50720
rect 47535 50680 47584 50708
rect 47535 50677 47547 50680
rect 47489 50671 47547 50677
rect 47578 50668 47584 50680
rect 47636 50668 47642 50720
rect 1104 50618 98808 50640
rect 1104 50566 19606 50618
rect 19658 50566 19670 50618
rect 19722 50566 19734 50618
rect 19786 50566 19798 50618
rect 19850 50566 50326 50618
rect 50378 50566 50390 50618
rect 50442 50566 50454 50618
rect 50506 50566 50518 50618
rect 50570 50566 81046 50618
rect 81098 50566 81110 50618
rect 81162 50566 81174 50618
rect 81226 50566 81238 50618
rect 81290 50566 98808 50618
rect 1104 50544 98808 50566
rect 21729 50507 21787 50513
rect 21729 50473 21741 50507
rect 21775 50504 21787 50507
rect 21913 50507 21971 50513
rect 21913 50504 21925 50507
rect 21775 50476 21925 50504
rect 21775 50473 21787 50476
rect 21729 50467 21787 50473
rect 21913 50473 21925 50476
rect 21959 50504 21971 50507
rect 60090 50504 60096 50516
rect 21959 50476 60096 50504
rect 21959 50473 21971 50476
rect 21913 50467 21971 50473
rect 60090 50464 60096 50476
rect 60148 50464 60154 50516
rect 32950 50396 32956 50448
rect 33008 50436 33014 50448
rect 48038 50436 48044 50448
rect 33008 50408 35894 50436
rect 47999 50408 48044 50436
rect 33008 50396 33014 50408
rect 18782 50328 18788 50380
rect 18840 50368 18846 50380
rect 19886 50368 19892 50380
rect 18840 50340 19892 50368
rect 18840 50328 18846 50340
rect 19886 50328 19892 50340
rect 19944 50368 19950 50380
rect 21821 50371 21879 50377
rect 21821 50368 21833 50371
rect 19944 50340 21833 50368
rect 19944 50328 19950 50340
rect 21821 50337 21833 50340
rect 21867 50337 21879 50371
rect 21821 50331 21879 50337
rect 22097 50371 22155 50377
rect 22097 50337 22109 50371
rect 22143 50368 22155 50371
rect 24486 50368 24492 50380
rect 22143 50340 24492 50368
rect 22143 50337 22155 50340
rect 22097 50331 22155 50337
rect 21836 50300 21864 50331
rect 24486 50328 24492 50340
rect 24544 50328 24550 50380
rect 27798 50328 27804 50380
rect 27856 50368 27862 50380
rect 28350 50368 28356 50380
rect 27856 50340 28356 50368
rect 27856 50328 27862 50340
rect 28350 50328 28356 50340
rect 28408 50328 28414 50380
rect 33594 50368 33600 50380
rect 31956 50340 33600 50368
rect 22462 50300 22468 50312
rect 21836 50272 22468 50300
rect 22462 50260 22468 50272
rect 22520 50260 22526 50312
rect 30374 50260 30380 50312
rect 30432 50300 30438 50312
rect 31956 50309 31984 50340
rect 33594 50328 33600 50340
rect 33652 50328 33658 50380
rect 35866 50368 35894 50408
rect 48038 50396 48044 50408
rect 48096 50396 48102 50448
rect 53374 50396 53380 50448
rect 53432 50436 53438 50448
rect 53742 50436 53748 50448
rect 53432 50408 53748 50436
rect 53432 50396 53438 50408
rect 53742 50396 53748 50408
rect 53800 50396 53806 50448
rect 63770 50396 63776 50448
rect 63828 50436 63834 50448
rect 64690 50436 64696 50448
rect 63828 50408 64696 50436
rect 63828 50396 63834 50408
rect 64690 50396 64696 50408
rect 64748 50436 64754 50448
rect 75362 50436 75368 50448
rect 64748 50408 75368 50436
rect 64748 50396 64754 50408
rect 75362 50396 75368 50408
rect 75420 50396 75426 50448
rect 90637 50439 90695 50445
rect 90637 50436 90649 50439
rect 84166 50408 90649 50436
rect 37829 50371 37887 50377
rect 35866 50340 37688 50368
rect 31941 50303 31999 50309
rect 31941 50300 31953 50303
rect 30432 50272 31953 50300
rect 30432 50260 30438 50272
rect 31941 50269 31953 50272
rect 31987 50269 31999 50303
rect 32214 50300 32220 50312
rect 32175 50272 32220 50300
rect 31941 50263 31999 50269
rect 32214 50260 32220 50272
rect 32272 50260 32278 50312
rect 8294 50192 8300 50244
rect 8352 50232 8358 50244
rect 19518 50232 19524 50244
rect 8352 50204 19524 50232
rect 8352 50192 8358 50204
rect 19518 50192 19524 50204
rect 19576 50192 19582 50244
rect 22646 50232 22652 50244
rect 19628 50204 22652 50232
rect 2038 50124 2044 50176
rect 2096 50164 2102 50176
rect 19628 50164 19656 50204
rect 22646 50192 22652 50204
rect 22704 50192 22710 50244
rect 37660 50241 37688 50340
rect 37829 50337 37841 50371
rect 37875 50368 37887 50371
rect 49605 50371 49663 50377
rect 37875 50340 45554 50368
rect 37875 50337 37887 50340
rect 37829 50331 37887 50337
rect 45526 50300 45554 50340
rect 49605 50337 49617 50371
rect 49651 50368 49663 50371
rect 58621 50371 58679 50377
rect 58621 50368 58633 50371
rect 49651 50340 58633 50368
rect 49651 50337 49663 50340
rect 49605 50331 49663 50337
rect 58621 50337 58633 50340
rect 58667 50337 58679 50371
rect 58621 50331 58679 50337
rect 72605 50371 72663 50377
rect 72605 50337 72617 50371
rect 72651 50368 72663 50371
rect 84166 50368 84194 50408
rect 90637 50405 90649 50408
rect 90683 50405 90695 50439
rect 90637 50399 90695 50405
rect 90450 50368 90456 50380
rect 72651 50340 84194 50368
rect 90411 50340 90456 50368
rect 72651 50337 72663 50340
rect 72605 50331 72663 50337
rect 49620 50300 49648 50331
rect 90450 50328 90456 50340
rect 90508 50328 90514 50380
rect 45526 50272 49648 50300
rect 65058 50260 65064 50312
rect 65116 50300 65122 50312
rect 73065 50303 73123 50309
rect 73065 50300 73077 50303
rect 65116 50272 73077 50300
rect 65116 50260 65122 50272
rect 73065 50269 73077 50272
rect 73111 50300 73123 50303
rect 75178 50300 75184 50312
rect 73111 50272 75184 50300
rect 73111 50269 73123 50272
rect 73065 50263 73123 50269
rect 75178 50260 75184 50272
rect 75236 50260 75242 50312
rect 37645 50235 37703 50241
rect 32876 50204 37596 50232
rect 22278 50164 22284 50176
rect 2096 50136 19656 50164
rect 22239 50136 22284 50164
rect 2096 50124 2102 50136
rect 22278 50124 22284 50136
rect 22336 50124 22342 50176
rect 23842 50124 23848 50176
rect 23900 50164 23906 50176
rect 32876 50164 32904 50204
rect 23900 50136 32904 50164
rect 23900 50124 23906 50136
rect 33410 50124 33416 50176
rect 33468 50164 33474 50176
rect 33505 50167 33563 50173
rect 33505 50164 33517 50167
rect 33468 50136 33517 50164
rect 33468 50124 33474 50136
rect 33505 50133 33517 50136
rect 33551 50133 33563 50167
rect 33505 50127 33563 50133
rect 36173 50167 36231 50173
rect 36173 50133 36185 50167
rect 36219 50164 36231 50167
rect 36449 50167 36507 50173
rect 36449 50164 36461 50167
rect 36219 50136 36461 50164
rect 36219 50133 36231 50136
rect 36173 50127 36231 50133
rect 36449 50133 36461 50136
rect 36495 50164 36507 50167
rect 36814 50164 36820 50176
rect 36495 50136 36820 50164
rect 36495 50133 36507 50136
rect 36449 50127 36507 50133
rect 36814 50124 36820 50136
rect 36872 50124 36878 50176
rect 37568 50164 37596 50204
rect 37645 50201 37657 50235
rect 37691 50201 37703 50235
rect 58437 50235 58495 50241
rect 37645 50195 37703 50201
rect 45526 50204 55214 50232
rect 45526 50164 45554 50204
rect 37568 50136 45554 50164
rect 55186 50164 55214 50204
rect 58437 50201 58449 50235
rect 58483 50232 58495 50235
rect 71590 50232 71596 50244
rect 58483 50204 71596 50232
rect 58483 50201 58495 50204
rect 58437 50195 58495 50201
rect 71590 50192 71596 50204
rect 71648 50192 71654 50244
rect 84562 50164 84568 50176
rect 55186 50136 84568 50164
rect 84562 50124 84568 50136
rect 84620 50124 84626 50176
rect 1104 50074 98808 50096
rect 1104 50022 4246 50074
rect 4298 50022 4310 50074
rect 4362 50022 4374 50074
rect 4426 50022 4438 50074
rect 4490 50022 34966 50074
rect 35018 50022 35030 50074
rect 35082 50022 35094 50074
rect 35146 50022 35158 50074
rect 35210 50022 65686 50074
rect 65738 50022 65750 50074
rect 65802 50022 65814 50074
rect 65866 50022 65878 50074
rect 65930 50022 96406 50074
rect 96458 50022 96470 50074
rect 96522 50022 96534 50074
rect 96586 50022 96598 50074
rect 96650 50022 98808 50074
rect 1104 50000 98808 50022
rect 13446 49960 13452 49972
rect 13407 49932 13452 49960
rect 13446 49920 13452 49932
rect 13504 49920 13510 49972
rect 17862 49920 17868 49972
rect 17920 49960 17926 49972
rect 22922 49960 22928 49972
rect 17920 49932 22928 49960
rect 17920 49920 17926 49932
rect 22922 49920 22928 49932
rect 22980 49920 22986 49972
rect 23014 49920 23020 49972
rect 23072 49960 23078 49972
rect 84838 49960 84844 49972
rect 23072 49932 84844 49960
rect 23072 49920 23078 49932
rect 84838 49920 84844 49932
rect 84896 49920 84902 49972
rect 15102 49892 15108 49904
rect 12636 49864 15108 49892
rect 1394 49756 1400 49768
rect 1355 49728 1400 49756
rect 1394 49716 1400 49728
rect 1452 49716 1458 49768
rect 12250 49756 12256 49768
rect 12211 49728 12256 49756
rect 12250 49716 12256 49728
rect 12308 49716 12314 49768
rect 12636 49765 12664 49864
rect 15102 49852 15108 49864
rect 15160 49852 15166 49904
rect 22281 49895 22339 49901
rect 22281 49861 22293 49895
rect 22327 49892 22339 49895
rect 24026 49892 24032 49904
rect 22327 49864 24032 49892
rect 22327 49861 22339 49864
rect 22281 49855 22339 49861
rect 24026 49852 24032 49864
rect 24084 49852 24090 49904
rect 49510 49852 49516 49904
rect 49568 49892 49574 49904
rect 63770 49892 63776 49904
rect 49568 49864 63776 49892
rect 49568 49852 49574 49864
rect 63770 49852 63776 49864
rect 63828 49852 63834 49904
rect 67634 49852 67640 49904
rect 67692 49892 67698 49904
rect 70121 49895 70179 49901
rect 70121 49892 70133 49895
rect 67692 49864 70133 49892
rect 67692 49852 67698 49864
rect 70121 49861 70133 49864
rect 70167 49861 70179 49895
rect 70121 49855 70179 49861
rect 12713 49827 12771 49833
rect 12713 49793 12725 49827
rect 12759 49824 12771 49827
rect 82262 49824 82268 49836
rect 12759 49796 82268 49824
rect 12759 49793 12771 49796
rect 12713 49787 12771 49793
rect 82262 49784 82268 49796
rect 82320 49784 82326 49836
rect 12621 49759 12679 49765
rect 12621 49725 12633 49759
rect 12667 49725 12679 49759
rect 12986 49756 12992 49768
rect 12947 49728 12992 49756
rect 12621 49719 12679 49725
rect 12986 49716 12992 49728
rect 13044 49716 13050 49768
rect 13173 49759 13231 49765
rect 13173 49725 13185 49759
rect 13219 49756 13231 49759
rect 17402 49756 17408 49768
rect 13219 49728 17408 49756
rect 13219 49725 13231 49728
rect 13173 49719 13231 49725
rect 17402 49716 17408 49728
rect 17460 49716 17466 49768
rect 19518 49716 19524 49768
rect 19576 49756 19582 49768
rect 22281 49759 22339 49765
rect 22281 49756 22293 49759
rect 19576 49728 22293 49756
rect 19576 49716 19582 49728
rect 22281 49725 22293 49728
rect 22327 49756 22339 49759
rect 22557 49759 22615 49765
rect 22557 49756 22569 49759
rect 22327 49728 22569 49756
rect 22327 49725 22339 49728
rect 22281 49719 22339 49725
rect 22557 49725 22569 49728
rect 22603 49725 22615 49759
rect 22557 49719 22615 49725
rect 22646 49716 22652 49768
rect 22704 49756 22710 49768
rect 22741 49759 22799 49765
rect 22741 49756 22753 49759
rect 22704 49728 22753 49756
rect 22704 49716 22710 49728
rect 22741 49725 22753 49728
rect 22787 49725 22799 49759
rect 22922 49756 22928 49768
rect 22883 49728 22928 49756
rect 22741 49719 22799 49725
rect 22922 49716 22928 49728
rect 22980 49716 22986 49768
rect 23014 49716 23020 49768
rect 23072 49756 23078 49768
rect 23201 49759 23259 49765
rect 23201 49756 23213 49759
rect 23072 49728 23213 49756
rect 23072 49716 23078 49728
rect 23201 49725 23213 49728
rect 23247 49725 23259 49759
rect 23201 49719 23259 49725
rect 23290 49716 23296 49768
rect 23348 49756 23354 49768
rect 23842 49756 23848 49768
rect 23348 49728 23393 49756
rect 23803 49728 23848 49756
rect 23348 49716 23354 49728
rect 23842 49716 23848 49728
rect 23900 49716 23906 49768
rect 30285 49759 30343 49765
rect 30285 49725 30297 49759
rect 30331 49756 30343 49759
rect 30374 49756 30380 49768
rect 30331 49728 30380 49756
rect 30331 49725 30343 49728
rect 30285 49719 30343 49725
rect 30374 49716 30380 49728
rect 30432 49716 30438 49768
rect 30558 49756 30564 49768
rect 30519 49728 30564 49756
rect 30558 49716 30564 49728
rect 30616 49716 30622 49768
rect 31754 49716 31760 49768
rect 31812 49756 31818 49768
rect 31941 49759 31999 49765
rect 31941 49756 31953 49759
rect 31812 49728 31953 49756
rect 31812 49716 31818 49728
rect 31941 49725 31953 49728
rect 31987 49725 31999 49759
rect 31941 49719 31999 49725
rect 48406 49716 48412 49768
rect 48464 49756 48470 49768
rect 48777 49759 48835 49765
rect 48777 49756 48789 49759
rect 48464 49728 48789 49756
rect 48464 49716 48470 49728
rect 48777 49725 48789 49728
rect 48823 49725 48835 49759
rect 48777 49719 48835 49725
rect 49510 49716 49516 49768
rect 49568 49756 49574 49768
rect 49605 49759 49663 49765
rect 49605 49756 49617 49759
rect 49568 49728 49617 49756
rect 49568 49716 49574 49728
rect 49605 49725 49617 49728
rect 49651 49725 49663 49759
rect 55950 49756 55956 49768
rect 55911 49728 55956 49756
rect 49605 49719 49663 49725
rect 55950 49716 55956 49728
rect 56008 49716 56014 49768
rect 71409 49759 71467 49765
rect 71409 49756 71421 49759
rect 69860 49728 71421 49756
rect 13004 49688 13032 49716
rect 43346 49688 43352 49700
rect 13004 49660 26234 49688
rect 22370 49620 22376 49632
rect 22331 49592 22376 49620
rect 22370 49580 22376 49592
rect 22428 49620 22434 49632
rect 23014 49620 23020 49632
rect 22428 49592 23020 49620
rect 22428 49580 22434 49592
rect 23014 49580 23020 49592
rect 23072 49580 23078 49632
rect 26206 49620 26234 49660
rect 31220 49660 43352 49688
rect 31220 49620 31248 49660
rect 43346 49648 43352 49660
rect 43404 49648 43410 49700
rect 48222 49648 48228 49700
rect 48280 49688 48286 49700
rect 56689 49691 56747 49697
rect 56689 49688 56701 49691
rect 48280 49660 56701 49688
rect 48280 49648 48286 49660
rect 56689 49657 56701 49660
rect 56735 49657 56747 49691
rect 56689 49651 56747 49657
rect 26206 49592 31248 49620
rect 31570 49580 31576 49632
rect 31628 49620 31634 49632
rect 69860 49629 69888 49728
rect 71409 49725 71421 49728
rect 71455 49725 71467 49759
rect 71682 49756 71688 49768
rect 71643 49728 71688 49756
rect 71409 49719 71467 49725
rect 71682 49716 71688 49728
rect 71740 49716 71746 49768
rect 69845 49623 69903 49629
rect 69845 49620 69857 49623
rect 31628 49592 69857 49620
rect 31628 49580 31634 49592
rect 69845 49589 69857 49592
rect 69891 49589 69903 49623
rect 69845 49583 69903 49589
rect 1104 49530 98808 49552
rect 1104 49478 19606 49530
rect 19658 49478 19670 49530
rect 19722 49478 19734 49530
rect 19786 49478 19798 49530
rect 19850 49478 50326 49530
rect 50378 49478 50390 49530
rect 50442 49478 50454 49530
rect 50506 49478 50518 49530
rect 50570 49478 81046 49530
rect 81098 49478 81110 49530
rect 81162 49478 81174 49530
rect 81226 49478 81238 49530
rect 81290 49478 98808 49530
rect 1104 49456 98808 49478
rect 24026 49376 24032 49428
rect 24084 49416 24090 49428
rect 69658 49416 69664 49428
rect 24084 49388 69664 49416
rect 24084 49376 24090 49388
rect 69658 49376 69664 49388
rect 69716 49376 69722 49428
rect 70118 49376 70124 49428
rect 70176 49416 70182 49428
rect 82722 49416 82728 49428
rect 70176 49388 82728 49416
rect 70176 49376 70182 49388
rect 82722 49376 82728 49388
rect 82780 49376 82786 49428
rect 28442 49308 28448 49360
rect 28500 49348 28506 49360
rect 31570 49348 31576 49360
rect 28500 49320 31576 49348
rect 28500 49308 28506 49320
rect 31570 49308 31576 49320
rect 31628 49308 31634 49360
rect 69676 49348 69704 49376
rect 81986 49348 81992 49360
rect 69676 49320 81992 49348
rect 81986 49308 81992 49320
rect 82044 49348 82050 49360
rect 82044 49320 84194 49348
rect 82044 49308 82050 49320
rect 15010 49240 15016 49292
rect 15068 49280 15074 49292
rect 76190 49280 76196 49292
rect 15068 49252 76196 49280
rect 15068 49240 15074 49252
rect 76190 49240 76196 49252
rect 76248 49240 76254 49292
rect 84166 49280 84194 49320
rect 92842 49280 92848 49292
rect 84166 49252 92848 49280
rect 92842 49240 92848 49252
rect 92900 49240 92906 49292
rect 36722 49172 36728 49224
rect 36780 49212 36786 49224
rect 38194 49212 38200 49224
rect 36780 49184 38200 49212
rect 36780 49172 36786 49184
rect 38194 49172 38200 49184
rect 38252 49172 38258 49224
rect 42334 49212 42340 49224
rect 42295 49184 42340 49212
rect 42334 49172 42340 49184
rect 42392 49172 42398 49224
rect 42613 49215 42671 49221
rect 42613 49181 42625 49215
rect 42659 49212 42671 49215
rect 46198 49212 46204 49224
rect 42659 49184 46204 49212
rect 42659 49181 42671 49184
rect 42613 49175 42671 49181
rect 46198 49172 46204 49184
rect 46256 49172 46262 49224
rect 58802 49172 58808 49224
rect 58860 49212 58866 49224
rect 78030 49212 78036 49224
rect 58860 49184 78036 49212
rect 58860 49172 58866 49184
rect 78030 49172 78036 49184
rect 78088 49172 78094 49224
rect 84194 49172 84200 49224
rect 84252 49212 84258 49224
rect 85669 49215 85727 49221
rect 85669 49212 85681 49215
rect 84252 49184 85681 49212
rect 84252 49172 84258 49184
rect 85669 49181 85681 49184
rect 85715 49181 85727 49215
rect 85942 49212 85948 49224
rect 85903 49184 85948 49212
rect 85669 49175 85727 49181
rect 85942 49172 85948 49184
rect 86000 49172 86006 49224
rect 3694 49104 3700 49156
rect 3752 49144 3758 49156
rect 12986 49144 12992 49156
rect 3752 49116 12992 49144
rect 3752 49104 3758 49116
rect 12986 49104 12992 49116
rect 13044 49104 13050 49156
rect 19242 49104 19248 49156
rect 19300 49144 19306 49156
rect 25866 49144 25872 49156
rect 19300 49116 25872 49144
rect 19300 49104 19306 49116
rect 25866 49104 25872 49116
rect 25924 49144 25930 49156
rect 36078 49144 36084 49156
rect 25924 49116 36084 49144
rect 25924 49104 25930 49116
rect 36078 49104 36084 49116
rect 36136 49104 36142 49156
rect 43346 49104 43352 49156
rect 43404 49144 43410 49156
rect 47026 49144 47032 49156
rect 43404 49116 47032 49144
rect 43404 49104 43410 49116
rect 47026 49104 47032 49116
rect 47084 49144 47090 49156
rect 48222 49144 48228 49156
rect 47084 49116 48228 49144
rect 47084 49104 47090 49116
rect 48222 49104 48228 49116
rect 48280 49104 48286 49156
rect 53742 49104 53748 49156
rect 53800 49144 53806 49156
rect 55398 49144 55404 49156
rect 53800 49116 55404 49144
rect 53800 49104 53806 49116
rect 55398 49104 55404 49116
rect 55456 49144 55462 49156
rect 84381 49147 84439 49153
rect 84381 49144 84393 49147
rect 55456 49116 84393 49144
rect 55456 49104 55462 49116
rect 84381 49113 84393 49116
rect 84427 49113 84439 49147
rect 84381 49107 84439 49113
rect 1489 49079 1547 49085
rect 1489 49045 1501 49079
rect 1535 49076 1547 49079
rect 1765 49079 1823 49085
rect 1765 49076 1777 49079
rect 1535 49048 1777 49076
rect 1535 49045 1547 49048
rect 1489 49039 1547 49045
rect 1765 49045 1777 49048
rect 1811 49076 1823 49079
rect 16114 49076 16120 49088
rect 1811 49048 16120 49076
rect 1811 49045 1823 49048
rect 1765 49039 1823 49045
rect 16114 49036 16120 49048
rect 16172 49036 16178 49088
rect 22373 49079 22431 49085
rect 22373 49045 22385 49079
rect 22419 49076 22431 49079
rect 22646 49076 22652 49088
rect 22419 49048 22652 49076
rect 22419 49045 22431 49048
rect 22373 49039 22431 49045
rect 22646 49036 22652 49048
rect 22704 49036 22710 49088
rect 24029 49079 24087 49085
rect 24029 49045 24041 49079
rect 24075 49076 24087 49079
rect 24302 49076 24308 49088
rect 24075 49048 24308 49076
rect 24075 49045 24087 49048
rect 24029 49039 24087 49045
rect 24302 49036 24308 49048
rect 24360 49036 24366 49088
rect 43714 49076 43720 49088
rect 43675 49048 43720 49076
rect 43714 49036 43720 49048
rect 43772 49036 43778 49088
rect 1104 48986 98808 49008
rect 1104 48934 4246 48986
rect 4298 48934 4310 48986
rect 4362 48934 4374 48986
rect 4426 48934 4438 48986
rect 4490 48934 34966 48986
rect 35018 48934 35030 48986
rect 35082 48934 35094 48986
rect 35146 48934 35158 48986
rect 35210 48934 65686 48986
rect 65738 48934 65750 48986
rect 65802 48934 65814 48986
rect 65866 48934 65878 48986
rect 65930 48934 96406 48986
rect 96458 48934 96470 48986
rect 96522 48934 96534 48986
rect 96586 48934 96598 48986
rect 96650 48934 98808 48986
rect 1104 48912 98808 48934
rect 24302 48832 24308 48884
rect 24360 48872 24366 48884
rect 30098 48872 30104 48884
rect 24360 48844 30104 48872
rect 24360 48832 24366 48844
rect 30098 48832 30104 48844
rect 30156 48832 30162 48884
rect 48958 48832 48964 48884
rect 49016 48872 49022 48884
rect 84194 48872 84200 48884
rect 49016 48844 84200 48872
rect 49016 48832 49022 48844
rect 84194 48832 84200 48844
rect 84252 48832 84258 48884
rect 18598 48764 18604 48816
rect 18656 48804 18662 48816
rect 18656 48776 21036 48804
rect 18656 48764 18662 48776
rect 15378 48696 15384 48748
rect 15436 48736 15442 48748
rect 18877 48739 18935 48745
rect 18877 48736 18889 48739
rect 15436 48708 18889 48736
rect 15436 48696 15442 48708
rect 18877 48705 18889 48708
rect 18923 48736 18935 48739
rect 21008 48736 21036 48776
rect 22646 48764 22652 48816
rect 22704 48804 22710 48816
rect 87506 48804 87512 48816
rect 22704 48776 87512 48804
rect 22704 48764 22710 48776
rect 87506 48764 87512 48776
rect 87564 48764 87570 48816
rect 18923 48708 19380 48736
rect 21008 48708 34284 48736
rect 18923 48705 18935 48708
rect 18877 48699 18935 48705
rect 18966 48668 18972 48680
rect 18927 48640 18972 48668
rect 18966 48628 18972 48640
rect 19024 48628 19030 48680
rect 19242 48668 19248 48680
rect 19203 48640 19248 48668
rect 19242 48628 19248 48640
rect 19300 48628 19306 48680
rect 19352 48677 19380 48708
rect 34256 48677 34284 48708
rect 67542 48696 67548 48748
rect 67600 48736 67606 48748
rect 68005 48739 68063 48745
rect 68005 48736 68017 48739
rect 67600 48708 68017 48736
rect 67600 48696 67606 48708
rect 68005 48705 68017 48708
rect 68051 48705 68063 48739
rect 68005 48699 68063 48705
rect 19337 48671 19395 48677
rect 19337 48637 19349 48671
rect 19383 48668 19395 48671
rect 34241 48671 34299 48677
rect 19383 48640 26234 48668
rect 19383 48637 19395 48640
rect 19337 48631 19395 48637
rect 19153 48603 19211 48609
rect 19153 48569 19165 48603
rect 19199 48569 19211 48603
rect 22830 48600 22836 48612
rect 19153 48563 19211 48569
rect 19352 48572 22836 48600
rect 19168 48532 19196 48563
rect 19352 48532 19380 48572
rect 22830 48560 22836 48572
rect 22888 48560 22894 48612
rect 23934 48560 23940 48612
rect 23992 48600 23998 48612
rect 24210 48600 24216 48612
rect 23992 48572 24216 48600
rect 23992 48560 23998 48572
rect 24210 48560 24216 48572
rect 24268 48560 24274 48612
rect 26206 48600 26234 48640
rect 34241 48637 34253 48671
rect 34287 48637 34299 48671
rect 65058 48668 65064 48680
rect 34241 48631 34299 48637
rect 34348 48640 65064 48668
rect 34348 48600 34376 48640
rect 65058 48628 65064 48640
rect 65116 48628 65122 48680
rect 67726 48668 67732 48680
rect 67687 48640 67732 48668
rect 67726 48628 67732 48640
rect 67784 48628 67790 48680
rect 26206 48572 34376 48600
rect 35069 48603 35127 48609
rect 35069 48569 35081 48603
rect 35115 48600 35127 48603
rect 52454 48600 52460 48612
rect 35115 48572 52460 48600
rect 35115 48569 35127 48572
rect 35069 48563 35127 48569
rect 52454 48560 52460 48572
rect 52512 48560 52518 48612
rect 19168 48504 19380 48532
rect 19521 48535 19579 48541
rect 19521 48501 19533 48535
rect 19567 48532 19579 48535
rect 20530 48532 20536 48544
rect 19567 48504 20536 48532
rect 19567 48501 19579 48504
rect 19521 48495 19579 48501
rect 20530 48492 20536 48504
rect 20588 48492 20594 48544
rect 1104 48442 98808 48464
rect 1104 48390 19606 48442
rect 19658 48390 19670 48442
rect 19722 48390 19734 48442
rect 19786 48390 19798 48442
rect 19850 48390 50326 48442
rect 50378 48390 50390 48442
rect 50442 48390 50454 48442
rect 50506 48390 50518 48442
rect 50570 48390 81046 48442
rect 81098 48390 81110 48442
rect 81162 48390 81174 48442
rect 81226 48390 81238 48442
rect 81290 48390 98808 48442
rect 1104 48368 98808 48390
rect 45278 48328 45284 48340
rect 42720 48300 45284 48328
rect 34054 48260 34060 48272
rect 5276 48232 34060 48260
rect 4890 48192 4896 48204
rect 4851 48164 4896 48192
rect 4890 48152 4896 48164
rect 4948 48152 4954 48204
rect 5276 48201 5304 48232
rect 34054 48220 34060 48232
rect 34112 48220 34118 48272
rect 5261 48195 5319 48201
rect 5261 48161 5273 48195
rect 5307 48161 5319 48195
rect 5261 48155 5319 48161
rect 5445 48195 5503 48201
rect 5445 48161 5457 48195
rect 5491 48161 5503 48195
rect 41785 48195 41843 48201
rect 5445 48155 5503 48161
rect 8312 48164 12434 48192
rect 4985 48127 5043 48133
rect 4985 48093 4997 48127
rect 5031 48093 5043 48127
rect 5460 48124 5488 48155
rect 8312 48124 8340 48164
rect 5460 48096 8340 48124
rect 12406 48124 12434 48164
rect 41785 48161 41797 48195
rect 41831 48192 41843 48195
rect 42334 48192 42340 48204
rect 41831 48164 42340 48192
rect 41831 48161 41843 48164
rect 41785 48155 41843 48161
rect 42334 48152 42340 48164
rect 42392 48152 42398 48204
rect 36630 48124 36636 48136
rect 12406 48096 36636 48124
rect 4985 48087 5043 48093
rect 5000 48056 5028 48087
rect 36630 48084 36636 48096
rect 36688 48084 36694 48136
rect 42061 48127 42119 48133
rect 42061 48093 42073 48127
rect 42107 48124 42119 48127
rect 42720 48124 42748 48300
rect 45278 48288 45284 48300
rect 45336 48288 45342 48340
rect 58250 48260 58256 48272
rect 57716 48232 58256 48260
rect 52454 48152 52460 48204
rect 52512 48192 52518 48204
rect 53190 48192 53196 48204
rect 52512 48164 53196 48192
rect 52512 48152 52518 48164
rect 53190 48152 53196 48164
rect 53248 48192 53254 48204
rect 57716 48201 57744 48232
rect 58250 48220 58256 48232
rect 58308 48220 58314 48272
rect 63586 48220 63592 48272
rect 63644 48260 63650 48272
rect 64506 48260 64512 48272
rect 63644 48232 64512 48260
rect 63644 48220 63650 48232
rect 64506 48220 64512 48232
rect 64564 48260 64570 48272
rect 91738 48260 91744 48272
rect 64564 48232 91744 48260
rect 64564 48220 64570 48232
rect 91738 48220 91744 48232
rect 91796 48220 91802 48272
rect 57716 48195 57799 48201
rect 57716 48192 57753 48195
rect 53248 48164 57753 48192
rect 53248 48152 53254 48164
rect 57741 48161 57753 48164
rect 57787 48161 57799 48195
rect 57882 48192 57888 48204
rect 57843 48164 57888 48192
rect 57741 48155 57799 48161
rect 57882 48152 57888 48164
rect 57940 48152 57946 48204
rect 57977 48195 58035 48201
rect 57977 48161 57989 48195
rect 58023 48161 58035 48195
rect 57977 48155 58035 48161
rect 42107 48096 42748 48124
rect 43441 48127 43499 48133
rect 42107 48093 42119 48096
rect 42061 48087 42119 48093
rect 43441 48093 43453 48127
rect 43487 48124 43499 48127
rect 51994 48124 52000 48136
rect 43487 48096 52000 48124
rect 43487 48093 43499 48096
rect 43441 48087 43499 48093
rect 51994 48084 52000 48096
rect 52052 48084 52058 48136
rect 57992 48124 58020 48155
rect 58066 48152 58072 48204
rect 58124 48192 58130 48204
rect 58161 48195 58219 48201
rect 58161 48192 58173 48195
rect 58124 48164 58173 48192
rect 58124 48152 58130 48164
rect 58161 48161 58173 48164
rect 58207 48192 58219 48195
rect 83642 48192 83648 48204
rect 58207 48164 83648 48192
rect 58207 48161 58219 48164
rect 58161 48155 58219 48161
rect 83642 48152 83648 48164
rect 83700 48152 83706 48204
rect 57348 48096 58020 48124
rect 8294 48056 8300 48068
rect 5000 48028 8300 48056
rect 8294 48016 8300 48028
rect 8352 48016 8358 48068
rect 8386 48016 8392 48068
rect 8444 48056 8450 48068
rect 8444 48028 16574 48056
rect 8444 48016 8450 48028
rect 4525 47991 4583 47997
rect 4525 47957 4537 47991
rect 4571 47988 4583 47991
rect 11790 47988 11796 48000
rect 4571 47960 11796 47988
rect 4571 47957 4583 47960
rect 4525 47951 4583 47957
rect 11790 47948 11796 47960
rect 11848 47948 11854 48000
rect 16546 47988 16574 48028
rect 26206 48028 40724 48056
rect 26206 47988 26234 48028
rect 16546 47960 26234 47988
rect 37553 47991 37611 47997
rect 37553 47957 37565 47991
rect 37599 47988 37611 47991
rect 37826 47988 37832 48000
rect 37599 47960 37832 47988
rect 37599 47957 37611 47960
rect 37553 47951 37611 47957
rect 37826 47948 37832 47960
rect 37884 47948 37890 48000
rect 40696 47988 40724 48028
rect 42720 48028 55214 48056
rect 42720 47988 42748 48028
rect 46014 47988 46020 48000
rect 40696 47960 42748 47988
rect 45975 47960 46020 47988
rect 46014 47948 46020 47960
rect 46072 47988 46078 48000
rect 46201 47991 46259 47997
rect 46201 47988 46213 47991
rect 46072 47960 46213 47988
rect 46072 47948 46078 47960
rect 46201 47957 46213 47960
rect 46247 47957 46259 47991
rect 55186 47988 55214 48028
rect 57348 47997 57376 48096
rect 57333 47991 57391 47997
rect 57333 47988 57345 47991
rect 55186 47960 57345 47988
rect 46201 47951 46259 47957
rect 57333 47957 57345 47960
rect 57379 47957 57391 47991
rect 57333 47951 57391 47957
rect 57422 47948 57428 48000
rect 57480 47988 57486 48000
rect 57609 47991 57667 47997
rect 57609 47988 57621 47991
rect 57480 47960 57621 47988
rect 57480 47948 57486 47960
rect 57609 47957 57621 47960
rect 57655 47957 57667 47991
rect 58250 47988 58256 48000
rect 58211 47960 58256 47988
rect 57609 47951 57667 47957
rect 58250 47948 58256 47960
rect 58308 47948 58314 48000
rect 71682 47948 71688 48000
rect 71740 47988 71746 48000
rect 83090 47988 83096 48000
rect 71740 47960 83096 47988
rect 71740 47948 71746 47960
rect 83090 47948 83096 47960
rect 83148 47988 83154 48000
rect 92474 47988 92480 48000
rect 83148 47960 92480 47988
rect 83148 47948 83154 47960
rect 92474 47948 92480 47960
rect 92532 47948 92538 48000
rect 1104 47898 98808 47920
rect 1104 47846 4246 47898
rect 4298 47846 4310 47898
rect 4362 47846 4374 47898
rect 4426 47846 4438 47898
rect 4490 47846 34966 47898
rect 35018 47846 35030 47898
rect 35082 47846 35094 47898
rect 35146 47846 35158 47898
rect 35210 47846 65686 47898
rect 65738 47846 65750 47898
rect 65802 47846 65814 47898
rect 65866 47846 65878 47898
rect 65930 47846 96406 47898
rect 96458 47846 96470 47898
rect 96522 47846 96534 47898
rect 96586 47846 96598 47898
rect 96650 47846 98808 47898
rect 1104 47824 98808 47846
rect 5718 47744 5724 47796
rect 5776 47784 5782 47796
rect 8386 47784 8392 47796
rect 5776 47756 8392 47784
rect 5776 47744 5782 47756
rect 8386 47744 8392 47756
rect 8444 47744 8450 47796
rect 28442 47784 28448 47796
rect 28403 47756 28448 47784
rect 28442 47744 28448 47756
rect 28500 47744 28506 47796
rect 28810 47744 28816 47796
rect 28868 47784 28874 47796
rect 57422 47784 57428 47796
rect 28868 47756 57428 47784
rect 28868 47744 28874 47756
rect 57422 47744 57428 47756
rect 57480 47744 57486 47796
rect 73982 47744 73988 47796
rect 74040 47784 74046 47796
rect 86954 47784 86960 47796
rect 74040 47756 86960 47784
rect 74040 47744 74046 47756
rect 86954 47744 86960 47756
rect 87012 47744 87018 47796
rect 91738 47744 91744 47796
rect 91796 47784 91802 47796
rect 92937 47787 92995 47793
rect 92937 47784 92949 47787
rect 91796 47756 92949 47784
rect 91796 47744 91802 47756
rect 92937 47753 92949 47756
rect 92983 47753 92995 47787
rect 92937 47747 92995 47753
rect 7098 47676 7104 47728
rect 7156 47716 7162 47728
rect 57882 47716 57888 47728
rect 7156 47688 57888 47716
rect 7156 47676 7162 47688
rect 57882 47676 57888 47688
rect 57940 47676 57946 47728
rect 71222 47676 71228 47728
rect 71280 47716 71286 47728
rect 71280 47688 92612 47716
rect 71280 47676 71286 47688
rect 27522 47608 27528 47660
rect 27580 47648 27586 47660
rect 28166 47648 28172 47660
rect 27580 47620 27844 47648
rect 28127 47620 28172 47648
rect 27580 47608 27586 47620
rect 7466 47540 7472 47592
rect 7524 47580 7530 47592
rect 21818 47580 21824 47592
rect 7524 47552 21824 47580
rect 7524 47540 7530 47552
rect 21818 47540 21824 47552
rect 21876 47580 21882 47592
rect 27816 47589 27844 47620
rect 28166 47608 28172 47620
rect 28224 47608 28230 47660
rect 54754 47648 54760 47660
rect 35866 47620 54760 47648
rect 27801 47583 27859 47589
rect 21876 47552 27752 47580
rect 21876 47540 21882 47552
rect 27522 47404 27528 47456
rect 27580 47444 27586 47456
rect 27617 47447 27675 47453
rect 27617 47444 27629 47447
rect 27580 47416 27629 47444
rect 27580 47404 27586 47416
rect 27617 47413 27629 47416
rect 27663 47413 27675 47447
rect 27724 47444 27752 47552
rect 27801 47549 27813 47583
rect 27847 47549 27859 47583
rect 27982 47580 27988 47592
rect 27943 47552 27988 47580
rect 27801 47543 27859 47549
rect 27982 47540 27988 47552
rect 28040 47540 28046 47592
rect 28077 47583 28135 47589
rect 28077 47549 28089 47583
rect 28123 47549 28135 47583
rect 28077 47543 28135 47549
rect 28353 47583 28411 47589
rect 28353 47549 28365 47583
rect 28399 47580 28411 47583
rect 35866 47580 35894 47620
rect 54754 47608 54760 47620
rect 54812 47608 54818 47660
rect 63402 47608 63408 47660
rect 63460 47648 63466 47660
rect 63460 47620 86632 47648
rect 63460 47608 63466 47620
rect 28399 47552 35894 47580
rect 28399 47549 28411 47552
rect 28353 47543 28411 47549
rect 28092 47512 28120 47543
rect 73890 47540 73896 47592
rect 73948 47580 73954 47592
rect 76650 47580 76656 47592
rect 73948 47552 76656 47580
rect 73948 47540 73954 47552
rect 76650 47540 76656 47552
rect 76708 47580 76714 47592
rect 77294 47580 77300 47592
rect 76708 47552 77300 47580
rect 76708 47540 76714 47552
rect 77294 47540 77300 47552
rect 77352 47540 77358 47592
rect 86604 47580 86632 47620
rect 86678 47608 86684 47660
rect 86736 47648 86742 47660
rect 92109 47651 92167 47657
rect 92109 47648 92121 47651
rect 86736 47620 92121 47648
rect 86736 47608 86742 47620
rect 92109 47617 92121 47620
rect 92155 47617 92167 47651
rect 92474 47648 92480 47660
rect 92435 47620 92480 47648
rect 92109 47611 92167 47617
rect 92474 47608 92480 47620
rect 92532 47608 92538 47660
rect 92584 47657 92612 47688
rect 92569 47651 92627 47657
rect 92569 47617 92581 47651
rect 92615 47617 92627 47651
rect 92569 47611 92627 47617
rect 86862 47580 86868 47592
rect 86604 47552 86868 47580
rect 86862 47540 86868 47552
rect 86920 47540 86926 47592
rect 86954 47540 86960 47592
rect 87012 47580 87018 47592
rect 87141 47583 87199 47589
rect 87012 47552 87057 47580
rect 87012 47540 87018 47552
rect 87141 47549 87153 47583
rect 87187 47549 87199 47583
rect 87322 47580 87328 47592
rect 87283 47552 87328 47580
rect 87141 47543 87199 47549
rect 36722 47512 36728 47524
rect 28092 47484 36728 47512
rect 36722 47472 36728 47484
rect 36780 47512 36786 47524
rect 36906 47512 36912 47524
rect 36780 47484 36912 47512
rect 36780 47472 36786 47484
rect 36906 47472 36912 47484
rect 36964 47472 36970 47524
rect 62390 47472 62396 47524
rect 62448 47512 62454 47524
rect 86678 47512 86684 47524
rect 62448 47484 86684 47512
rect 62448 47472 62454 47484
rect 86678 47472 86684 47484
rect 86736 47472 86742 47524
rect 87156 47512 87184 47543
rect 87322 47540 87328 47552
rect 87380 47540 87386 47592
rect 87414 47540 87420 47592
rect 87472 47580 87478 47592
rect 87693 47583 87751 47589
rect 87693 47580 87705 47583
rect 87472 47552 87705 47580
rect 87472 47540 87478 47552
rect 87693 47549 87705 47552
rect 87739 47549 87751 47583
rect 87693 47543 87751 47549
rect 87877 47583 87935 47589
rect 87877 47549 87889 47583
rect 87923 47580 87935 47583
rect 87966 47580 87972 47592
rect 87923 47552 87972 47580
rect 87923 47549 87935 47552
rect 87877 47543 87935 47549
rect 86788 47484 87184 47512
rect 86788 47453 86816 47484
rect 87598 47472 87604 47524
rect 87656 47512 87662 47524
rect 87892 47512 87920 47543
rect 87966 47540 87972 47552
rect 88024 47540 88030 47592
rect 91738 47540 91744 47592
rect 91796 47580 91802 47592
rect 92293 47583 92351 47589
rect 92293 47580 92305 47583
rect 91796 47552 92305 47580
rect 91796 47540 91802 47552
rect 92293 47549 92305 47552
rect 92339 47549 92351 47583
rect 92662 47583 92720 47589
rect 92662 47580 92674 47583
rect 92293 47543 92351 47549
rect 92400 47552 92674 47580
rect 91925 47515 91983 47521
rect 91925 47512 91937 47515
rect 87656 47484 87920 47512
rect 87984 47484 91937 47512
rect 87656 47472 87662 47484
rect 86773 47447 86831 47453
rect 86773 47444 86785 47447
rect 27724 47416 86785 47444
rect 27617 47407 27675 47413
rect 86773 47413 86785 47416
rect 86819 47413 86831 47447
rect 86773 47407 86831 47413
rect 86862 47404 86868 47456
rect 86920 47444 86926 47456
rect 87984 47444 88012 47484
rect 91925 47481 91937 47484
rect 91971 47512 91983 47515
rect 92400 47512 92428 47552
rect 92662 47549 92674 47552
rect 92708 47549 92720 47583
rect 92842 47580 92848 47592
rect 92803 47552 92848 47580
rect 92662 47543 92720 47549
rect 92842 47540 92848 47552
rect 92900 47540 92906 47592
rect 91971 47484 92428 47512
rect 91971 47481 91983 47484
rect 91925 47475 91983 47481
rect 88150 47444 88156 47456
rect 86920 47416 88012 47444
rect 88111 47416 88156 47444
rect 86920 47404 86926 47416
rect 88150 47404 88156 47416
rect 88208 47404 88214 47456
rect 1104 47354 98808 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 50326 47354
rect 50378 47302 50390 47354
rect 50442 47302 50454 47354
rect 50506 47302 50518 47354
rect 50570 47302 81046 47354
rect 81098 47302 81110 47354
rect 81162 47302 81174 47354
rect 81226 47302 81238 47354
rect 81290 47302 98808 47354
rect 1104 47280 98808 47302
rect 8202 47200 8208 47252
rect 8260 47240 8266 47252
rect 17681 47243 17739 47249
rect 17681 47240 17693 47243
rect 8260 47212 17693 47240
rect 8260 47200 8266 47212
rect 17681 47209 17693 47212
rect 17727 47209 17739 47243
rect 17681 47203 17739 47209
rect 31478 47200 31484 47252
rect 31536 47240 31542 47252
rect 88150 47240 88156 47252
rect 31536 47212 88156 47240
rect 31536 47200 31542 47212
rect 88150 47200 88156 47212
rect 88208 47200 88214 47252
rect 38010 47132 38016 47184
rect 38068 47172 38074 47184
rect 64969 47175 65027 47181
rect 64969 47172 64981 47175
rect 38068 47144 64981 47172
rect 38068 47132 38074 47144
rect 64969 47141 64981 47144
rect 65015 47141 65027 47175
rect 64969 47135 65027 47141
rect 74074 47132 74080 47184
rect 74132 47172 74138 47184
rect 74132 47144 77156 47172
rect 74132 47132 74138 47144
rect 77128 47116 77156 47144
rect 77294 47132 77300 47184
rect 77352 47172 77358 47184
rect 87414 47172 87420 47184
rect 77352 47144 87420 47172
rect 77352 47132 77358 47144
rect 87414 47132 87420 47144
rect 87472 47132 87478 47184
rect 14734 47064 14740 47116
rect 14792 47104 14798 47116
rect 16301 47107 16359 47113
rect 16301 47104 16313 47107
rect 14792 47076 16313 47104
rect 14792 47064 14798 47076
rect 16301 47073 16313 47076
rect 16347 47073 16359 47107
rect 16301 47067 16359 47073
rect 37090 47064 37096 47116
rect 37148 47104 37154 47116
rect 64509 47107 64567 47113
rect 64509 47104 64521 47107
rect 37148 47076 64521 47104
rect 37148 47064 37154 47076
rect 64509 47073 64521 47076
rect 64555 47073 64567 47107
rect 64690 47104 64696 47116
rect 64651 47076 64696 47104
rect 64509 47067 64567 47073
rect 16577 47039 16635 47045
rect 16577 47005 16589 47039
rect 16623 47036 16635 47039
rect 50798 47036 50804 47048
rect 16623 47008 50804 47036
rect 16623 47005 16635 47008
rect 16577 46999 16635 47005
rect 50798 46996 50804 47008
rect 50856 46996 50862 47048
rect 64524 47036 64552 47067
rect 64690 47064 64696 47076
rect 64748 47064 64754 47116
rect 64877 47107 64935 47113
rect 64877 47073 64889 47107
rect 64923 47073 64935 47107
rect 65058 47104 65064 47116
rect 65116 47113 65122 47116
rect 65024 47076 65064 47104
rect 64877 47067 64935 47073
rect 64892 47036 64920 47067
rect 65058 47064 65064 47076
rect 65116 47067 65124 47113
rect 75825 47107 75883 47113
rect 75825 47073 75837 47107
rect 75871 47104 75883 47107
rect 76006 47104 76012 47116
rect 75871 47076 76012 47104
rect 75871 47073 75883 47076
rect 75825 47067 75883 47073
rect 65116 47064 65122 47067
rect 76006 47064 76012 47076
rect 76064 47104 76070 47116
rect 76282 47104 76288 47116
rect 76064 47076 76288 47104
rect 76064 47064 76070 47076
rect 76282 47064 76288 47076
rect 76340 47064 76346 47116
rect 77110 47104 77116 47116
rect 77023 47076 77116 47104
rect 77110 47064 77116 47076
rect 77168 47104 77174 47116
rect 87322 47104 87328 47116
rect 77168 47076 87328 47104
rect 77168 47064 77174 47076
rect 87322 47064 87328 47076
rect 87380 47064 87386 47116
rect 64524 47008 64920 47036
rect 68922 46996 68928 47048
rect 68980 47036 68986 47048
rect 76101 47039 76159 47045
rect 76101 47036 76113 47039
rect 68980 47008 76113 47036
rect 68980 46996 68986 47008
rect 76101 47005 76113 47008
rect 76147 47005 76159 47039
rect 76101 46999 76159 47005
rect 17604 46940 17816 46968
rect 9950 46860 9956 46912
rect 10008 46900 10014 46912
rect 17604 46900 17632 46940
rect 10008 46872 17632 46900
rect 17788 46900 17816 46940
rect 27062 46928 27068 46980
rect 27120 46968 27126 46980
rect 27522 46968 27528 46980
rect 27120 46940 27528 46968
rect 27120 46928 27126 46940
rect 27522 46928 27528 46940
rect 27580 46968 27586 46980
rect 58894 46968 58900 46980
rect 27580 46940 58900 46968
rect 27580 46928 27586 46940
rect 58894 46928 58900 46940
rect 58952 46928 58958 46980
rect 65242 46968 65248 46980
rect 64432 46940 64644 46968
rect 65203 46940 65248 46968
rect 34330 46900 34336 46912
rect 17788 46872 34336 46900
rect 10008 46860 10014 46872
rect 34330 46860 34336 46872
rect 34388 46860 34394 46912
rect 45370 46860 45376 46912
rect 45428 46900 45434 46912
rect 64432 46900 64460 46940
rect 45428 46872 64460 46900
rect 64616 46900 64644 46940
rect 65242 46928 65248 46940
rect 65300 46928 65306 46980
rect 73246 46900 73252 46912
rect 64616 46872 73252 46900
rect 45428 46860 45434 46872
rect 73246 46860 73252 46872
rect 73304 46860 73310 46912
rect 79502 46860 79508 46912
rect 79560 46900 79566 46912
rect 81526 46900 81532 46912
rect 79560 46872 81532 46900
rect 79560 46860 79566 46872
rect 81526 46860 81532 46872
rect 81584 46860 81590 46912
rect 1104 46810 98808 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 65686 46810
rect 65738 46758 65750 46810
rect 65802 46758 65814 46810
rect 65866 46758 65878 46810
rect 65930 46758 96406 46810
rect 96458 46758 96470 46810
rect 96522 46758 96534 46810
rect 96586 46758 96598 46810
rect 96650 46758 98808 46810
rect 1104 46736 98808 46758
rect 11882 46656 11888 46708
rect 11940 46696 11946 46708
rect 14826 46696 14832 46708
rect 11940 46668 14832 46696
rect 11940 46656 11946 46668
rect 14826 46656 14832 46668
rect 14884 46656 14890 46708
rect 25682 46656 25688 46708
rect 25740 46696 25746 46708
rect 75822 46696 75828 46708
rect 25740 46668 75828 46696
rect 25740 46656 25746 46668
rect 75822 46656 75828 46668
rect 75880 46656 75886 46708
rect 76006 46656 76012 46708
rect 76064 46696 76070 46708
rect 86957 46699 87015 46705
rect 86957 46696 86969 46699
rect 76064 46668 86969 46696
rect 76064 46656 76070 46668
rect 86957 46665 86969 46668
rect 87003 46665 87015 46699
rect 86957 46659 87015 46665
rect 18414 46628 18420 46640
rect 14660 46600 18420 46628
rect 14660 46569 14688 46600
rect 18414 46588 18420 46600
rect 18472 46628 18478 46640
rect 96890 46628 96896 46640
rect 18472 46600 96896 46628
rect 18472 46588 18478 46600
rect 96890 46588 96896 46600
rect 96948 46588 96954 46640
rect 13357 46563 13415 46569
rect 13357 46529 13369 46563
rect 13403 46560 13415 46563
rect 14645 46563 14703 46569
rect 14645 46560 14657 46563
rect 13403 46532 14657 46560
rect 13403 46529 13415 46532
rect 13357 46523 13415 46529
rect 14645 46529 14657 46532
rect 14691 46529 14703 46563
rect 19242 46560 19248 46572
rect 19203 46532 19248 46560
rect 14645 46523 14703 46529
rect 19242 46520 19248 46532
rect 19300 46520 19306 46572
rect 43254 46520 43260 46572
rect 43312 46560 43318 46572
rect 71774 46560 71780 46572
rect 43312 46532 71780 46560
rect 43312 46520 43318 46532
rect 71774 46520 71780 46532
rect 71832 46520 71838 46572
rect 74258 46520 74264 46572
rect 74316 46560 74322 46572
rect 87325 46563 87383 46569
rect 87325 46560 87337 46563
rect 74316 46532 87337 46560
rect 74316 46520 74322 46532
rect 87325 46529 87337 46532
rect 87371 46529 87383 46563
rect 87325 46523 87383 46529
rect 87432 46532 87920 46560
rect 14093 46495 14151 46501
rect 14093 46461 14105 46495
rect 14139 46461 14151 46495
rect 14093 46455 14151 46461
rect 14185 46495 14243 46501
rect 14185 46461 14197 46495
rect 14231 46461 14243 46495
rect 14185 46455 14243 46461
rect 14461 46495 14519 46501
rect 14461 46461 14473 46495
rect 14507 46492 14519 46495
rect 14734 46492 14740 46504
rect 14507 46464 14740 46492
rect 14507 46461 14519 46464
rect 14461 46455 14519 46461
rect 13630 46356 13636 46368
rect 13591 46328 13636 46356
rect 13630 46316 13636 46328
rect 13688 46316 13694 46368
rect 14108 46356 14136 46455
rect 14200 46424 14228 46455
rect 14734 46452 14740 46464
rect 14792 46452 14798 46504
rect 14826 46452 14832 46504
rect 14884 46492 14890 46504
rect 18690 46492 18696 46504
rect 14884 46464 14929 46492
rect 18651 46464 18696 46492
rect 14884 46452 14890 46464
rect 18690 46452 18696 46464
rect 18748 46452 18754 46504
rect 86957 46495 87015 46501
rect 19444 46464 26234 46492
rect 19444 46424 19472 46464
rect 14200 46396 19472 46424
rect 26206 46424 26234 46464
rect 86957 46461 86969 46495
rect 87003 46492 87015 46495
rect 87141 46495 87199 46501
rect 87141 46492 87153 46495
rect 87003 46464 87153 46492
rect 87003 46461 87015 46464
rect 86957 46455 87015 46461
rect 87141 46461 87153 46464
rect 87187 46461 87199 46495
rect 87141 46455 87199 46461
rect 66162 46424 66168 46436
rect 26206 46396 66168 46424
rect 66162 46384 66168 46396
rect 66220 46384 66226 46436
rect 81526 46384 81532 46436
rect 81584 46424 81590 46436
rect 87432 46424 87460 46532
rect 87509 46495 87567 46501
rect 87509 46461 87521 46495
rect 87555 46461 87567 46495
rect 87782 46492 87788 46504
rect 87743 46464 87788 46492
rect 87509 46455 87567 46461
rect 81584 46396 87460 46424
rect 81584 46384 81590 46396
rect 16482 46356 16488 46368
rect 14108 46328 16488 46356
rect 16482 46316 16488 46328
rect 16540 46316 16546 46368
rect 71222 46316 71228 46368
rect 71280 46356 71286 46368
rect 74258 46356 74264 46368
rect 71280 46328 74264 46356
rect 71280 46316 71286 46328
rect 74258 46316 74264 46328
rect 74316 46316 74322 46368
rect 84838 46316 84844 46368
rect 84896 46356 84902 46368
rect 87524 46356 87552 46455
rect 87782 46452 87788 46464
rect 87840 46452 87846 46504
rect 87892 46501 87920 46532
rect 88150 46520 88156 46572
rect 88208 46560 88214 46572
rect 88245 46563 88303 46569
rect 88245 46560 88257 46563
rect 88208 46532 88257 46560
rect 88208 46520 88214 46532
rect 88245 46529 88257 46532
rect 88291 46529 88303 46563
rect 88245 46523 88303 46529
rect 87877 46495 87935 46501
rect 87877 46461 87889 46495
rect 87923 46461 87935 46495
rect 87877 46455 87935 46461
rect 84896 46328 87552 46356
rect 84896 46316 84902 46328
rect 1104 46266 98808 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 50326 46266
rect 50378 46214 50390 46266
rect 50442 46214 50454 46266
rect 50506 46214 50518 46266
rect 50570 46214 81046 46266
rect 81098 46214 81110 46266
rect 81162 46214 81174 46266
rect 81226 46214 81238 46266
rect 81290 46214 98808 46266
rect 1104 46192 98808 46214
rect 11238 46112 11244 46164
rect 11296 46152 11302 46164
rect 11606 46152 11612 46164
rect 11296 46124 11612 46152
rect 11296 46112 11302 46124
rect 11606 46112 11612 46124
rect 11664 46112 11670 46164
rect 14734 46112 14740 46164
rect 14792 46152 14798 46164
rect 16942 46152 16948 46164
rect 14792 46124 16948 46152
rect 14792 46112 14798 46124
rect 16942 46112 16948 46124
rect 17000 46112 17006 46164
rect 53558 46112 53564 46164
rect 53616 46152 53622 46164
rect 60366 46152 60372 46164
rect 53616 46124 60372 46152
rect 53616 46112 53622 46124
rect 60366 46112 60372 46124
rect 60424 46112 60430 46164
rect 9674 46044 9680 46096
rect 9732 46084 9738 46096
rect 18690 46084 18696 46096
rect 9732 46056 18696 46084
rect 9732 46044 9738 46056
rect 18690 46044 18696 46056
rect 18748 46044 18754 46096
rect 34330 46044 34336 46096
rect 34388 46084 34394 46096
rect 87782 46084 87788 46096
rect 34388 46056 87788 46084
rect 34388 46044 34394 46056
rect 87782 46044 87788 46056
rect 87840 46044 87846 46096
rect 13630 45976 13636 46028
rect 13688 46016 13694 46028
rect 90542 46016 90548 46028
rect 13688 45988 90548 46016
rect 13688 45976 13694 45988
rect 90542 45976 90548 45988
rect 90600 45976 90606 46028
rect 77662 45772 77668 45824
rect 77720 45812 77726 45824
rect 85942 45812 85948 45824
rect 77720 45784 85948 45812
rect 77720 45772 77726 45784
rect 85942 45772 85948 45784
rect 86000 45772 86006 45824
rect 1104 45722 98808 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 65686 45722
rect 65738 45670 65750 45722
rect 65802 45670 65814 45722
rect 65866 45670 65878 45722
rect 65930 45670 96406 45722
rect 96458 45670 96470 45722
rect 96522 45670 96534 45722
rect 96586 45670 96598 45722
rect 96650 45670 98808 45722
rect 1104 45648 98808 45670
rect 76300 45580 77248 45608
rect 3050 45500 3056 45552
rect 3108 45540 3114 45552
rect 76300 45540 76328 45580
rect 3108 45512 12434 45540
rect 3108 45500 3114 45512
rect 7469 45475 7527 45481
rect 7469 45441 7481 45475
rect 7515 45472 7527 45475
rect 10318 45472 10324 45484
rect 7515 45444 10324 45472
rect 7515 45441 7527 45444
rect 7469 45435 7527 45441
rect 10318 45432 10324 45444
rect 10376 45432 10382 45484
rect 12406 45472 12434 45512
rect 76208 45512 76328 45540
rect 77220 45540 77248 45580
rect 77846 45568 77852 45620
rect 77904 45608 77910 45620
rect 77904 45580 86954 45608
rect 77904 45568 77910 45580
rect 77662 45540 77668 45552
rect 77220 45512 77668 45540
rect 17310 45472 17316 45484
rect 12406 45444 17316 45472
rect 17310 45432 17316 45444
rect 17368 45432 17374 45484
rect 41874 45432 41880 45484
rect 41932 45472 41938 45484
rect 76208 45472 76236 45512
rect 77662 45500 77668 45512
rect 77720 45500 77726 45552
rect 86926 45540 86954 45580
rect 90450 45540 90456 45552
rect 86926 45512 90456 45540
rect 90450 45500 90456 45512
rect 90508 45500 90514 45552
rect 76285 45475 76343 45481
rect 76285 45472 76297 45475
rect 41932 45444 70394 45472
rect 76208 45444 76297 45472
rect 41932 45432 41938 45444
rect 6638 45364 6644 45416
rect 6696 45404 6702 45416
rect 6917 45407 6975 45413
rect 6917 45404 6929 45407
rect 6696 45376 6929 45404
rect 6696 45364 6702 45376
rect 6917 45373 6929 45376
rect 6963 45373 6975 45407
rect 6917 45367 6975 45373
rect 26878 45364 26884 45416
rect 26936 45404 26942 45416
rect 47578 45404 47584 45416
rect 26936 45376 47584 45404
rect 26936 45364 26942 45376
rect 47578 45364 47584 45376
rect 47636 45364 47642 45416
rect 70366 45404 70394 45444
rect 76285 45441 76297 45444
rect 76331 45441 76343 45475
rect 77846 45472 77852 45484
rect 76285 45435 76343 45441
rect 76392 45444 77852 45472
rect 76392 45404 76420 45444
rect 77846 45432 77852 45444
rect 77904 45432 77910 45484
rect 70366 45376 76420 45404
rect 76561 45407 76619 45413
rect 76561 45373 76573 45407
rect 76607 45404 76619 45407
rect 76607 45376 77248 45404
rect 76607 45373 76619 45376
rect 76561 45367 76619 45373
rect 7650 45296 7656 45348
rect 7708 45336 7714 45348
rect 18138 45336 18144 45348
rect 7708 45308 18144 45336
rect 7708 45296 7714 45308
rect 18138 45296 18144 45308
rect 18196 45336 18202 45348
rect 40310 45336 40316 45348
rect 18196 45308 40316 45336
rect 18196 45296 18202 45308
rect 40310 45296 40316 45308
rect 40368 45296 40374 45348
rect 63126 45296 63132 45348
rect 63184 45336 63190 45348
rect 74258 45336 74264 45348
rect 63184 45308 74264 45336
rect 63184 45296 63190 45308
rect 74258 45296 74264 45308
rect 74316 45296 74322 45348
rect 77220 45336 77248 45376
rect 82262 45336 82268 45348
rect 77220 45308 82268 45336
rect 82262 45296 82268 45308
rect 82320 45296 82326 45348
rect 15102 45228 15108 45280
rect 15160 45268 15166 45280
rect 21358 45268 21364 45280
rect 15160 45240 21364 45268
rect 15160 45228 15166 45240
rect 21358 45228 21364 45240
rect 21416 45228 21422 45280
rect 23290 45228 23296 45280
rect 23348 45268 23354 45280
rect 44266 45268 44272 45280
rect 23348 45240 44272 45268
rect 23348 45228 23354 45240
rect 44266 45228 44272 45240
rect 44324 45228 44330 45280
rect 57882 45228 57888 45280
rect 57940 45268 57946 45280
rect 77665 45271 77723 45277
rect 77665 45268 77677 45271
rect 57940 45240 77677 45268
rect 57940 45228 57946 45240
rect 77665 45237 77677 45240
rect 77711 45268 77723 45271
rect 82446 45268 82452 45280
rect 77711 45240 82452 45268
rect 77711 45237 77723 45240
rect 77665 45231 77723 45237
rect 82446 45228 82452 45240
rect 82504 45228 82510 45280
rect 1104 45178 98808 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 50326 45178
rect 50378 45126 50390 45178
rect 50442 45126 50454 45178
rect 50506 45126 50518 45178
rect 50570 45126 81046 45178
rect 81098 45126 81110 45178
rect 81162 45126 81174 45178
rect 81226 45126 81238 45178
rect 81290 45126 98808 45178
rect 1104 45104 98808 45126
rect 8110 45024 8116 45076
rect 8168 45064 8174 45076
rect 58894 45064 58900 45076
rect 8168 45036 58900 45064
rect 8168 45024 8174 45036
rect 58894 45024 58900 45036
rect 58952 45064 58958 45076
rect 70670 45064 70676 45076
rect 58952 45036 70676 45064
rect 58952 45024 58958 45036
rect 70670 45024 70676 45036
rect 70728 45064 70734 45076
rect 70728 45036 72648 45064
rect 70728 45024 70734 45036
rect 4798 44956 4804 45008
rect 4856 44996 4862 45008
rect 4856 44968 16574 44996
rect 4856 44956 4862 44968
rect 6457 44931 6515 44937
rect 6457 44897 6469 44931
rect 6503 44928 6515 44931
rect 6825 44931 6883 44937
rect 6825 44928 6837 44931
rect 6503 44900 6837 44928
rect 6503 44897 6515 44900
rect 6457 44891 6515 44897
rect 6825 44897 6837 44900
rect 6871 44928 6883 44931
rect 7650 44928 7656 44940
rect 6871 44900 7656 44928
rect 6871 44897 6883 44900
rect 6825 44891 6883 44897
rect 7650 44888 7656 44900
rect 7708 44888 7714 44940
rect 16546 44860 16574 44968
rect 17310 44956 17316 45008
rect 17368 44996 17374 45008
rect 18049 44999 18107 45005
rect 18049 44996 18061 44999
rect 17368 44968 18061 44996
rect 17368 44956 17374 44968
rect 18049 44965 18061 44968
rect 18095 44965 18107 44999
rect 18049 44959 18107 44965
rect 21358 44956 21364 45008
rect 21416 44996 21422 45008
rect 72510 44996 72516 45008
rect 21416 44968 72516 44996
rect 21416 44956 21422 44968
rect 72510 44956 72516 44968
rect 72568 44956 72574 45008
rect 17860 44931 17918 44937
rect 17860 44897 17872 44931
rect 17906 44897 17918 44931
rect 17860 44891 17918 44897
rect 17880 44860 17908 44891
rect 17954 44888 17960 44940
rect 18012 44928 18018 44940
rect 18230 44928 18236 44940
rect 18012 44900 18057 44928
rect 18143 44900 18236 44928
rect 18012 44888 18018 44900
rect 18230 44888 18236 44900
rect 18288 44928 18294 44940
rect 19242 44928 19248 44940
rect 18288 44900 19248 44928
rect 18288 44888 18294 44900
rect 19242 44888 19248 44900
rect 19300 44928 19306 44940
rect 57974 44928 57980 44940
rect 19300 44900 57980 44928
rect 19300 44888 19306 44900
rect 57974 44888 57980 44900
rect 58032 44888 58038 44940
rect 72620 44928 72648 45036
rect 74258 44996 74264 45008
rect 74219 44968 74264 44996
rect 74258 44956 74264 44968
rect 74316 44956 74322 45008
rect 73154 44928 73160 44940
rect 72620 44900 73160 44928
rect 73154 44888 73160 44900
rect 73212 44928 73218 44940
rect 74077 44931 74135 44937
rect 74077 44928 74089 44931
rect 73212 44900 74089 44928
rect 73212 44888 73218 44900
rect 74077 44897 74089 44900
rect 74123 44897 74135 44931
rect 74077 44891 74135 44897
rect 74353 44931 74411 44937
rect 74353 44897 74365 44931
rect 74399 44897 74411 44931
rect 74353 44891 74411 44897
rect 18598 44860 18604 44872
rect 16546 44832 17816 44860
rect 17880 44832 18604 44860
rect 4614 44752 4620 44804
rect 4672 44792 4678 44804
rect 17681 44795 17739 44801
rect 17681 44792 17693 44795
rect 4672 44764 12434 44792
rect 4672 44752 4678 44764
rect 1670 44724 1676 44736
rect 1631 44696 1676 44724
rect 1670 44684 1676 44696
rect 1728 44724 1734 44736
rect 1949 44727 2007 44733
rect 1949 44724 1961 44727
rect 1728 44696 1961 44724
rect 1728 44684 1734 44696
rect 1949 44693 1961 44696
rect 1995 44693 2007 44727
rect 6638 44724 6644 44736
rect 6599 44696 6644 44724
rect 1949 44687 2007 44693
rect 6638 44684 6644 44696
rect 6696 44684 6702 44736
rect 12406 44724 12434 44764
rect 16546 44764 17693 44792
rect 16546 44724 16574 44764
rect 17681 44761 17693 44764
rect 17727 44761 17739 44795
rect 17788 44792 17816 44832
rect 18598 44820 18604 44832
rect 18656 44820 18662 44872
rect 32398 44820 32404 44872
rect 32456 44860 32462 44872
rect 54754 44860 54760 44872
rect 32456 44832 54760 44860
rect 32456 44820 32462 44832
rect 54754 44820 54760 44832
rect 54812 44820 54818 44872
rect 64782 44820 64788 44872
rect 64840 44860 64846 44872
rect 74368 44860 74396 44891
rect 74442 44888 74448 44940
rect 74500 44937 74506 44940
rect 74500 44928 74508 44937
rect 74500 44900 74545 44928
rect 74500 44891 74508 44900
rect 74500 44888 74506 44891
rect 64840 44832 74396 44860
rect 64840 44820 64846 44832
rect 17954 44792 17960 44804
rect 17788 44764 17960 44792
rect 17681 44755 17739 44761
rect 17954 44752 17960 44764
rect 18012 44752 18018 44804
rect 12406 44696 16574 44724
rect 17497 44727 17555 44733
rect 17497 44693 17509 44727
rect 17543 44724 17555 44727
rect 18230 44724 18236 44736
rect 17543 44696 18236 44724
rect 17543 44693 17555 44696
rect 17497 44687 17555 44693
rect 18230 44684 18236 44696
rect 18288 44684 18294 44736
rect 21729 44727 21787 44733
rect 21729 44693 21741 44727
rect 21775 44724 21787 44727
rect 22005 44727 22063 44733
rect 22005 44724 22017 44727
rect 21775 44696 22017 44724
rect 21775 44693 21787 44696
rect 21729 44687 21787 44693
rect 22005 44693 22017 44696
rect 22051 44724 22063 44727
rect 45922 44724 45928 44736
rect 22051 44696 45928 44724
rect 22051 44693 22063 44696
rect 22005 44687 22063 44693
rect 45922 44684 45928 44696
rect 45980 44684 45986 44736
rect 74626 44724 74632 44736
rect 74587 44696 74632 44724
rect 74626 44684 74632 44696
rect 74684 44684 74690 44736
rect 1104 44634 98808 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 65686 44634
rect 65738 44582 65750 44634
rect 65802 44582 65814 44634
rect 65866 44582 65878 44634
rect 65930 44582 96406 44634
rect 96458 44582 96470 44634
rect 96522 44582 96534 44634
rect 96586 44582 96598 44634
rect 96650 44582 98808 44634
rect 1104 44560 98808 44582
rect 40310 44412 40316 44464
rect 40368 44452 40374 44464
rect 41874 44452 41880 44464
rect 40368 44424 41880 44452
rect 40368 44412 40374 44424
rect 41874 44412 41880 44424
rect 41932 44412 41938 44464
rect 70486 44384 70492 44396
rect 64846 44356 70492 44384
rect 17678 44276 17684 44328
rect 17736 44316 17742 44328
rect 23293 44319 23351 44325
rect 23293 44316 23305 44319
rect 17736 44288 23305 44316
rect 17736 44276 17742 44288
rect 23293 44285 23305 44288
rect 23339 44285 23351 44319
rect 23566 44316 23572 44328
rect 23527 44288 23572 44316
rect 23293 44279 23351 44285
rect 23566 44276 23572 44288
rect 23624 44276 23630 44328
rect 58069 44319 58127 44325
rect 58069 44285 58081 44319
rect 58115 44316 58127 44319
rect 58345 44319 58403 44325
rect 58345 44316 58357 44319
rect 58115 44288 58357 44316
rect 58115 44285 58127 44288
rect 58069 44279 58127 44285
rect 58345 44285 58357 44288
rect 58391 44316 58403 44319
rect 62850 44316 62856 44328
rect 58391 44288 62856 44316
rect 58391 44285 58403 44288
rect 58345 44279 58403 44285
rect 62850 44276 62856 44288
rect 62908 44276 62914 44328
rect 44266 44208 44272 44260
rect 44324 44248 44330 44260
rect 45094 44248 45100 44260
rect 44324 44220 45100 44248
rect 44324 44208 44330 44220
rect 45094 44208 45100 44220
rect 45152 44248 45158 44260
rect 64846 44248 64874 44356
rect 70486 44344 70492 44356
rect 70544 44384 70550 44396
rect 71682 44384 71688 44396
rect 70544 44356 71688 44384
rect 70544 44344 70550 44356
rect 71682 44344 71688 44356
rect 71740 44344 71746 44396
rect 69753 44319 69811 44325
rect 69753 44285 69765 44319
rect 69799 44285 69811 44319
rect 69753 44279 69811 44285
rect 45152 44220 64874 44248
rect 45152 44208 45158 44220
rect 24854 44180 24860 44192
rect 24815 44152 24860 44180
rect 24854 44140 24860 44152
rect 24912 44140 24918 44192
rect 46842 44140 46848 44192
rect 46900 44180 46906 44192
rect 53742 44180 53748 44192
rect 46900 44152 53748 44180
rect 46900 44140 46906 44152
rect 53742 44140 53748 44152
rect 53800 44140 53806 44192
rect 69566 44180 69572 44192
rect 69527 44152 69572 44180
rect 69566 44140 69572 44152
rect 69624 44180 69630 44192
rect 69768 44180 69796 44279
rect 69624 44152 69796 44180
rect 69624 44140 69630 44152
rect 84930 44140 84936 44192
rect 84988 44180 84994 44192
rect 86494 44180 86500 44192
rect 84988 44152 86500 44180
rect 84988 44140 84994 44152
rect 86494 44140 86500 44152
rect 86552 44140 86558 44192
rect 1104 44090 98808 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 50326 44090
rect 50378 44038 50390 44090
rect 50442 44038 50454 44090
rect 50506 44038 50518 44090
rect 50570 44038 81046 44090
rect 81098 44038 81110 44090
rect 81162 44038 81174 44090
rect 81226 44038 81238 44090
rect 81290 44038 98808 44090
rect 1104 44016 98808 44038
rect 10410 43936 10416 43988
rect 10468 43976 10474 43988
rect 39758 43976 39764 43988
rect 10468 43948 39764 43976
rect 10468 43936 10474 43948
rect 39758 43936 39764 43948
rect 39816 43936 39822 43988
rect 72418 43936 72424 43988
rect 72476 43976 72482 43988
rect 72970 43976 72976 43988
rect 72476 43948 72976 43976
rect 72476 43936 72482 43948
rect 72970 43936 72976 43948
rect 73028 43936 73034 43988
rect 74074 43936 74080 43988
rect 74132 43976 74138 43988
rect 78122 43976 78128 43988
rect 74132 43948 78128 43976
rect 74132 43936 74138 43948
rect 78122 43936 78128 43948
rect 78180 43936 78186 43988
rect 64322 43868 64328 43920
rect 64380 43908 64386 43920
rect 66714 43908 66720 43920
rect 64380 43880 66720 43908
rect 64380 43868 64386 43880
rect 66714 43868 66720 43880
rect 66772 43868 66778 43920
rect 24578 43800 24584 43852
rect 24636 43840 24642 43852
rect 25225 43843 25283 43849
rect 25225 43840 25237 43843
rect 24636 43812 25237 43840
rect 24636 43800 24642 43812
rect 25225 43809 25237 43812
rect 25271 43809 25283 43843
rect 25225 43803 25283 43809
rect 26206 43812 45554 43840
rect 24486 43732 24492 43784
rect 24544 43772 24550 43784
rect 25593 43775 25651 43781
rect 25593 43772 25605 43775
rect 24544 43744 25605 43772
rect 24544 43732 24550 43744
rect 25593 43741 25605 43744
rect 25639 43772 25651 43775
rect 26206 43772 26234 43812
rect 25639 43744 26234 43772
rect 25639 43741 25651 43744
rect 25593 43735 25651 43741
rect 31018 43732 31024 43784
rect 31076 43772 31082 43784
rect 37277 43775 37335 43781
rect 37277 43772 37289 43775
rect 31076 43744 37289 43772
rect 31076 43732 31082 43744
rect 37277 43741 37289 43744
rect 37323 43741 37335 43775
rect 37550 43772 37556 43784
rect 37511 43744 37556 43772
rect 37277 43735 37335 43741
rect 37550 43732 37556 43744
rect 37608 43732 37614 43784
rect 45526 43772 45554 43812
rect 59538 43772 59544 43784
rect 45526 43744 59544 43772
rect 59538 43732 59544 43744
rect 59596 43732 59602 43784
rect 38838 43704 38844 43716
rect 38799 43676 38844 43704
rect 38838 43664 38844 43676
rect 38896 43664 38902 43716
rect 40034 43664 40040 43716
rect 40092 43704 40098 43716
rect 69198 43704 69204 43716
rect 40092 43676 69204 43704
rect 40092 43664 40098 43676
rect 69198 43664 69204 43676
rect 69256 43664 69262 43716
rect 23201 43639 23259 43645
rect 23201 43605 23213 43639
rect 23247 43636 23259 43639
rect 23477 43639 23535 43645
rect 23477 43636 23489 43639
rect 23247 43608 23489 43636
rect 23247 43605 23259 43608
rect 23201 43599 23259 43605
rect 23477 43605 23489 43608
rect 23523 43636 23535 43639
rect 63126 43636 63132 43648
rect 23523 43608 63132 43636
rect 23523 43605 23535 43608
rect 23477 43599 23535 43605
rect 63126 43596 63132 43608
rect 63184 43596 63190 43648
rect 1104 43546 98808 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 65686 43546
rect 65738 43494 65750 43546
rect 65802 43494 65814 43546
rect 65866 43494 65878 43546
rect 65930 43494 96406 43546
rect 96458 43494 96470 43546
rect 96522 43494 96534 43546
rect 96586 43494 96598 43546
rect 96650 43494 98808 43546
rect 1104 43472 98808 43494
rect 7650 43392 7656 43444
rect 7708 43432 7714 43444
rect 35250 43432 35256 43444
rect 7708 43404 35256 43432
rect 7708 43392 7714 43404
rect 35250 43392 35256 43404
rect 35308 43392 35314 43444
rect 38838 43392 38844 43444
rect 38896 43432 38902 43444
rect 50798 43432 50804 43444
rect 38896 43404 50804 43432
rect 38896 43392 38902 43404
rect 50798 43392 50804 43404
rect 50856 43392 50862 43444
rect 52178 43392 52184 43444
rect 52236 43432 52242 43444
rect 82354 43432 82360 43444
rect 52236 43404 82360 43432
rect 52236 43392 52242 43404
rect 82354 43392 82360 43404
rect 82412 43392 82418 43444
rect 16482 43324 16488 43376
rect 16540 43364 16546 43376
rect 38654 43364 38660 43376
rect 16540 43336 38660 43364
rect 16540 43324 16546 43336
rect 38654 43324 38660 43336
rect 38712 43324 38718 43376
rect 29822 43256 29828 43308
rect 29880 43296 29886 43308
rect 38856 43296 38884 43392
rect 40034 43364 40040 43376
rect 39995 43336 40040 43364
rect 40034 43324 40040 43336
rect 40092 43324 40098 43376
rect 45094 43296 45100 43308
rect 29880 43268 38884 43296
rect 45055 43268 45100 43296
rect 29880 43256 29886 43268
rect 45094 43256 45100 43268
rect 45152 43256 45158 43308
rect 59357 43299 59415 43305
rect 59357 43265 59369 43299
rect 59403 43296 59415 43299
rect 82538 43296 82544 43308
rect 59403 43268 82544 43296
rect 59403 43265 59415 43268
rect 59357 43259 59415 43265
rect 82538 43256 82544 43268
rect 82596 43256 82602 43308
rect 94038 43296 94044 43308
rect 84166 43268 94044 43296
rect 40218 43228 40224 43240
rect 40179 43200 40224 43228
rect 40218 43188 40224 43200
rect 40276 43188 40282 43240
rect 40405 43231 40463 43237
rect 40405 43197 40417 43231
rect 40451 43228 40463 43231
rect 44726 43228 44732 43240
rect 40451 43200 41828 43228
rect 44687 43200 44732 43228
rect 40451 43197 40463 43200
rect 40405 43191 40463 43197
rect 40494 43160 40500 43172
rect 40455 43132 40500 43160
rect 40494 43120 40500 43132
rect 40552 43120 40558 43172
rect 41800 43160 41828 43200
rect 44726 43188 44732 43200
rect 44784 43188 44790 43240
rect 59538 43228 59544 43240
rect 59451 43200 59544 43228
rect 59538 43188 59544 43200
rect 59596 43228 59602 43240
rect 84166 43228 84194 43268
rect 94038 43256 94044 43268
rect 94096 43256 94102 43308
rect 59596 43200 84194 43228
rect 88705 43231 88763 43237
rect 59596 43188 59602 43200
rect 88705 43197 88717 43231
rect 88751 43197 88763 43231
rect 88705 43191 88763 43197
rect 53650 43160 53656 43172
rect 41800 43132 53656 43160
rect 53650 43120 53656 43132
rect 53708 43120 53714 43172
rect 56042 43120 56048 43172
rect 56100 43160 56106 43172
rect 59817 43163 59875 43169
rect 59817 43160 59829 43163
rect 56100 43132 59829 43160
rect 56100 43120 56106 43132
rect 59817 43129 59829 43132
rect 59863 43129 59875 43163
rect 59817 43123 59875 43129
rect 40512 43092 40540 43120
rect 55122 43092 55128 43104
rect 40512 43064 55128 43092
rect 55122 43052 55128 43064
rect 55180 43052 55186 43104
rect 58342 43052 58348 43104
rect 58400 43092 58406 43104
rect 58618 43092 58624 43104
rect 58400 43064 58624 43092
rect 58400 43052 58406 43064
rect 58618 43052 58624 43064
rect 58676 43092 58682 43104
rect 59725 43095 59783 43101
rect 59725 43092 59737 43095
rect 58676 43064 59737 43092
rect 58676 43052 58682 43064
rect 59725 43061 59737 43064
rect 59771 43061 59783 43095
rect 59725 43055 59783 43061
rect 71130 43052 71136 43104
rect 71188 43092 71194 43104
rect 88521 43095 88579 43101
rect 88521 43092 88533 43095
rect 71188 43064 88533 43092
rect 71188 43052 71194 43064
rect 88521 43061 88533 43064
rect 88567 43092 88579 43095
rect 88720 43092 88748 43191
rect 88567 43064 88748 43092
rect 88567 43061 88579 43064
rect 88521 43055 88579 43061
rect 1104 43002 98808 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 50326 43002
rect 50378 42950 50390 43002
rect 50442 42950 50454 43002
rect 50506 42950 50518 43002
rect 50570 42950 81046 43002
rect 81098 42950 81110 43002
rect 81162 42950 81174 43002
rect 81226 42950 81238 43002
rect 81290 42950 98808 43002
rect 1104 42928 98808 42950
rect 38654 42848 38660 42900
rect 38712 42888 38718 42900
rect 42886 42888 42892 42900
rect 38712 42860 42892 42888
rect 38712 42848 38718 42860
rect 42886 42848 42892 42860
rect 42944 42888 42950 42900
rect 72418 42888 72424 42900
rect 42944 42860 72424 42888
rect 42944 42848 42950 42860
rect 72418 42848 72424 42860
rect 72476 42848 72482 42900
rect 17402 42780 17408 42832
rect 17460 42820 17466 42832
rect 80882 42820 80888 42832
rect 17460 42792 80888 42820
rect 17460 42780 17466 42792
rect 80882 42780 80888 42792
rect 80940 42820 80946 42832
rect 85574 42820 85580 42832
rect 80940 42792 85580 42820
rect 80940 42780 80946 42792
rect 85574 42780 85580 42792
rect 85632 42780 85638 42832
rect 12066 42712 12072 42764
rect 12124 42752 12130 42764
rect 12250 42752 12256 42764
rect 12124 42724 12256 42752
rect 12124 42712 12130 42724
rect 12250 42712 12256 42724
rect 12308 42752 12314 42764
rect 46106 42752 46112 42764
rect 12308 42724 46112 42752
rect 12308 42712 12314 42724
rect 46106 42712 46112 42724
rect 46164 42752 46170 42764
rect 49418 42752 49424 42764
rect 46164 42724 49424 42752
rect 46164 42712 46170 42724
rect 49418 42712 49424 42724
rect 49476 42712 49482 42764
rect 60734 42712 60740 42764
rect 60792 42752 60798 42764
rect 73157 42755 73215 42761
rect 73157 42752 73169 42755
rect 60792 42724 73169 42752
rect 60792 42712 60798 42724
rect 73157 42721 73169 42724
rect 73203 42721 73215 42755
rect 73522 42752 73528 42764
rect 73483 42724 73528 42752
rect 73157 42715 73215 42721
rect 73522 42712 73528 42724
rect 73580 42712 73586 42764
rect 73709 42755 73767 42761
rect 73709 42721 73721 42755
rect 73755 42752 73767 42755
rect 74442 42752 74448 42764
rect 73755 42724 74448 42752
rect 73755 42721 73767 42724
rect 73709 42715 73767 42721
rect 74442 42712 74448 42724
rect 74500 42712 74506 42764
rect 78674 42712 78680 42764
rect 78732 42752 78738 42764
rect 79962 42752 79968 42764
rect 78732 42724 79968 42752
rect 78732 42712 78738 42724
rect 79962 42712 79968 42724
rect 80020 42752 80026 42764
rect 80517 42755 80575 42761
rect 80517 42752 80529 42755
rect 80020 42724 80529 42752
rect 80020 42712 80026 42724
rect 80517 42721 80529 42724
rect 80563 42721 80575 42755
rect 80517 42715 80575 42721
rect 86218 42712 86224 42764
rect 86276 42752 86282 42764
rect 91649 42755 91707 42761
rect 91649 42752 91661 42755
rect 86276 42724 91661 42752
rect 86276 42712 86282 42724
rect 91649 42721 91661 42724
rect 91695 42721 91707 42755
rect 91649 42715 91707 42721
rect 21542 42644 21548 42696
rect 21600 42684 21606 42696
rect 72510 42684 72516 42696
rect 21600 42656 45554 42684
rect 72471 42656 72516 42684
rect 21600 42644 21606 42656
rect 45526 42548 45554 42656
rect 72510 42644 72516 42656
rect 72568 42644 72574 42696
rect 73062 42684 73068 42696
rect 73023 42656 73068 42684
rect 73062 42644 73068 42656
rect 73120 42644 73126 42696
rect 73172 42656 77294 42684
rect 55950 42576 55956 42628
rect 56008 42616 56014 42628
rect 73172 42616 73200 42656
rect 56008 42588 73200 42616
rect 56008 42576 56014 42588
rect 62206 42548 62212 42560
rect 45526 42520 62212 42548
rect 62206 42508 62212 42520
rect 62264 42548 62270 42560
rect 73522 42548 73528 42560
rect 62264 42520 73528 42548
rect 62264 42508 62270 42520
rect 73522 42508 73528 42520
rect 73580 42508 73586 42560
rect 77266 42548 77294 42656
rect 80698 42616 80704 42628
rect 80659 42588 80704 42616
rect 80698 42576 80704 42588
rect 80756 42576 80762 42628
rect 91833 42619 91891 42625
rect 91833 42585 91845 42619
rect 91879 42616 91891 42619
rect 91922 42616 91928 42628
rect 91879 42588 91928 42616
rect 91879 42585 91891 42588
rect 91833 42579 91891 42585
rect 91922 42576 91928 42588
rect 91980 42576 91986 42628
rect 86586 42548 86592 42560
rect 77266 42520 86592 42548
rect 86586 42508 86592 42520
rect 86644 42548 86650 42560
rect 86862 42548 86868 42560
rect 86644 42520 86868 42548
rect 86644 42508 86650 42520
rect 86862 42508 86868 42520
rect 86920 42508 86926 42560
rect 1104 42458 98808 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 65686 42458
rect 65738 42406 65750 42458
rect 65802 42406 65814 42458
rect 65866 42406 65878 42458
rect 65930 42406 96406 42458
rect 96458 42406 96470 42458
rect 96522 42406 96534 42458
rect 96586 42406 96598 42458
rect 96650 42406 98808 42458
rect 1104 42384 98808 42406
rect 72510 42304 72516 42356
rect 72568 42344 72574 42356
rect 72878 42344 72884 42356
rect 72568 42316 72884 42344
rect 72568 42304 72574 42316
rect 72878 42304 72884 42316
rect 72936 42304 72942 42356
rect 95694 42236 95700 42288
rect 95752 42276 95758 42288
rect 96522 42276 96528 42288
rect 95752 42248 96528 42276
rect 95752 42236 95758 42248
rect 96522 42236 96528 42248
rect 96580 42236 96586 42288
rect 39758 42168 39764 42220
rect 39816 42208 39822 42220
rect 92842 42208 92848 42220
rect 39816 42180 45554 42208
rect 92803 42180 92848 42208
rect 39816 42168 39822 42180
rect 16942 42100 16948 42152
rect 17000 42140 17006 42152
rect 42794 42140 42800 42152
rect 17000 42112 42800 42140
rect 17000 42100 17006 42112
rect 42794 42100 42800 42112
rect 42852 42100 42858 42152
rect 44729 42143 44787 42149
rect 44729 42109 44741 42143
rect 44775 42109 44787 42143
rect 44729 42103 44787 42109
rect 16206 42032 16212 42084
rect 16264 42072 16270 42084
rect 21542 42072 21548 42084
rect 16264 42044 21548 42072
rect 16264 42032 16270 42044
rect 21542 42032 21548 42044
rect 21600 42032 21606 42084
rect 44358 42004 44364 42016
rect 44319 41976 44364 42004
rect 44358 41964 44364 41976
rect 44416 42004 44422 42016
rect 44744 42004 44772 42103
rect 45526 42072 45554 42180
rect 92842 42168 92848 42180
rect 92900 42168 92906 42220
rect 92566 42140 92572 42152
rect 92527 42112 92572 42140
rect 92566 42100 92572 42112
rect 92624 42100 92630 42152
rect 78674 42072 78680 42084
rect 45526 42044 78680 42072
rect 78674 42032 78680 42044
rect 78732 42032 78738 42084
rect 44416 41976 44772 42004
rect 44416 41964 44422 41976
rect 1104 41914 98808 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 50326 41914
rect 50378 41862 50390 41914
rect 50442 41862 50454 41914
rect 50506 41862 50518 41914
rect 50570 41862 81046 41914
rect 81098 41862 81110 41914
rect 81162 41862 81174 41914
rect 81226 41862 81238 41914
rect 81290 41862 98808 41914
rect 1104 41840 98808 41862
rect 80054 41760 80060 41812
rect 80112 41800 80118 41812
rect 80422 41800 80428 41812
rect 80112 41772 80428 41800
rect 80112 41760 80118 41772
rect 80422 41760 80428 41772
rect 80480 41800 80486 41812
rect 80480 41772 97304 41800
rect 80480 41760 80486 41772
rect 42794 41692 42800 41744
rect 42852 41732 42858 41744
rect 42978 41732 42984 41744
rect 42852 41704 42984 41732
rect 42852 41692 42858 41704
rect 42978 41692 42984 41704
rect 43036 41732 43042 41744
rect 72510 41732 72516 41744
rect 43036 41704 72516 41732
rect 43036 41692 43042 41704
rect 72510 41692 72516 41704
rect 72568 41692 72574 41744
rect 86862 41692 86868 41744
rect 86920 41732 86926 41744
rect 86920 41704 97120 41732
rect 86920 41692 86926 41704
rect 29270 41624 29276 41676
rect 29328 41664 29334 41676
rect 30469 41667 30527 41673
rect 30469 41664 30481 41667
rect 29328 41636 30481 41664
rect 29328 41624 29334 41636
rect 30469 41633 30481 41636
rect 30515 41633 30527 41667
rect 30469 41627 30527 41633
rect 48777 41667 48835 41673
rect 48777 41633 48789 41667
rect 48823 41664 48835 41667
rect 95510 41664 95516 41676
rect 48823 41636 95516 41664
rect 48823 41633 48835 41636
rect 48777 41627 48835 41633
rect 95510 41624 95516 41636
rect 95568 41664 95574 41676
rect 97092 41673 97120 41704
rect 97276 41673 97304 41772
rect 96341 41667 96399 41673
rect 96341 41664 96353 41667
rect 95568 41636 96353 41664
rect 95568 41624 95574 41636
rect 96341 41633 96353 41636
rect 96387 41633 96399 41667
rect 96709 41667 96767 41673
rect 96709 41664 96721 41667
rect 96341 41627 96399 41633
rect 96448 41636 96721 41664
rect 31294 41596 31300 41608
rect 31255 41568 31300 41596
rect 31294 41556 31300 41568
rect 31352 41556 31358 41608
rect 49418 41596 49424 41608
rect 49379 41568 49424 41596
rect 49418 41556 49424 41568
rect 49476 41556 49482 41608
rect 96154 41596 96160 41608
rect 96115 41568 96160 41596
rect 96154 41556 96160 41568
rect 96212 41596 96218 41608
rect 96448 41596 96476 41636
rect 96709 41633 96721 41636
rect 96755 41633 96767 41667
rect 96709 41627 96767 41633
rect 97077 41667 97135 41673
rect 97077 41633 97089 41667
rect 97123 41633 97135 41667
rect 97077 41627 97135 41633
rect 97261 41667 97319 41673
rect 97261 41633 97273 41667
rect 97307 41633 97319 41667
rect 97261 41627 97319 41633
rect 96212 41568 96476 41596
rect 96212 41556 96218 41568
rect 96522 41556 96528 41608
rect 96580 41596 96586 41608
rect 96580 41568 96625 41596
rect 96580 41556 96586 41568
rect 18138 41488 18144 41540
rect 18196 41528 18202 41540
rect 97445 41531 97503 41537
rect 97445 41528 97457 41531
rect 18196 41500 97457 41528
rect 18196 41488 18202 41500
rect 97445 41497 97457 41500
rect 97491 41497 97503 41531
rect 97445 41491 97503 41497
rect 18782 41420 18788 41472
rect 18840 41460 18846 41472
rect 80054 41460 80060 41472
rect 18840 41432 80060 41460
rect 18840 41420 18846 41432
rect 80054 41420 80060 41432
rect 80112 41420 80118 41472
rect 1104 41370 98808 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 65686 41370
rect 65738 41318 65750 41370
rect 65802 41318 65814 41370
rect 65866 41318 65878 41370
rect 65930 41318 96406 41370
rect 96458 41318 96470 41370
rect 96522 41318 96534 41370
rect 96586 41318 96598 41370
rect 96650 41318 98808 41370
rect 1104 41296 98808 41318
rect 12342 41216 12348 41268
rect 12400 41256 12406 41268
rect 24854 41256 24860 41268
rect 12400 41228 24860 41256
rect 12400 41216 12406 41228
rect 24854 41216 24860 41228
rect 24912 41216 24918 41268
rect 44266 41216 44272 41268
rect 44324 41256 44330 41268
rect 66898 41256 66904 41268
rect 44324 41228 66904 41256
rect 44324 41216 44330 41228
rect 66898 41216 66904 41228
rect 66956 41216 66962 41268
rect 25590 41148 25596 41200
rect 25648 41188 25654 41200
rect 34422 41188 34428 41200
rect 25648 41160 34428 41188
rect 25648 41148 25654 41160
rect 34422 41148 34428 41160
rect 34480 41148 34486 41200
rect 44634 41148 44640 41200
rect 44692 41188 44698 41200
rect 48130 41188 48136 41200
rect 44692 41160 48136 41188
rect 44692 41148 44698 41160
rect 48130 41148 48136 41160
rect 48188 41148 48194 41200
rect 14366 41080 14372 41132
rect 14424 41120 14430 41132
rect 26970 41120 26976 41132
rect 14424 41092 26976 41120
rect 14424 41080 14430 41092
rect 26970 41080 26976 41092
rect 27028 41080 27034 41132
rect 8294 41012 8300 41064
rect 8352 41052 8358 41064
rect 36538 41052 36544 41064
rect 8352 41024 36544 41052
rect 8352 41012 8358 41024
rect 36538 41012 36544 41024
rect 36596 41012 36602 41064
rect 14826 40944 14832 40996
rect 14884 40984 14890 40996
rect 42518 40984 42524 40996
rect 14884 40956 42524 40984
rect 14884 40944 14890 40956
rect 42518 40944 42524 40956
rect 42576 40944 42582 40996
rect 86862 40944 86868 40996
rect 86920 40984 86926 40996
rect 92106 40984 92112 40996
rect 86920 40956 92112 40984
rect 86920 40944 86926 40956
rect 92106 40944 92112 40956
rect 92164 40944 92170 40996
rect 11882 40876 11888 40928
rect 11940 40916 11946 40928
rect 12342 40916 12348 40928
rect 11940 40888 12348 40916
rect 11940 40876 11946 40888
rect 12342 40876 12348 40888
rect 12400 40876 12406 40928
rect 24854 40876 24860 40928
rect 24912 40916 24918 40928
rect 53742 40916 53748 40928
rect 24912 40888 53748 40916
rect 24912 40876 24918 40888
rect 53742 40876 53748 40888
rect 53800 40876 53806 40928
rect 66898 40876 66904 40928
rect 66956 40916 66962 40928
rect 88426 40916 88432 40928
rect 66956 40888 88432 40916
rect 66956 40876 66962 40888
rect 88426 40876 88432 40888
rect 88484 40876 88490 40928
rect 1104 40826 98808 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 50326 40826
rect 50378 40774 50390 40826
rect 50442 40774 50454 40826
rect 50506 40774 50518 40826
rect 50570 40774 81046 40826
rect 81098 40774 81110 40826
rect 81162 40774 81174 40826
rect 81226 40774 81238 40826
rect 81290 40774 98808 40826
rect 1104 40752 98808 40774
rect 19978 40672 19984 40724
rect 20036 40712 20042 40724
rect 68554 40712 68560 40724
rect 20036 40684 68560 40712
rect 20036 40672 20042 40684
rect 68554 40672 68560 40684
rect 68612 40672 68618 40724
rect 86402 40712 86408 40724
rect 70366 40684 86408 40712
rect 31754 40536 31760 40588
rect 31812 40576 31818 40588
rect 32398 40576 32404 40588
rect 31812 40548 32404 40576
rect 31812 40536 31818 40548
rect 32398 40536 32404 40548
rect 32456 40576 32462 40588
rect 70366 40576 70394 40684
rect 86402 40672 86408 40684
rect 86460 40712 86466 40724
rect 86862 40712 86868 40724
rect 86460 40684 86868 40712
rect 86460 40672 86466 40684
rect 86862 40672 86868 40684
rect 86920 40672 86926 40724
rect 90542 40712 90548 40724
rect 90503 40684 90548 40712
rect 90542 40672 90548 40684
rect 90600 40672 90606 40724
rect 95510 40712 95516 40724
rect 95471 40684 95516 40712
rect 95510 40672 95516 40684
rect 95568 40672 95574 40724
rect 32456 40548 70394 40576
rect 90560 40576 90588 40672
rect 92109 40579 92167 40585
rect 92109 40576 92121 40579
rect 90560 40548 92121 40576
rect 32456 40536 32462 40548
rect 92109 40545 92121 40548
rect 92155 40545 92167 40579
rect 95421 40579 95479 40585
rect 95421 40576 95433 40579
rect 92109 40539 92167 40545
rect 92216 40548 95433 40576
rect 36354 40468 36360 40520
rect 36412 40508 36418 40520
rect 36538 40508 36544 40520
rect 36412 40480 36544 40508
rect 36412 40468 36418 40480
rect 36538 40468 36544 40480
rect 36596 40508 36602 40520
rect 67726 40508 67732 40520
rect 36596 40480 67732 40508
rect 36596 40468 36602 40480
rect 67726 40468 67732 40480
rect 67784 40468 67790 40520
rect 68554 40468 68560 40520
rect 68612 40508 68618 40520
rect 68922 40508 68928 40520
rect 68612 40480 68928 40508
rect 68612 40468 68618 40480
rect 68922 40468 68928 40480
rect 68980 40468 68986 40520
rect 74074 40508 74080 40520
rect 70366 40480 74080 40508
rect 34422 40400 34428 40452
rect 34480 40440 34486 40452
rect 70366 40440 70394 40480
rect 74074 40468 74080 40480
rect 74132 40468 74138 40520
rect 92014 40468 92020 40520
rect 92072 40508 92078 40520
rect 92216 40508 92244 40548
rect 95421 40545 95433 40548
rect 95467 40545 95479 40579
rect 95421 40539 95479 40545
rect 92382 40508 92388 40520
rect 92072 40480 92244 40508
rect 92343 40480 92388 40508
rect 92072 40468 92078 40480
rect 92382 40468 92388 40480
rect 92440 40468 92446 40520
rect 90821 40443 90879 40449
rect 90821 40440 90833 40443
rect 34480 40412 70394 40440
rect 71240 40412 90833 40440
rect 34480 40400 34486 40412
rect 66162 40332 66168 40384
rect 66220 40372 66226 40384
rect 71240 40372 71268 40412
rect 90821 40409 90833 40412
rect 90867 40409 90879 40443
rect 90821 40403 90879 40409
rect 77662 40372 77668 40384
rect 66220 40344 71268 40372
rect 77623 40344 77668 40372
rect 66220 40332 66226 40344
rect 77662 40332 77668 40344
rect 77720 40372 77726 40384
rect 77849 40375 77907 40381
rect 77849 40372 77861 40375
rect 77720 40344 77861 40372
rect 77720 40332 77726 40344
rect 77849 40341 77861 40344
rect 77895 40341 77907 40375
rect 77849 40335 77907 40341
rect 1104 40282 98808 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 65686 40282
rect 65738 40230 65750 40282
rect 65802 40230 65814 40282
rect 65866 40230 65878 40282
rect 65930 40230 96406 40282
rect 96458 40230 96470 40282
rect 96522 40230 96534 40282
rect 96586 40230 96598 40282
rect 96650 40230 98808 40282
rect 1104 40208 98808 40230
rect 53650 40128 53656 40180
rect 53708 40168 53714 40180
rect 77662 40168 77668 40180
rect 53708 40140 77668 40168
rect 53708 40128 53714 40140
rect 77662 40128 77668 40140
rect 77720 40128 77726 40180
rect 32953 40103 33011 40109
rect 32953 40069 32965 40103
rect 32999 40100 33011 40103
rect 33229 40103 33287 40109
rect 33229 40100 33241 40103
rect 32999 40072 33241 40100
rect 32999 40069 33011 40072
rect 32953 40063 33011 40069
rect 33229 40069 33241 40072
rect 33275 40100 33287 40103
rect 34238 40100 34244 40112
rect 33275 40072 34244 40100
rect 33275 40069 33287 40072
rect 33229 40063 33287 40069
rect 34238 40060 34244 40072
rect 34296 40060 34302 40112
rect 35802 40060 35808 40112
rect 35860 40100 35866 40112
rect 39758 40100 39764 40112
rect 35860 40072 39764 40100
rect 35860 40060 35866 40072
rect 39758 40060 39764 40072
rect 39816 40060 39822 40112
rect 43806 40060 43812 40112
rect 43864 40100 43870 40112
rect 44818 40100 44824 40112
rect 43864 40072 44824 40100
rect 43864 40060 43870 40072
rect 44818 40060 44824 40072
rect 44876 40060 44882 40112
rect 47026 40060 47032 40112
rect 47084 40100 47090 40112
rect 48958 40100 48964 40112
rect 47084 40072 48964 40100
rect 47084 40060 47090 40072
rect 48958 40060 48964 40072
rect 49016 40060 49022 40112
rect 67726 40060 67732 40112
rect 67784 40100 67790 40112
rect 68646 40100 68652 40112
rect 67784 40072 68652 40100
rect 67784 40060 67790 40072
rect 68646 40060 68652 40072
rect 68704 40060 68710 40112
rect 12986 39992 12992 40044
rect 13044 40032 13050 40044
rect 14642 40032 14648 40044
rect 13044 40004 14648 40032
rect 13044 39992 13050 40004
rect 14642 39992 14648 40004
rect 14700 39992 14706 40044
rect 41056 40035 41114 40041
rect 14752 40004 40264 40032
rect 2777 39967 2835 39973
rect 2777 39933 2789 39967
rect 2823 39933 2835 39967
rect 2777 39927 2835 39933
rect 2792 39828 2820 39927
rect 10870 39924 10876 39976
rect 10928 39964 10934 39976
rect 14752 39964 14780 40004
rect 18966 39964 18972 39976
rect 10928 39936 14780 39964
rect 16546 39936 18972 39964
rect 10928 39924 10934 39936
rect 3329 39899 3387 39905
rect 3329 39865 3341 39899
rect 3375 39896 3387 39899
rect 7742 39896 7748 39908
rect 3375 39868 7748 39896
rect 3375 39865 3387 39868
rect 3329 39859 3387 39865
rect 7742 39856 7748 39868
rect 7800 39856 7806 39908
rect 10042 39856 10048 39908
rect 10100 39896 10106 39908
rect 16546 39896 16574 39936
rect 18966 39924 18972 39936
rect 19024 39924 19030 39976
rect 28353 39967 28411 39973
rect 28353 39933 28365 39967
rect 28399 39933 28411 39967
rect 28353 39927 28411 39933
rect 28629 39967 28687 39973
rect 28629 39933 28641 39967
rect 28675 39964 28687 39967
rect 28718 39964 28724 39976
rect 28675 39936 28724 39964
rect 28675 39933 28687 39936
rect 28629 39927 28687 39933
rect 10100 39868 16574 39896
rect 10100 39856 10106 39868
rect 28258 39828 28264 39840
rect 2792 39800 28264 39828
rect 28258 39788 28264 39800
rect 28316 39788 28322 39840
rect 28368 39828 28396 39927
rect 28718 39924 28724 39936
rect 28776 39924 28782 39976
rect 34422 39964 34428 39976
rect 34383 39936 34428 39964
rect 34422 39924 34428 39936
rect 34480 39924 34486 39976
rect 34606 39964 34612 39976
rect 34567 39936 34612 39964
rect 34606 39924 34612 39936
rect 34664 39924 34670 39976
rect 34845 39967 34903 39973
rect 34845 39933 34857 39967
rect 34891 39964 34903 39967
rect 35250 39964 35256 39976
rect 34891 39936 35256 39964
rect 34891 39933 34903 39936
rect 34845 39927 34903 39933
rect 35250 39924 35256 39936
rect 35308 39924 35314 39976
rect 40236 39964 40264 40004
rect 41056 40001 41068 40035
rect 41102 40001 41114 40035
rect 41056 39995 41114 40001
rect 41509 40035 41567 40041
rect 41509 40001 41521 40035
rect 41555 40032 41567 40035
rect 49694 40032 49700 40044
rect 41555 40004 49700 40032
rect 41555 40001 41567 40004
rect 41509 39995 41567 40001
rect 40770 39964 40776 39976
rect 40236 39936 40776 39964
rect 40770 39924 40776 39936
rect 40828 39924 40834 39976
rect 40956 39967 41014 39973
rect 40956 39933 40968 39967
rect 41002 39933 41014 39967
rect 40956 39927 41014 39933
rect 31018 39896 31024 39908
rect 29288 39868 31024 39896
rect 29288 39828 29316 39868
rect 31018 39856 31024 39868
rect 31076 39856 31082 39908
rect 34698 39896 34704 39908
rect 34659 39868 34704 39896
rect 34698 39856 34704 39868
rect 34756 39856 34762 39908
rect 40972 39896 41000 39927
rect 41064 39908 41092 39995
rect 49694 39992 49700 40004
rect 49752 39992 49758 40044
rect 50062 40032 50068 40044
rect 50023 40004 50068 40032
rect 50062 39992 50068 40004
rect 50120 39992 50126 40044
rect 50249 40035 50307 40041
rect 50249 40001 50261 40035
rect 50295 40032 50307 40035
rect 59265 40035 59323 40041
rect 59265 40032 59277 40035
rect 50295 40004 59277 40032
rect 50295 40001 50307 40004
rect 50249 39995 50307 40001
rect 59265 40001 59277 40004
rect 59311 40032 59323 40035
rect 60918 40032 60924 40044
rect 59311 40004 60734 40032
rect 60879 40004 60924 40032
rect 59311 40001 59323 40004
rect 59265 39995 59323 40001
rect 41141 39967 41199 39973
rect 41141 39933 41153 39967
rect 41187 39933 41199 39967
rect 41141 39927 41199 39933
rect 41325 39967 41383 39973
rect 41325 39933 41337 39967
rect 41371 39964 41383 39967
rect 41598 39964 41604 39976
rect 41371 39936 41604 39964
rect 41371 39933 41383 39936
rect 41325 39927 41383 39933
rect 40604 39868 41000 39896
rect 40604 39840 40632 39868
rect 41046 39856 41052 39908
rect 41104 39856 41110 39908
rect 29730 39828 29736 39840
rect 28368 39800 29316 39828
rect 29691 39800 29736 39828
rect 29730 39788 29736 39800
rect 29788 39788 29794 39840
rect 32858 39788 32864 39840
rect 32916 39828 32922 39840
rect 34054 39828 34060 39840
rect 32916 39800 34060 39828
rect 32916 39788 32922 39800
rect 34054 39788 34060 39800
rect 34112 39788 34118 39840
rect 34790 39788 34796 39840
rect 34848 39828 34854 39840
rect 34985 39831 35043 39837
rect 34985 39828 34997 39831
rect 34848 39800 34997 39828
rect 34848 39788 34854 39800
rect 34985 39797 34997 39800
rect 35031 39797 35043 39831
rect 40586 39828 40592 39840
rect 40547 39800 40592 39828
rect 34985 39791 35043 39797
rect 40586 39788 40592 39800
rect 40644 39788 40650 39840
rect 41156 39828 41184 39927
rect 41598 39924 41604 39936
rect 41656 39924 41662 39976
rect 44818 39924 44824 39976
rect 44876 39964 44882 39976
rect 45186 39964 45192 39976
rect 44876 39936 45192 39964
rect 44876 39924 44882 39936
rect 45186 39924 45192 39936
rect 45244 39924 45250 39976
rect 50080 39964 50108 39992
rect 50525 39967 50583 39973
rect 50525 39964 50537 39967
rect 50080 39936 50537 39964
rect 50525 39933 50537 39936
rect 50571 39933 50583 39967
rect 50525 39927 50583 39933
rect 57330 39924 57336 39976
rect 57388 39964 57394 39976
rect 59081 39967 59139 39973
rect 59081 39964 59093 39967
rect 57388 39936 59093 39964
rect 57388 39924 57394 39936
rect 59081 39933 59093 39936
rect 59127 39964 59139 39967
rect 59541 39967 59599 39973
rect 59541 39964 59553 39967
rect 59127 39936 59553 39964
rect 59127 39933 59139 39936
rect 59081 39927 59139 39933
rect 59541 39933 59553 39936
rect 59587 39933 59599 39967
rect 60706 39964 60734 40004
rect 60918 39992 60924 40004
rect 60976 39992 60982 40044
rect 71777 40035 71835 40041
rect 71777 40001 71789 40035
rect 71823 40032 71835 40035
rect 73614 40032 73620 40044
rect 71823 40004 73620 40032
rect 71823 40001 71835 40004
rect 71777 39995 71835 40001
rect 73614 39992 73620 40004
rect 73672 39992 73678 40044
rect 61562 39964 61568 39976
rect 60706 39936 61568 39964
rect 59541 39927 59599 39933
rect 61562 39924 61568 39936
rect 61620 39924 61626 39976
rect 67729 39967 67787 39973
rect 67729 39933 67741 39967
rect 67775 39964 67787 39967
rect 68005 39967 68063 39973
rect 68005 39964 68017 39967
rect 67775 39936 68017 39964
rect 67775 39933 67787 39936
rect 67729 39927 67787 39933
rect 68005 39933 68017 39936
rect 68051 39964 68063 39967
rect 71498 39964 71504 39976
rect 68051 39936 71504 39964
rect 68051 39933 68063 39936
rect 68005 39927 68063 39933
rect 71498 39924 71504 39936
rect 71556 39924 71562 39976
rect 72050 39964 72056 39976
rect 72011 39936 72056 39964
rect 72050 39924 72056 39936
rect 72108 39924 72114 39976
rect 41230 39856 41236 39908
rect 41288 39896 41294 39908
rect 73338 39896 73344 39908
rect 41288 39868 50200 39896
rect 41288 39856 41294 39868
rect 44818 39828 44824 39840
rect 41156 39800 44824 39828
rect 44818 39788 44824 39800
rect 44876 39788 44882 39840
rect 50172 39828 50200 39868
rect 72988 39868 73344 39896
rect 51629 39831 51687 39837
rect 51629 39828 51641 39831
rect 50172 39800 51641 39828
rect 51629 39797 51641 39800
rect 51675 39797 51687 39831
rect 51629 39791 51687 39797
rect 64046 39788 64052 39840
rect 64104 39828 64110 39840
rect 72988 39828 73016 39868
rect 73338 39856 73344 39868
rect 73396 39856 73402 39908
rect 73154 39828 73160 39840
rect 64104 39800 73016 39828
rect 73115 39800 73160 39828
rect 64104 39788 64110 39800
rect 73154 39788 73160 39800
rect 73212 39788 73218 39840
rect 1104 39738 98808 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 50326 39738
rect 50378 39686 50390 39738
rect 50442 39686 50454 39738
rect 50506 39686 50518 39738
rect 50570 39686 81046 39738
rect 81098 39686 81110 39738
rect 81162 39686 81174 39738
rect 81226 39686 81238 39738
rect 81290 39686 98808 39738
rect 1104 39664 98808 39686
rect 6178 39624 6184 39636
rect 6139 39596 6184 39624
rect 6178 39584 6184 39596
rect 6236 39584 6242 39636
rect 28258 39584 28264 39636
rect 28316 39624 28322 39636
rect 31110 39624 31116 39636
rect 28316 39596 31116 39624
rect 28316 39584 28322 39596
rect 31110 39584 31116 39596
rect 31168 39584 31174 39636
rect 33137 39627 33195 39633
rect 33137 39593 33149 39627
rect 33183 39624 33195 39627
rect 33321 39627 33379 39633
rect 33321 39624 33333 39627
rect 33183 39596 33333 39624
rect 33183 39593 33195 39596
rect 33137 39587 33195 39593
rect 33321 39593 33333 39596
rect 33367 39624 33379 39627
rect 33686 39624 33692 39636
rect 33367 39596 33692 39624
rect 33367 39593 33379 39596
rect 33321 39587 33379 39593
rect 33686 39584 33692 39596
rect 33744 39584 33750 39636
rect 34146 39624 34152 39636
rect 34107 39596 34152 39624
rect 34146 39584 34152 39596
rect 34204 39584 34210 39636
rect 40770 39584 40776 39636
rect 40828 39624 40834 39636
rect 42058 39624 42064 39636
rect 40828 39596 42064 39624
rect 40828 39584 40834 39596
rect 42058 39584 42064 39596
rect 42116 39584 42122 39636
rect 49694 39584 49700 39636
rect 49752 39624 49758 39636
rect 50982 39624 50988 39636
rect 49752 39596 50988 39624
rect 49752 39584 49758 39596
rect 50982 39584 50988 39596
rect 51040 39584 51046 39636
rect 70026 39584 70032 39636
rect 70084 39624 70090 39636
rect 76834 39624 76840 39636
rect 70084 39596 76840 39624
rect 70084 39584 70090 39596
rect 76834 39584 76840 39596
rect 76892 39584 76898 39636
rect 31665 39559 31723 39565
rect 31665 39525 31677 39559
rect 31711 39556 31723 39559
rect 31711 39528 33824 39556
rect 31711 39525 31723 39528
rect 31665 39519 31723 39525
rect 5074 39488 5080 39500
rect 5035 39460 5080 39488
rect 5074 39448 5080 39460
rect 5132 39448 5138 39500
rect 29546 39448 29552 39500
rect 29604 39488 29610 39500
rect 31113 39491 31171 39497
rect 31113 39488 31125 39491
rect 29604 39460 31125 39488
rect 29604 39448 29610 39460
rect 31113 39457 31125 39460
rect 31159 39488 31171 39491
rect 31570 39488 31576 39500
rect 31159 39460 31576 39488
rect 31159 39457 31171 39460
rect 31113 39451 31171 39457
rect 31570 39448 31576 39460
rect 31628 39448 31634 39500
rect 32125 39491 32183 39497
rect 32125 39457 32137 39491
rect 32171 39488 32183 39491
rect 32677 39491 32735 39497
rect 32677 39488 32689 39491
rect 32171 39460 32689 39488
rect 32171 39457 32183 39460
rect 32125 39451 32183 39457
rect 32677 39457 32689 39460
rect 32723 39457 32735 39491
rect 32950 39488 32956 39500
rect 32911 39460 32956 39488
rect 32677 39451 32735 39457
rect 4801 39423 4859 39429
rect 4801 39389 4813 39423
rect 4847 39420 4859 39423
rect 6086 39420 6092 39432
rect 4847 39392 6092 39420
rect 4847 39389 4859 39392
rect 4801 39383 4859 39389
rect 6086 39380 6092 39392
rect 6144 39380 6150 39432
rect 32490 39420 32496 39432
rect 32451 39392 32496 39420
rect 32490 39380 32496 39392
rect 32548 39380 32554 39432
rect 32692 39420 32720 39451
rect 32950 39448 32956 39460
rect 33008 39448 33014 39500
rect 33413 39491 33471 39497
rect 33413 39457 33425 39491
rect 33459 39457 33471 39491
rect 33594 39488 33600 39500
rect 33555 39460 33600 39488
rect 33413 39451 33471 39457
rect 33428 39420 33456 39451
rect 33594 39448 33600 39460
rect 33652 39448 33658 39500
rect 33502 39420 33508 39432
rect 32692 39392 33272 39420
rect 33428 39392 33508 39420
rect 32858 39352 32864 39364
rect 32819 39324 32864 39352
rect 32858 39312 32864 39324
rect 32916 39312 32922 39364
rect 24210 39244 24216 39296
rect 24268 39284 24274 39296
rect 33137 39287 33195 39293
rect 33137 39284 33149 39287
rect 24268 39256 33149 39284
rect 24268 39244 24274 39256
rect 33137 39253 33149 39256
rect 33183 39253 33195 39287
rect 33244 39284 33272 39392
rect 33502 39380 33508 39392
rect 33560 39380 33566 39432
rect 33686 39420 33692 39432
rect 33647 39392 33692 39420
rect 33686 39380 33692 39392
rect 33744 39380 33750 39432
rect 33796 39429 33824 39528
rect 34054 39516 34060 39568
rect 34112 39556 34118 39568
rect 44266 39556 44272 39568
rect 34112 39528 44272 39556
rect 34112 39516 34118 39528
rect 44266 39516 44272 39528
rect 44324 39516 44330 39568
rect 53742 39516 53748 39568
rect 53800 39556 53806 39568
rect 78306 39556 78312 39568
rect 53800 39528 78312 39556
rect 53800 39516 53806 39528
rect 78306 39516 78312 39528
rect 78364 39516 78370 39568
rect 33962 39488 33968 39500
rect 33923 39460 33968 39488
rect 33962 39448 33968 39460
rect 34020 39448 34026 39500
rect 34698 39448 34704 39500
rect 34756 39488 34762 39500
rect 44910 39488 44916 39500
rect 34756 39460 44916 39488
rect 34756 39448 34762 39460
rect 44910 39448 44916 39460
rect 44968 39488 44974 39500
rect 55490 39488 55496 39500
rect 44968 39460 55496 39488
rect 44968 39448 44974 39460
rect 55490 39448 55496 39460
rect 55548 39448 55554 39500
rect 69014 39488 69020 39500
rect 68975 39460 69020 39488
rect 69014 39448 69020 39460
rect 69072 39448 69078 39500
rect 33781 39423 33839 39429
rect 33781 39389 33793 39423
rect 33827 39420 33839 39423
rect 63402 39420 63408 39432
rect 33827 39392 63408 39420
rect 33827 39389 33839 39392
rect 33781 39383 33839 39389
rect 63402 39380 63408 39392
rect 63460 39420 63466 39432
rect 97442 39420 97448 39432
rect 63460 39392 97448 39420
rect 63460 39380 63466 39392
rect 97442 39380 97448 39392
rect 97500 39380 97506 39432
rect 33612 39324 41414 39352
rect 33612 39284 33640 39324
rect 33244 39256 33640 39284
rect 33137 39247 33195 39253
rect 35710 39244 35716 39296
rect 35768 39284 35774 39296
rect 41230 39284 41236 39296
rect 35768 39256 41236 39284
rect 35768 39244 35774 39256
rect 41230 39244 41236 39256
rect 41288 39244 41294 39296
rect 41386 39284 41414 39324
rect 69198 39312 69204 39364
rect 69256 39352 69262 39364
rect 78398 39352 78404 39364
rect 69256 39324 78404 39352
rect 69256 39312 69262 39324
rect 78398 39312 78404 39324
rect 78456 39312 78462 39364
rect 66990 39284 66996 39296
rect 41386 39256 66996 39284
rect 66990 39244 66996 39256
rect 67048 39244 67054 39296
rect 68922 39284 68928 39296
rect 68883 39256 68928 39284
rect 68922 39244 68928 39256
rect 68980 39244 68986 39296
rect 1104 39194 98808 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 65686 39194
rect 65738 39142 65750 39194
rect 65802 39142 65814 39194
rect 65866 39142 65878 39194
rect 65930 39142 96406 39194
rect 96458 39142 96470 39194
rect 96522 39142 96534 39194
rect 96586 39142 96598 39194
rect 96650 39142 98808 39194
rect 1104 39120 98808 39142
rect 33502 39040 33508 39092
rect 33560 39080 33566 39092
rect 34514 39080 34520 39092
rect 33560 39052 34520 39080
rect 33560 39040 33566 39052
rect 34514 39040 34520 39052
rect 34572 39080 34578 39092
rect 35526 39080 35532 39092
rect 34572 39052 35532 39080
rect 34572 39040 34578 39052
rect 35526 39040 35532 39052
rect 35584 39040 35590 39092
rect 40034 39040 40040 39092
rect 40092 39080 40098 39092
rect 41138 39080 41144 39092
rect 40092 39052 41144 39080
rect 40092 39040 40098 39052
rect 41138 39040 41144 39052
rect 41196 39080 41202 39092
rect 68922 39080 68928 39092
rect 41196 39052 68928 39080
rect 41196 39040 41202 39052
rect 68922 39040 68928 39052
rect 68980 39040 68986 39092
rect 7558 38972 7564 39024
rect 7616 39012 7622 39024
rect 40586 39012 40592 39024
rect 7616 38984 40592 39012
rect 7616 38972 7622 38984
rect 40586 38972 40592 38984
rect 40644 38972 40650 39024
rect 60366 38972 60372 39024
rect 60424 39012 60430 39024
rect 73154 39012 73160 39024
rect 60424 38984 73160 39012
rect 60424 38972 60430 38984
rect 73154 38972 73160 38984
rect 73212 38972 73218 39024
rect 18230 38904 18236 38956
rect 18288 38944 18294 38956
rect 18966 38944 18972 38956
rect 18288 38916 18972 38944
rect 18288 38904 18294 38916
rect 18966 38904 18972 38916
rect 19024 38944 19030 38956
rect 33594 38944 33600 38956
rect 19024 38916 33600 38944
rect 19024 38904 19030 38916
rect 33594 38904 33600 38916
rect 33652 38904 33658 38956
rect 33042 38808 33048 38820
rect 33003 38780 33048 38808
rect 33042 38768 33048 38780
rect 33100 38768 33106 38820
rect 33873 38811 33931 38817
rect 33873 38777 33885 38811
rect 33919 38808 33931 38811
rect 43530 38808 43536 38820
rect 33919 38780 43536 38808
rect 33919 38777 33931 38780
rect 33873 38771 33931 38777
rect 43530 38768 43536 38780
rect 43588 38768 43594 38820
rect 1104 38650 98808 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 50326 38650
rect 50378 38598 50390 38650
rect 50442 38598 50454 38650
rect 50506 38598 50518 38650
rect 50570 38598 81046 38650
rect 81098 38598 81110 38650
rect 81162 38598 81174 38650
rect 81226 38598 81238 38650
rect 81290 38598 98808 38650
rect 1104 38576 98808 38598
rect 33042 38536 33048 38548
rect 10244 38508 33048 38536
rect 10244 38400 10272 38508
rect 33042 38496 33048 38508
rect 33100 38536 33106 38548
rect 33321 38539 33379 38545
rect 33321 38536 33333 38539
rect 33100 38508 33333 38536
rect 33100 38496 33106 38508
rect 33321 38505 33333 38508
rect 33367 38505 33379 38539
rect 33321 38499 33379 38505
rect 43165 38539 43223 38545
rect 43165 38505 43177 38539
rect 43211 38536 43223 38539
rect 43254 38536 43260 38548
rect 43211 38508 43260 38536
rect 43211 38505 43223 38508
rect 43165 38499 43223 38505
rect 43254 38496 43260 38508
rect 43312 38496 43318 38548
rect 43346 38496 43352 38548
rect 43404 38536 43410 38548
rect 94222 38536 94228 38548
rect 43404 38508 94228 38536
rect 43404 38496 43410 38508
rect 94222 38496 94228 38508
rect 94280 38496 94286 38548
rect 11330 38468 11336 38480
rect 11072 38440 11336 38468
rect 10401 38403 10459 38409
rect 10401 38400 10413 38403
rect 10244 38372 10413 38400
rect 10401 38369 10413 38372
rect 10447 38369 10459 38403
rect 10401 38363 10459 38369
rect 10689 38403 10747 38409
rect 10689 38369 10701 38403
rect 10735 38369 10747 38403
rect 10689 38363 10747 38369
rect 10781 38403 10839 38409
rect 10781 38369 10793 38403
rect 10827 38400 10839 38403
rect 10962 38400 10968 38412
rect 10827 38372 10968 38400
rect 10827 38369 10839 38372
rect 10781 38363 10839 38369
rect 10502 38292 10508 38344
rect 10560 38332 10566 38344
rect 10704 38332 10732 38363
rect 10962 38360 10968 38372
rect 11020 38360 11026 38412
rect 11072 38409 11100 38440
rect 11330 38428 11336 38440
rect 11388 38428 11394 38480
rect 32677 38471 32735 38477
rect 32677 38437 32689 38471
rect 32723 38468 32735 38471
rect 73249 38471 73307 38477
rect 32723 38440 60734 38468
rect 32723 38437 32735 38440
rect 32677 38431 32735 38437
rect 11057 38403 11115 38409
rect 11057 38369 11069 38403
rect 11103 38369 11115 38403
rect 11057 38363 11115 38369
rect 11241 38403 11299 38409
rect 11241 38369 11253 38403
rect 11287 38400 11299 38403
rect 16022 38400 16028 38412
rect 11287 38372 16028 38400
rect 11287 38369 11299 38372
rect 11241 38363 11299 38369
rect 16022 38360 16028 38372
rect 16080 38360 16086 38412
rect 33229 38403 33287 38409
rect 33229 38369 33241 38403
rect 33275 38400 33287 38403
rect 38102 38400 38108 38412
rect 33275 38372 38108 38400
rect 33275 38369 33287 38372
rect 33229 38363 33287 38369
rect 38102 38360 38108 38372
rect 38160 38360 38166 38412
rect 42518 38400 42524 38412
rect 42479 38372 42524 38400
rect 42518 38360 42524 38372
rect 42576 38360 42582 38412
rect 42704 38403 42762 38409
rect 42704 38369 42716 38403
rect 42750 38369 42762 38403
rect 42886 38400 42892 38412
rect 42847 38372 42892 38400
rect 42704 38363 42762 38369
rect 20162 38332 20168 38344
rect 10560 38304 20168 38332
rect 10560 38292 10566 38304
rect 20162 38292 20168 38304
rect 20220 38292 20226 38344
rect 31018 38332 31024 38344
rect 30979 38304 31024 38332
rect 31018 38292 31024 38304
rect 31076 38292 31082 38344
rect 31297 38335 31355 38341
rect 31297 38301 31309 38335
rect 31343 38332 31355 38335
rect 31478 38332 31484 38344
rect 31343 38304 31484 38332
rect 31343 38301 31355 38304
rect 31297 38295 31355 38301
rect 31478 38292 31484 38304
rect 31536 38292 31542 38344
rect 41322 38292 41328 38344
rect 41380 38332 41386 38344
rect 42720 38332 42748 38363
rect 42886 38360 42892 38372
rect 42944 38360 42950 38412
rect 43070 38400 43076 38412
rect 43031 38372 43076 38400
rect 43070 38360 43076 38372
rect 43128 38360 43134 38412
rect 46385 38403 46443 38409
rect 46385 38400 46397 38403
rect 45526 38372 46397 38400
rect 41380 38304 42748 38332
rect 42804 38335 42862 38341
rect 41380 38292 41386 38304
rect 42804 38301 42816 38335
rect 42850 38332 42862 38335
rect 42978 38332 42984 38344
rect 42850 38304 42984 38332
rect 42850 38301 42862 38304
rect 42804 38295 42862 38301
rect 42978 38292 42984 38304
rect 43036 38292 43042 38344
rect 10045 38267 10103 38273
rect 10045 38233 10057 38267
rect 10091 38264 10103 38267
rect 11238 38264 11244 38276
rect 10091 38236 11244 38264
rect 10091 38233 10103 38236
rect 10045 38227 10103 38233
rect 11238 38224 11244 38236
rect 11296 38224 11302 38276
rect 42518 38224 42524 38276
rect 42576 38264 42582 38276
rect 45526 38264 45554 38372
rect 46385 38369 46397 38372
rect 46431 38400 46443 38403
rect 46750 38400 46756 38412
rect 46431 38372 46756 38400
rect 46431 38369 46443 38372
rect 46385 38363 46443 38369
rect 46750 38360 46756 38372
rect 46808 38360 46814 38412
rect 48130 38400 48136 38412
rect 48091 38372 48136 38400
rect 48130 38360 48136 38372
rect 48188 38360 48194 38412
rect 48498 38360 48504 38412
rect 48556 38400 48562 38412
rect 49602 38400 49608 38412
rect 48556 38372 49608 38400
rect 48556 38360 48562 38372
rect 49602 38360 49608 38372
rect 49660 38360 49666 38412
rect 60706 38400 60734 38440
rect 73249 38437 73261 38471
rect 73295 38468 73307 38471
rect 73338 38468 73344 38480
rect 73295 38440 73344 38468
rect 73295 38437 73307 38440
rect 73249 38431 73307 38437
rect 73338 38428 73344 38440
rect 73396 38428 73402 38480
rect 87598 38468 87604 38480
rect 80026 38440 87604 38468
rect 80026 38400 80054 38440
rect 87598 38428 87604 38440
rect 87656 38428 87662 38480
rect 60706 38372 80054 38400
rect 46661 38335 46719 38341
rect 46661 38301 46673 38335
rect 46707 38332 46719 38335
rect 72234 38332 72240 38344
rect 46707 38304 72240 38332
rect 46707 38301 46719 38304
rect 46661 38295 46719 38301
rect 72234 38292 72240 38304
rect 72292 38332 72298 38344
rect 73062 38332 73068 38344
rect 72292 38304 73068 38332
rect 72292 38292 72298 38304
rect 73062 38292 73068 38304
rect 73120 38292 73126 38344
rect 73341 38335 73399 38341
rect 73341 38301 73353 38335
rect 73387 38301 73399 38335
rect 73341 38295 73399 38301
rect 42576 38236 45554 38264
rect 48317 38267 48375 38273
rect 42576 38224 42582 38236
rect 48317 38233 48329 38267
rect 48363 38264 48375 38267
rect 48406 38264 48412 38276
rect 48363 38236 48412 38264
rect 48363 38233 48375 38236
rect 48317 38227 48375 38233
rect 48406 38224 48412 38236
rect 48464 38224 48470 38276
rect 7285 38199 7343 38205
rect 7285 38165 7297 38199
rect 7331 38196 7343 38199
rect 7561 38199 7619 38205
rect 7561 38196 7573 38199
rect 7331 38168 7573 38196
rect 7331 38165 7343 38168
rect 7285 38159 7343 38165
rect 7561 38165 7573 38168
rect 7607 38196 7619 38199
rect 10870 38196 10876 38208
rect 7607 38168 10876 38196
rect 7607 38165 7619 38168
rect 7561 38159 7619 38165
rect 10870 38156 10876 38168
rect 10928 38156 10934 38208
rect 24394 38156 24400 38208
rect 24452 38196 24458 38208
rect 26234 38196 26240 38208
rect 24452 38168 26240 38196
rect 24452 38156 24458 38168
rect 26234 38156 26240 38168
rect 26292 38156 26298 38208
rect 33781 38199 33839 38205
rect 33781 38165 33793 38199
rect 33827 38196 33839 38199
rect 34054 38196 34060 38208
rect 33827 38168 34060 38196
rect 33827 38165 33839 38168
rect 33781 38159 33839 38165
rect 34054 38156 34060 38168
rect 34112 38156 34118 38208
rect 73356 38196 73384 38295
rect 73522 38292 73528 38344
rect 73580 38332 73586 38344
rect 73617 38335 73675 38341
rect 73617 38332 73629 38335
rect 73580 38304 73629 38332
rect 73580 38292 73586 38304
rect 73617 38301 73629 38304
rect 73663 38301 73675 38335
rect 74718 38332 74724 38344
rect 74679 38304 74724 38332
rect 73617 38295 73675 38301
rect 74718 38292 74724 38304
rect 74776 38292 74782 38344
rect 74442 38224 74448 38276
rect 74500 38264 74506 38276
rect 91830 38264 91836 38276
rect 74500 38236 91836 38264
rect 74500 38224 74506 38236
rect 91830 38224 91836 38236
rect 91888 38224 91894 38276
rect 73614 38196 73620 38208
rect 73356 38168 73620 38196
rect 73614 38156 73620 38168
rect 73672 38196 73678 38208
rect 77570 38196 77576 38208
rect 73672 38168 77576 38196
rect 73672 38156 73678 38168
rect 77570 38156 77576 38168
rect 77628 38196 77634 38208
rect 81158 38196 81164 38208
rect 77628 38168 81164 38196
rect 77628 38156 77634 38168
rect 81158 38156 81164 38168
rect 81216 38156 81222 38208
rect 1104 38106 98808 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 65686 38106
rect 65738 38054 65750 38106
rect 65802 38054 65814 38106
rect 65866 38054 65878 38106
rect 65930 38054 96406 38106
rect 96458 38054 96470 38106
rect 96522 38054 96534 38106
rect 96586 38054 96598 38106
rect 96650 38054 98808 38106
rect 1104 38032 98808 38054
rect 11238 37992 11244 38004
rect 9140 37964 11244 37992
rect 9140 37865 9168 37964
rect 11238 37952 11244 37964
rect 11296 37992 11302 38004
rect 17678 37992 17684 38004
rect 11296 37964 17684 37992
rect 11296 37952 11302 37964
rect 17678 37952 17684 37964
rect 17736 37952 17742 38004
rect 17788 37964 26096 37992
rect 17494 37884 17500 37936
rect 17552 37924 17558 37936
rect 17788 37924 17816 37964
rect 17552 37896 17816 37924
rect 17552 37884 17558 37896
rect 17862 37884 17868 37936
rect 17920 37924 17926 37936
rect 25869 37927 25927 37933
rect 25869 37924 25881 37927
rect 17920 37896 25881 37924
rect 17920 37884 17926 37896
rect 25869 37893 25881 37896
rect 25915 37893 25927 37927
rect 26068 37924 26096 37964
rect 26234 37952 26240 38004
rect 26292 37992 26298 38004
rect 78398 37992 78404 38004
rect 26292 37964 48636 37992
rect 78359 37964 78404 37992
rect 26292 37952 26298 37964
rect 42886 37924 42892 37936
rect 26068 37896 42892 37924
rect 25869 37887 25927 37893
rect 42886 37884 42892 37896
rect 42944 37924 42950 37936
rect 43346 37924 43352 37936
rect 42944 37896 43352 37924
rect 42944 37884 42950 37896
rect 43346 37884 43352 37896
rect 43404 37884 43410 37936
rect 47026 37924 47032 37936
rect 45526 37896 46796 37924
rect 46987 37896 47032 37924
rect 9125 37859 9183 37865
rect 9125 37825 9137 37859
rect 9171 37825 9183 37859
rect 9125 37819 9183 37825
rect 6086 37748 6092 37800
rect 6144 37788 6150 37800
rect 6730 37788 6736 37800
rect 6144 37760 6736 37788
rect 6144 37748 6150 37760
rect 6730 37748 6736 37760
rect 6788 37788 6794 37800
rect 9140 37788 9168 37819
rect 10962 37816 10968 37868
rect 11020 37856 11026 37868
rect 45526 37856 45554 37896
rect 46658 37856 46664 37868
rect 11020 37828 45554 37856
rect 46124 37828 46520 37856
rect 46619 37828 46664 37856
rect 11020 37816 11026 37828
rect 9398 37788 9404 37800
rect 6788 37760 9168 37788
rect 9359 37760 9404 37788
rect 6788 37748 6794 37760
rect 9398 37748 9404 37760
rect 9456 37748 9462 37800
rect 12434 37748 12440 37800
rect 12492 37788 12498 37800
rect 17034 37788 17040 37800
rect 12492 37760 17040 37788
rect 12492 37748 12498 37760
rect 17034 37748 17040 37760
rect 17092 37788 17098 37800
rect 17862 37788 17868 37800
rect 17092 37760 17868 37788
rect 17092 37748 17098 37760
rect 17862 37748 17868 37760
rect 17920 37748 17926 37800
rect 19613 37791 19671 37797
rect 19613 37757 19625 37791
rect 19659 37788 19671 37791
rect 19886 37788 19892 37800
rect 19659 37760 19892 37788
rect 19659 37757 19671 37760
rect 19613 37751 19671 37757
rect 19886 37748 19892 37760
rect 19944 37748 19950 37800
rect 26053 37791 26111 37797
rect 26053 37757 26065 37791
rect 26099 37788 26111 37791
rect 26326 37788 26332 37800
rect 26099 37760 26332 37788
rect 26099 37757 26111 37760
rect 26053 37751 26111 37757
rect 26326 37748 26332 37760
rect 26384 37748 26390 37800
rect 46124 37797 46152 37828
rect 27157 37791 27215 37797
rect 26436 37760 27108 37788
rect 10781 37723 10839 37729
rect 10428 37692 10640 37720
rect 5442 37612 5448 37664
rect 5500 37652 5506 37664
rect 10428 37652 10456 37692
rect 5500 37624 10456 37652
rect 10612 37652 10640 37692
rect 10781 37689 10793 37723
rect 10827 37720 10839 37723
rect 26436 37720 26464 37760
rect 10827 37692 26464 37720
rect 27080 37720 27108 37760
rect 27157 37757 27169 37791
rect 27203 37788 27215 37791
rect 46109 37791 46167 37797
rect 46109 37788 46121 37791
rect 27203 37760 46121 37788
rect 27203 37757 27215 37760
rect 27157 37751 27215 37757
rect 46109 37757 46121 37760
rect 46155 37757 46167 37791
rect 46290 37788 46296 37800
rect 46251 37760 46296 37788
rect 46109 37751 46167 37757
rect 46290 37748 46296 37760
rect 46348 37748 46354 37800
rect 46492 37797 46520 37828
rect 46658 37816 46664 37828
rect 46716 37816 46722 37868
rect 46768 37856 46796 37896
rect 47026 37884 47032 37896
rect 47084 37884 47090 37936
rect 48406 37856 48412 37868
rect 46768 37828 48412 37856
rect 48406 37816 48412 37828
rect 48464 37816 48470 37868
rect 46476 37791 46534 37797
rect 46476 37757 46488 37791
rect 46522 37757 46534 37791
rect 46476 37751 46534 37757
rect 46566 37748 46572 37800
rect 46624 37788 46630 37800
rect 46842 37788 46848 37800
rect 46624 37760 46717 37788
rect 46803 37760 46848 37788
rect 46624 37748 46630 37760
rect 43806 37720 43812 37732
rect 27080 37692 43812 37720
rect 10827 37689 10839 37692
rect 10781 37683 10839 37689
rect 43806 37680 43812 37692
rect 43864 37680 43870 37732
rect 46676 37720 46704 37760
rect 46842 37748 46848 37760
rect 46900 37748 46906 37800
rect 48608 37788 48636 37964
rect 78398 37952 78404 37964
rect 78456 37952 78462 38004
rect 81158 37952 81164 38004
rect 81216 37992 81222 38004
rect 87325 37995 87383 38001
rect 81216 37964 86954 37992
rect 81216 37952 81222 37964
rect 78416 37856 78444 37952
rect 86926 37924 86954 37964
rect 87325 37961 87337 37995
rect 87371 37992 87383 37995
rect 89806 37992 89812 38004
rect 87371 37964 89812 37992
rect 87371 37961 87383 37964
rect 87325 37955 87383 37961
rect 89806 37952 89812 37964
rect 89864 37952 89870 38004
rect 92382 37924 92388 37936
rect 86926 37896 92388 37924
rect 92382 37884 92388 37896
rect 92440 37884 92446 37936
rect 78950 37856 78956 37868
rect 78416 37828 78812 37856
rect 78911 37828 78956 37856
rect 49510 37788 49516 37800
rect 48608 37760 49516 37788
rect 49510 37748 49516 37760
rect 49568 37788 49574 37800
rect 50617 37791 50675 37797
rect 50617 37788 50629 37791
rect 49568 37760 50629 37788
rect 49568 37748 49574 37760
rect 50617 37757 50629 37760
rect 50663 37757 50675 37791
rect 50890 37788 50896 37800
rect 50851 37760 50896 37788
rect 50617 37751 50675 37757
rect 50890 37748 50896 37760
rect 50948 37748 50954 37800
rect 73709 37791 73767 37797
rect 73709 37757 73721 37791
rect 73755 37757 73767 37791
rect 78582 37788 78588 37800
rect 78543 37760 78588 37788
rect 73709 37751 73767 37757
rect 57330 37720 57336 37732
rect 46676 37692 57336 37720
rect 57330 37680 57336 37692
rect 57388 37720 57394 37732
rect 57698 37720 57704 37732
rect 57388 37692 57704 37720
rect 57388 37680 57394 37692
rect 57698 37680 57704 37692
rect 57756 37680 57762 37732
rect 18506 37652 18512 37664
rect 10612 37624 18512 37652
rect 5500 37612 5506 37624
rect 18506 37612 18512 37624
rect 18564 37612 18570 37664
rect 25869 37655 25927 37661
rect 25869 37621 25881 37655
rect 25915 37652 25927 37655
rect 27157 37655 27215 37661
rect 27157 37652 27169 37655
rect 25915 37624 27169 37652
rect 25915 37621 25927 37624
rect 25869 37615 25927 37621
rect 27157 37621 27169 37624
rect 27203 37621 27215 37655
rect 27157 37615 27215 37621
rect 50154 37612 50160 37664
rect 50212 37652 50218 37664
rect 50433 37655 50491 37661
rect 50433 37652 50445 37655
rect 50212 37624 50445 37652
rect 50212 37612 50218 37624
rect 50433 37621 50445 37624
rect 50479 37621 50491 37655
rect 50798 37652 50804 37664
rect 50759 37624 50804 37652
rect 50433 37615 50491 37621
rect 50798 37612 50804 37624
rect 50856 37612 50862 37664
rect 73522 37652 73528 37664
rect 73483 37624 73528 37652
rect 73522 37612 73528 37624
rect 73580 37652 73586 37664
rect 73724 37652 73752 37751
rect 78582 37748 78588 37760
rect 78640 37748 78646 37800
rect 78784 37797 78812 37828
rect 78950 37816 78956 37828
rect 79008 37816 79014 37868
rect 81158 37856 81164 37868
rect 81119 37828 81164 37856
rect 81158 37816 81164 37828
rect 81216 37816 81222 37868
rect 81437 37859 81495 37865
rect 81437 37825 81449 37859
rect 81483 37856 81495 37859
rect 87325 37859 87383 37865
rect 87325 37856 87337 37859
rect 81483 37828 87337 37856
rect 81483 37825 81495 37828
rect 81437 37819 81495 37825
rect 87325 37825 87337 37828
rect 87371 37825 87383 37859
rect 87690 37856 87696 37868
rect 87651 37828 87696 37856
rect 87325 37819 87383 37825
rect 87690 37816 87696 37828
rect 87748 37816 87754 37868
rect 87782 37816 87788 37868
rect 87840 37856 87846 37868
rect 87877 37859 87935 37865
rect 87877 37856 87889 37859
rect 87840 37828 87889 37856
rect 87840 37816 87846 37828
rect 87877 37825 87889 37828
rect 87923 37856 87935 37859
rect 88429 37859 88487 37865
rect 88429 37856 88441 37859
rect 87923 37828 88441 37856
rect 87923 37825 87935 37828
rect 87877 37819 87935 37825
rect 88429 37825 88441 37828
rect 88475 37825 88487 37859
rect 88429 37819 88487 37825
rect 78768 37791 78826 37797
rect 78768 37757 78780 37791
rect 78814 37757 78826 37791
rect 78768 37751 78826 37757
rect 78858 37748 78864 37800
rect 78916 37788 78922 37800
rect 79134 37797 79140 37800
rect 79110 37791 79140 37797
rect 78916 37760 78961 37788
rect 78916 37748 78922 37760
rect 79110 37757 79122 37791
rect 79192 37788 79198 37800
rect 93854 37788 93860 37800
rect 79192 37760 93860 37788
rect 79110 37751 79140 37757
rect 79134 37748 79140 37751
rect 79192 37748 79198 37760
rect 93854 37748 93860 37760
rect 93912 37748 93918 37800
rect 87506 37720 87512 37732
rect 87467 37692 87512 37720
rect 87506 37680 87512 37692
rect 87564 37720 87570 37732
rect 87969 37723 88027 37729
rect 87969 37720 87981 37723
rect 87564 37692 87981 37720
rect 87564 37680 87570 37692
rect 87969 37689 87981 37692
rect 88015 37689 88027 37723
rect 89622 37720 89628 37732
rect 87969 37683 88027 37689
rect 88076 37692 89628 37720
rect 79226 37652 79232 37664
rect 73580 37624 73752 37652
rect 79187 37624 79232 37652
rect 73580 37612 73586 37624
rect 79226 37612 79232 37624
rect 79284 37612 79290 37664
rect 82538 37652 82544 37664
rect 82499 37624 82544 37652
rect 82538 37612 82544 37624
rect 82596 37652 82602 37664
rect 88076 37652 88104 37692
rect 89622 37680 89628 37692
rect 89680 37680 89686 37732
rect 82596 37624 88104 37652
rect 88337 37655 88395 37661
rect 82596 37612 82602 37624
rect 88337 37621 88349 37655
rect 88383 37652 88395 37655
rect 92658 37652 92664 37664
rect 88383 37624 92664 37652
rect 88383 37621 88395 37624
rect 88337 37615 88395 37621
rect 92658 37612 92664 37624
rect 92716 37612 92722 37664
rect 1104 37562 98808 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 50326 37562
rect 50378 37510 50390 37562
rect 50442 37510 50454 37562
rect 50506 37510 50518 37562
rect 50570 37510 81046 37562
rect 81098 37510 81110 37562
rect 81162 37510 81174 37562
rect 81226 37510 81238 37562
rect 81290 37510 98808 37562
rect 1104 37488 98808 37510
rect 17589 37451 17647 37457
rect 17589 37417 17601 37451
rect 17635 37448 17647 37451
rect 17954 37448 17960 37460
rect 17635 37420 17960 37448
rect 17635 37417 17647 37420
rect 17589 37411 17647 37417
rect 17954 37408 17960 37420
rect 18012 37408 18018 37460
rect 20714 37448 20720 37460
rect 18340 37420 20720 37448
rect 12897 37383 12955 37389
rect 12897 37349 12909 37383
rect 12943 37380 12955 37383
rect 12986 37380 12992 37392
rect 12943 37352 12992 37380
rect 12943 37349 12955 37352
rect 12897 37343 12955 37349
rect 12986 37340 12992 37352
rect 13044 37340 13050 37392
rect 11238 37312 11244 37324
rect 11199 37284 11244 37312
rect 11238 37272 11244 37284
rect 11296 37272 11302 37324
rect 11514 37312 11520 37324
rect 11475 37284 11520 37312
rect 11514 37272 11520 37284
rect 11572 37272 11578 37324
rect 17770 37312 17776 37324
rect 17731 37284 17776 37312
rect 17770 37272 17776 37284
rect 17828 37272 17834 37324
rect 17972 37312 18000 37408
rect 18340 37321 18368 37420
rect 20714 37408 20720 37420
rect 20772 37448 20778 37460
rect 20990 37448 20996 37460
rect 20772 37420 20996 37448
rect 20772 37408 20778 37420
rect 20990 37408 20996 37420
rect 21048 37408 21054 37460
rect 52362 37408 52368 37460
rect 52420 37448 52426 37460
rect 52420 37420 84194 37448
rect 52420 37408 52426 37420
rect 18506 37340 18512 37392
rect 18564 37380 18570 37392
rect 36170 37380 36176 37392
rect 18564 37352 36176 37380
rect 18564 37340 18570 37352
rect 18141 37315 18199 37321
rect 18141 37312 18153 37315
rect 17972 37284 18153 37312
rect 18141 37281 18153 37284
rect 18187 37312 18199 37315
rect 18325 37315 18383 37321
rect 18187 37284 18276 37312
rect 18187 37281 18199 37284
rect 18141 37275 18199 37281
rect 18248 37244 18276 37284
rect 18325 37281 18337 37315
rect 18371 37281 18383 37315
rect 18598 37312 18604 37324
rect 18559 37284 18604 37312
rect 18325 37275 18383 37281
rect 18598 37272 18604 37284
rect 18656 37272 18662 37324
rect 18708 37321 18736 37352
rect 36170 37340 36176 37352
rect 36228 37380 36234 37392
rect 36228 37352 60734 37380
rect 36228 37340 36234 37352
rect 18693 37315 18751 37321
rect 18693 37281 18705 37315
rect 18739 37281 18751 37315
rect 18693 37275 18751 37281
rect 19061 37315 19119 37321
rect 19061 37281 19073 37315
rect 19107 37312 19119 37315
rect 19978 37312 19984 37324
rect 19107 37284 19984 37312
rect 19107 37281 19119 37284
rect 19061 37275 19119 37281
rect 19978 37272 19984 37284
rect 20036 37272 20042 37324
rect 60706 37312 60734 37352
rect 73246 37340 73252 37392
rect 73304 37380 73310 37392
rect 73525 37383 73583 37389
rect 73525 37380 73537 37383
rect 73304 37352 73537 37380
rect 73304 37340 73310 37352
rect 73525 37349 73537 37352
rect 73571 37349 73583 37383
rect 78677 37383 78735 37389
rect 78677 37380 78689 37383
rect 73525 37343 73583 37349
rect 73632 37352 78689 37380
rect 73632 37312 73660 37352
rect 78677 37349 78689 37352
rect 78723 37349 78735 37383
rect 78677 37343 78735 37349
rect 60706 37284 73660 37312
rect 73985 37315 74043 37321
rect 73985 37281 73997 37315
rect 74031 37312 74043 37315
rect 74074 37312 74080 37324
rect 74031 37284 74080 37312
rect 74031 37281 74043 37284
rect 73985 37275 74043 37281
rect 74074 37272 74080 37284
rect 74132 37272 74138 37324
rect 74169 37315 74227 37321
rect 74169 37281 74181 37315
rect 74215 37312 74227 37315
rect 74534 37312 74540 37324
rect 74215 37284 74304 37312
rect 74495 37284 74540 37312
rect 74215 37281 74227 37284
rect 74169 37275 74227 37281
rect 18506 37244 18512 37256
rect 18248 37216 18512 37244
rect 18506 37204 18512 37216
rect 18564 37204 18570 37256
rect 74276 37176 74304 37284
rect 74534 37272 74540 37284
rect 74592 37272 74598 37324
rect 76374 37312 76380 37324
rect 74644 37284 76380 37312
rect 74442 37244 74448 37256
rect 74403 37216 74448 37244
rect 74442 37204 74448 37216
rect 74500 37204 74506 37256
rect 74644 37176 74672 37284
rect 76374 37272 76380 37284
rect 76432 37272 76438 37324
rect 77941 37315 77999 37321
rect 77941 37281 77953 37315
rect 77987 37312 77999 37315
rect 79686 37312 79692 37324
rect 77987 37284 79692 37312
rect 77987 37281 77999 37284
rect 77941 37275 77999 37281
rect 79686 37272 79692 37284
rect 79744 37272 79750 37324
rect 84166 37312 84194 37420
rect 87506 37408 87512 37460
rect 87564 37448 87570 37460
rect 87966 37448 87972 37460
rect 87564 37420 87972 37448
rect 87564 37408 87570 37420
rect 87966 37408 87972 37420
rect 88024 37408 88030 37460
rect 93857 37315 93915 37321
rect 93857 37312 93869 37315
rect 84166 37284 93869 37312
rect 93857 37281 93869 37284
rect 93903 37281 93915 37315
rect 94222 37312 94228 37324
rect 94183 37284 94228 37312
rect 93857 37275 93915 37281
rect 94222 37272 94228 37284
rect 94280 37272 94286 37324
rect 78030 37204 78036 37256
rect 78088 37244 78094 37256
rect 94317 37247 94375 37253
rect 94317 37244 94329 37247
rect 78088 37216 94329 37244
rect 78088 37204 78094 37216
rect 94317 37213 94329 37216
rect 94363 37213 94375 37247
rect 94317 37207 94375 37213
rect 74276 37148 74672 37176
rect 93026 37136 93032 37188
rect 93084 37176 93090 37188
rect 93673 37179 93731 37185
rect 93673 37176 93685 37179
rect 93084 37148 93685 37176
rect 93084 37136 93090 37148
rect 93673 37145 93685 37148
rect 93719 37145 93731 37179
rect 93673 37139 93731 37145
rect 83642 37068 83648 37120
rect 83700 37108 83706 37120
rect 84749 37111 84807 37117
rect 84749 37108 84761 37111
rect 83700 37080 84761 37108
rect 83700 37068 83706 37080
rect 84749 37077 84761 37080
rect 84795 37108 84807 37111
rect 84841 37111 84899 37117
rect 84841 37108 84853 37111
rect 84795 37080 84853 37108
rect 84795 37077 84807 37080
rect 84749 37071 84807 37077
rect 84841 37077 84853 37080
rect 84887 37077 84899 37111
rect 84841 37071 84899 37077
rect 1104 37018 98808 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 65686 37018
rect 65738 36966 65750 37018
rect 65802 36966 65814 37018
rect 65866 36966 65878 37018
rect 65930 36966 96406 37018
rect 96458 36966 96470 37018
rect 96522 36966 96534 37018
rect 96586 36966 96598 37018
rect 96650 36966 98808 37018
rect 1104 36944 98808 36966
rect 3326 36904 3332 36916
rect 3287 36876 3332 36904
rect 3326 36864 3332 36876
rect 3384 36864 3390 36916
rect 49602 36864 49608 36916
rect 49660 36904 49666 36916
rect 76190 36904 76196 36916
rect 49660 36876 70394 36904
rect 76151 36876 76196 36904
rect 49660 36864 49666 36876
rect 33686 36796 33692 36848
rect 33744 36836 33750 36848
rect 63310 36836 63316 36848
rect 33744 36808 63316 36836
rect 33744 36796 33750 36808
rect 63310 36796 63316 36808
rect 63368 36796 63374 36848
rect 70366 36836 70394 36876
rect 76190 36864 76196 36876
rect 76248 36864 76254 36916
rect 70366 36808 90864 36836
rect 3145 36771 3203 36777
rect 3145 36737 3157 36771
rect 3191 36768 3203 36771
rect 5994 36768 6000 36780
rect 3191 36740 6000 36768
rect 3191 36737 3203 36740
rect 3145 36731 3203 36737
rect 3528 36709 3556 36740
rect 5994 36728 6000 36740
rect 6052 36768 6058 36780
rect 9950 36768 9956 36780
rect 6052 36740 9956 36768
rect 6052 36728 6058 36740
rect 9950 36728 9956 36740
rect 10008 36768 10014 36780
rect 52362 36768 52368 36780
rect 10008 36740 52368 36768
rect 10008 36728 10014 36740
rect 52362 36728 52368 36740
rect 52420 36728 52426 36780
rect 57330 36728 57336 36780
rect 57388 36768 57394 36780
rect 89254 36768 89260 36780
rect 57388 36740 89260 36768
rect 57388 36728 57394 36740
rect 89254 36728 89260 36740
rect 89312 36768 89318 36780
rect 89312 36740 89576 36768
rect 89312 36728 89318 36740
rect 3513 36703 3571 36709
rect 3513 36669 3525 36703
rect 3559 36669 3571 36703
rect 3513 36663 3571 36669
rect 3697 36703 3755 36709
rect 3697 36669 3709 36703
rect 3743 36700 3755 36703
rect 8202 36700 8208 36712
rect 3743 36672 8208 36700
rect 3743 36669 3755 36672
rect 3697 36663 3755 36669
rect 8202 36660 8208 36672
rect 8260 36660 8266 36712
rect 16022 36660 16028 36712
rect 16080 36700 16086 36712
rect 49602 36700 49608 36712
rect 16080 36672 49608 36700
rect 16080 36660 16086 36672
rect 49602 36660 49608 36672
rect 49660 36660 49666 36712
rect 74994 36700 75000 36712
rect 74955 36672 75000 36700
rect 74994 36660 75000 36672
rect 75052 36660 75058 36712
rect 75178 36700 75184 36712
rect 75139 36672 75184 36700
rect 75178 36660 75184 36672
rect 75236 36660 75242 36712
rect 75362 36700 75368 36712
rect 75323 36672 75368 36700
rect 75362 36660 75368 36672
rect 75420 36660 75426 36712
rect 75730 36700 75736 36712
rect 75691 36672 75736 36700
rect 75730 36660 75736 36672
rect 75788 36660 75794 36712
rect 75822 36660 75828 36712
rect 75880 36700 75886 36712
rect 75917 36703 75975 36709
rect 75917 36700 75929 36703
rect 75880 36672 75929 36700
rect 75880 36660 75886 36672
rect 75917 36669 75929 36672
rect 75963 36669 75975 36703
rect 87601 36703 87659 36709
rect 87601 36700 87613 36703
rect 75917 36663 75975 36669
rect 84166 36672 87613 36700
rect 3789 36635 3847 36641
rect 3789 36601 3801 36635
rect 3835 36601 3847 36635
rect 3789 36595 3847 36601
rect 3804 36564 3832 36595
rect 6454 36592 6460 36644
rect 6512 36632 6518 36644
rect 19426 36632 19432 36644
rect 6512 36604 19432 36632
rect 6512 36592 6518 36604
rect 19426 36592 19432 36604
rect 19484 36632 19490 36644
rect 20622 36632 20628 36644
rect 19484 36604 20628 36632
rect 19484 36592 19490 36604
rect 20622 36592 20628 36604
rect 20680 36592 20686 36644
rect 48406 36592 48412 36644
rect 48464 36632 48470 36644
rect 84166 36632 84194 36672
rect 87601 36669 87613 36672
rect 87647 36669 87659 36703
rect 88426 36700 88432 36712
rect 88387 36672 88432 36700
rect 87601 36663 87659 36669
rect 88426 36660 88432 36672
rect 88484 36660 88490 36712
rect 48464 36604 60734 36632
rect 48464 36592 48470 36604
rect 3973 36567 4031 36573
rect 3973 36564 3985 36567
rect 3804 36536 3985 36564
rect 3973 36533 3985 36536
rect 4019 36564 4031 36567
rect 8570 36564 8576 36576
rect 4019 36536 8576 36564
rect 4019 36533 4031 36536
rect 3973 36527 4031 36533
rect 8570 36524 8576 36536
rect 8628 36564 8634 36576
rect 59262 36564 59268 36576
rect 8628 36536 59268 36564
rect 8628 36524 8634 36536
rect 59262 36524 59268 36536
rect 59320 36524 59326 36576
rect 60706 36564 60734 36604
rect 75656 36604 84194 36632
rect 89548 36632 89576 36740
rect 90836 36709 90864 36808
rect 90821 36703 90879 36709
rect 90821 36669 90833 36703
rect 90867 36669 90879 36703
rect 90821 36663 90879 36669
rect 91189 36635 91247 36641
rect 91189 36632 91201 36635
rect 89548 36604 91201 36632
rect 75656 36564 75684 36604
rect 91189 36601 91201 36604
rect 91235 36601 91247 36635
rect 91189 36595 91247 36601
rect 88426 36564 88432 36576
rect 60706 36536 75684 36564
rect 88387 36536 88432 36564
rect 88426 36524 88432 36536
rect 88484 36524 88490 36576
rect 1104 36474 98808 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 50326 36474
rect 50378 36422 50390 36474
rect 50442 36422 50454 36474
rect 50506 36422 50518 36474
rect 50570 36422 81046 36474
rect 81098 36422 81110 36474
rect 81162 36422 81174 36474
rect 81226 36422 81238 36474
rect 81290 36422 98808 36474
rect 1104 36400 98808 36422
rect 20622 36320 20628 36372
rect 20680 36360 20686 36372
rect 51261 36363 51319 36369
rect 51261 36360 51273 36363
rect 20680 36332 51273 36360
rect 20680 36320 20686 36332
rect 51261 36329 51273 36332
rect 51307 36360 51319 36363
rect 51350 36360 51356 36372
rect 51307 36332 51356 36360
rect 51307 36329 51319 36332
rect 51261 36323 51319 36329
rect 51350 36320 51356 36332
rect 51408 36320 51414 36372
rect 51442 36320 51448 36372
rect 51500 36360 51506 36372
rect 66806 36360 66812 36372
rect 51500 36332 66812 36360
rect 51500 36320 51506 36332
rect 66806 36320 66812 36332
rect 66864 36360 66870 36372
rect 66864 36332 74304 36360
rect 66864 36320 66870 36332
rect 40862 36252 40868 36304
rect 40920 36292 40926 36304
rect 41322 36292 41328 36304
rect 40920 36264 41328 36292
rect 40920 36252 40926 36264
rect 41322 36252 41328 36264
rect 41380 36292 41386 36304
rect 41380 36264 63264 36292
rect 41380 36252 41386 36264
rect 35802 36224 35808 36236
rect 35763 36196 35808 36224
rect 35802 36184 35808 36196
rect 35860 36184 35866 36236
rect 42058 36184 42064 36236
rect 42116 36224 42122 36236
rect 51442 36224 51448 36236
rect 42116 36196 51448 36224
rect 42116 36184 42122 36196
rect 51442 36184 51448 36196
rect 51500 36184 51506 36236
rect 51626 36184 51632 36236
rect 51684 36224 51690 36236
rect 51810 36224 51816 36236
rect 51684 36196 51728 36224
rect 51771 36196 51816 36224
rect 51684 36184 51690 36196
rect 51810 36184 51816 36196
rect 51868 36184 51874 36236
rect 51997 36227 52055 36233
rect 51997 36224 52009 36227
rect 51920 36196 52009 36224
rect 51920 36168 51948 36196
rect 51997 36193 52009 36196
rect 52043 36193 52055 36227
rect 52178 36224 52184 36236
rect 52139 36196 52184 36224
rect 51997 36187 52055 36193
rect 52178 36184 52184 36196
rect 52236 36184 52242 36236
rect 63034 36224 63040 36236
rect 62995 36196 63040 36224
rect 63034 36184 63040 36196
rect 63092 36184 63098 36236
rect 63236 36233 63264 36264
rect 63220 36227 63278 36233
rect 63220 36193 63232 36227
rect 63266 36193 63278 36227
rect 63586 36224 63592 36236
rect 63499 36196 63592 36224
rect 63220 36187 63278 36193
rect 63586 36184 63592 36196
rect 63644 36224 63650 36236
rect 64690 36224 64696 36236
rect 63644 36196 64696 36224
rect 63644 36184 63650 36196
rect 64690 36184 64696 36196
rect 64748 36184 64754 36236
rect 74276 36224 74304 36332
rect 75730 36320 75736 36372
rect 75788 36360 75794 36372
rect 76006 36360 76012 36372
rect 75788 36332 76012 36360
rect 75788 36320 75794 36332
rect 76006 36320 76012 36332
rect 76064 36360 76070 36372
rect 76926 36360 76932 36372
rect 76064 36332 76932 36360
rect 76064 36320 76070 36332
rect 76926 36320 76932 36332
rect 76984 36320 76990 36372
rect 75362 36252 75368 36304
rect 75420 36292 75426 36304
rect 75914 36292 75920 36304
rect 75420 36264 75920 36292
rect 75420 36252 75426 36264
rect 75914 36252 75920 36264
rect 75972 36292 75978 36304
rect 76742 36292 76748 36304
rect 75972 36264 76748 36292
rect 75972 36252 75978 36264
rect 76742 36252 76748 36264
rect 76800 36252 76806 36304
rect 78953 36295 79011 36301
rect 78953 36292 78965 36295
rect 78140 36264 78965 36292
rect 77665 36227 77723 36233
rect 77665 36224 77677 36227
rect 74276 36196 77677 36224
rect 77665 36193 77677 36196
rect 77711 36193 77723 36227
rect 78033 36227 78091 36233
rect 78033 36224 78045 36227
rect 77665 36187 77723 36193
rect 77772 36196 78045 36224
rect 20714 36116 20720 36168
rect 20772 36156 20778 36168
rect 36541 36159 36599 36165
rect 36541 36156 36553 36159
rect 20772 36128 36553 36156
rect 20772 36116 20778 36128
rect 36541 36125 36553 36128
rect 36587 36156 36599 36159
rect 39758 36156 39764 36168
rect 36587 36128 39764 36156
rect 36587 36125 36599 36128
rect 36541 36119 36599 36125
rect 39758 36116 39764 36128
rect 39816 36116 39822 36168
rect 51718 36156 51724 36168
rect 51679 36128 51724 36156
rect 51718 36116 51724 36128
rect 51776 36116 51782 36168
rect 51902 36116 51908 36168
rect 51960 36116 51966 36168
rect 63310 36156 63316 36168
rect 63271 36128 63316 36156
rect 63310 36116 63316 36128
rect 63368 36116 63374 36168
rect 63402 36116 63408 36168
rect 63460 36156 63466 36168
rect 63460 36128 63505 36156
rect 63460 36116 63466 36128
rect 74258 36116 74264 36168
rect 74316 36156 74322 36168
rect 77772 36156 77800 36196
rect 78033 36193 78045 36196
rect 78079 36193 78091 36227
rect 78033 36187 78091 36193
rect 77938 36156 77944 36168
rect 74316 36128 77800 36156
rect 77899 36128 77944 36156
rect 74316 36116 74322 36128
rect 77938 36116 77944 36128
rect 77996 36116 78002 36168
rect 23566 36048 23572 36100
rect 23624 36088 23630 36100
rect 78140 36088 78168 36264
rect 78953 36261 78965 36264
rect 78999 36261 79011 36295
rect 78953 36255 79011 36261
rect 78306 36224 78312 36236
rect 78267 36196 78312 36224
rect 78306 36184 78312 36196
rect 78364 36184 78370 36236
rect 78401 36227 78459 36233
rect 78401 36193 78413 36227
rect 78447 36193 78459 36227
rect 78401 36187 78459 36193
rect 23624 36060 45554 36088
rect 23624 36048 23630 36060
rect 45526 36020 45554 36060
rect 60706 36060 78168 36088
rect 60706 36020 60734 36060
rect 63678 36020 63684 36032
rect 45526 35992 60734 36020
rect 63639 35992 63684 36020
rect 63678 35980 63684 35992
rect 63736 35980 63742 36032
rect 70302 35980 70308 36032
rect 70360 36020 70366 36032
rect 78416 36020 78444 36187
rect 70360 35992 78444 36020
rect 70360 35980 70366 35992
rect 1104 35930 98808 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 65686 35930
rect 65738 35878 65750 35930
rect 65802 35878 65814 35930
rect 65866 35878 65878 35930
rect 65930 35878 96406 35930
rect 96458 35878 96470 35930
rect 96522 35878 96534 35930
rect 96586 35878 96598 35930
rect 96650 35878 98808 35930
rect 1104 35856 98808 35878
rect 57330 35776 57336 35828
rect 57388 35816 57394 35828
rect 57606 35816 57612 35828
rect 57388 35788 57612 35816
rect 57388 35776 57394 35788
rect 57606 35776 57612 35788
rect 57664 35776 57670 35828
rect 73430 35776 73436 35828
rect 73488 35816 73494 35828
rect 73982 35816 73988 35828
rect 73488 35788 73988 35816
rect 73488 35776 73494 35788
rect 73982 35776 73988 35788
rect 74040 35776 74046 35828
rect 11790 35572 11796 35624
rect 11848 35612 11854 35624
rect 73798 35612 73804 35624
rect 11848 35584 73804 35612
rect 11848 35572 11854 35584
rect 73798 35572 73804 35584
rect 73856 35572 73862 35624
rect 74997 35615 75055 35621
rect 74997 35612 75009 35615
rect 74828 35584 75009 35612
rect 23934 35504 23940 35556
rect 23992 35544 23998 35556
rect 36262 35544 36268 35556
rect 23992 35516 36268 35544
rect 23992 35504 23998 35516
rect 36262 35504 36268 35516
rect 36320 35504 36326 35556
rect 9030 35436 9036 35488
rect 9088 35476 9094 35488
rect 31478 35476 31484 35488
rect 9088 35448 31484 35476
rect 9088 35436 9094 35448
rect 31478 35436 31484 35448
rect 31536 35436 31542 35488
rect 73890 35436 73896 35488
rect 73948 35476 73954 35488
rect 74828 35485 74856 35584
rect 74997 35581 75009 35584
rect 75043 35581 75055 35615
rect 74997 35575 75055 35581
rect 74813 35479 74871 35485
rect 74813 35476 74825 35479
rect 73948 35448 74825 35476
rect 73948 35436 73954 35448
rect 74813 35445 74825 35448
rect 74859 35445 74871 35479
rect 74813 35439 74871 35445
rect 1104 35386 98808 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 50326 35386
rect 50378 35334 50390 35386
rect 50442 35334 50454 35386
rect 50506 35334 50518 35386
rect 50570 35334 81046 35386
rect 81098 35334 81110 35386
rect 81162 35334 81174 35386
rect 81226 35334 81238 35386
rect 81290 35334 98808 35386
rect 1104 35312 98808 35334
rect 10042 35232 10048 35284
rect 10100 35272 10106 35284
rect 40034 35272 40040 35284
rect 10100 35244 40040 35272
rect 10100 35232 10106 35244
rect 40034 35232 40040 35244
rect 40092 35232 40098 35284
rect 42794 35164 42800 35216
rect 42852 35204 42858 35216
rect 51718 35204 51724 35216
rect 42852 35176 51724 35204
rect 42852 35164 42858 35176
rect 51718 35164 51724 35176
rect 51776 35164 51782 35216
rect 27709 35139 27767 35145
rect 27709 35105 27721 35139
rect 27755 35136 27767 35139
rect 39850 35136 39856 35148
rect 27755 35108 39856 35136
rect 27755 35105 27767 35108
rect 27709 35099 27767 35105
rect 39850 35096 39856 35108
rect 39908 35096 39914 35148
rect 63402 35096 63408 35148
rect 63460 35136 63466 35148
rect 72421 35139 72479 35145
rect 72421 35136 72433 35139
rect 63460 35108 72433 35136
rect 63460 35096 63466 35108
rect 72421 35105 72433 35108
rect 72467 35105 72479 35139
rect 72421 35099 72479 35105
rect 27433 35071 27491 35077
rect 27433 35037 27445 35071
rect 27479 35068 27491 35071
rect 31018 35068 31024 35080
rect 27479 35040 31024 35068
rect 27479 35037 27491 35040
rect 27433 35031 27491 35037
rect 31018 35028 31024 35040
rect 31076 35028 31082 35080
rect 31386 35028 31392 35080
rect 31444 35068 31450 35080
rect 72237 35071 72295 35077
rect 72237 35068 72249 35071
rect 31444 35040 72249 35068
rect 31444 35028 31450 35040
rect 72237 35037 72249 35040
rect 72283 35068 72295 35071
rect 72789 35071 72847 35077
rect 72789 35068 72801 35071
rect 72283 35040 72801 35068
rect 72283 35037 72295 35040
rect 72237 35031 72295 35037
rect 72789 35037 72801 35040
rect 72835 35037 72847 35071
rect 72789 35031 72847 35037
rect 66254 34960 66260 35012
rect 66312 35000 66318 35012
rect 66898 35000 66904 35012
rect 66312 34972 66904 35000
rect 66312 34960 66318 34972
rect 66898 34960 66904 34972
rect 66956 34960 66962 35012
rect 72697 35003 72755 35009
rect 72697 34969 72709 35003
rect 72743 35000 72755 35003
rect 73798 35000 73804 35012
rect 72743 34972 73804 35000
rect 72743 34969 72755 34972
rect 72697 34963 72755 34969
rect 73798 34960 73804 34972
rect 73856 34960 73862 35012
rect 28994 34932 29000 34944
rect 28955 34904 29000 34932
rect 28994 34892 29000 34904
rect 29052 34892 29058 34944
rect 65426 34892 65432 34944
rect 65484 34932 65490 34944
rect 66438 34932 66444 34944
rect 65484 34904 66444 34932
rect 65484 34892 65490 34904
rect 66438 34892 66444 34904
rect 66496 34892 66502 34944
rect 72326 34892 72332 34944
rect 72384 34932 72390 34944
rect 72559 34935 72617 34941
rect 72559 34932 72571 34935
rect 72384 34904 72571 34932
rect 72384 34892 72390 34904
rect 72559 34901 72571 34904
rect 72605 34901 72617 34935
rect 72559 34895 72617 34901
rect 73065 34935 73123 34941
rect 73065 34901 73077 34935
rect 73111 34932 73123 34935
rect 84378 34932 84384 34944
rect 73111 34904 84384 34932
rect 73111 34901 73123 34904
rect 73065 34895 73123 34901
rect 84378 34892 84384 34904
rect 84436 34892 84442 34944
rect 1104 34842 98808 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 65686 34842
rect 65738 34790 65750 34842
rect 65802 34790 65814 34842
rect 65866 34790 65878 34842
rect 65930 34790 96406 34842
rect 96458 34790 96470 34842
rect 96522 34790 96534 34842
rect 96586 34790 96598 34842
rect 96650 34790 98808 34842
rect 1104 34768 98808 34790
rect 28994 34688 29000 34740
rect 29052 34728 29058 34740
rect 53558 34728 53564 34740
rect 29052 34700 53564 34728
rect 29052 34688 29058 34700
rect 53558 34688 53564 34700
rect 53616 34728 53622 34740
rect 54662 34728 54668 34740
rect 53616 34700 54668 34728
rect 53616 34688 53622 34700
rect 54662 34688 54668 34700
rect 54720 34688 54726 34740
rect 57330 34688 57336 34740
rect 57388 34728 57394 34740
rect 65889 34731 65947 34737
rect 65889 34728 65901 34731
rect 57388 34700 65901 34728
rect 57388 34688 57394 34700
rect 65889 34697 65901 34700
rect 65935 34697 65947 34731
rect 65889 34691 65947 34697
rect 51810 34620 51816 34672
rect 51868 34660 51874 34672
rect 65426 34660 65432 34672
rect 51868 34632 65432 34660
rect 51868 34620 51874 34632
rect 65426 34620 65432 34632
rect 65484 34620 65490 34672
rect 65904 34660 65932 34691
rect 66438 34688 66444 34740
rect 66496 34728 66502 34740
rect 70302 34728 70308 34740
rect 66496 34700 70308 34728
rect 66496 34688 66502 34700
rect 70302 34688 70308 34700
rect 70360 34688 70366 34740
rect 66622 34660 66628 34672
rect 65904 34632 66628 34660
rect 66622 34620 66628 34632
rect 66680 34620 66686 34672
rect 66898 34620 66904 34672
rect 66956 34660 66962 34672
rect 66956 34632 67001 34660
rect 66956 34620 66962 34632
rect 43530 34552 43536 34604
rect 43588 34592 43594 34604
rect 48038 34592 48044 34604
rect 43588 34564 48044 34592
rect 43588 34552 43594 34564
rect 48038 34552 48044 34564
rect 48096 34552 48102 34604
rect 51718 34552 51724 34604
rect 51776 34592 51782 34604
rect 66533 34595 66591 34601
rect 66533 34592 66545 34595
rect 51776 34564 66545 34592
rect 51776 34552 51782 34564
rect 66533 34561 66545 34564
rect 66579 34592 66591 34595
rect 74258 34592 74264 34604
rect 66579 34564 74264 34592
rect 66579 34561 66591 34564
rect 66533 34555 66591 34561
rect 74258 34552 74264 34564
rect 74316 34552 74322 34604
rect 19886 34484 19892 34536
rect 19944 34524 19950 34536
rect 25682 34524 25688 34536
rect 19944 34496 25688 34524
rect 19944 34484 19950 34496
rect 25682 34484 25688 34496
rect 25740 34484 25746 34536
rect 33318 34484 33324 34536
rect 33376 34524 33382 34536
rect 66073 34527 66131 34533
rect 66073 34524 66085 34527
rect 33376 34496 66085 34524
rect 33376 34484 33382 34496
rect 66073 34493 66085 34496
rect 66119 34493 66131 34527
rect 66254 34524 66260 34536
rect 66215 34496 66260 34524
rect 66073 34487 66131 34493
rect 66254 34484 66260 34496
rect 66312 34484 66318 34536
rect 66438 34524 66444 34536
rect 66399 34496 66444 34524
rect 66438 34484 66444 34496
rect 66496 34484 66502 34536
rect 66622 34484 66628 34536
rect 66680 34524 66686 34536
rect 66812 34527 66870 34533
rect 66680 34496 66725 34524
rect 66680 34484 66686 34496
rect 66812 34493 66824 34527
rect 66858 34524 66870 34527
rect 66898 34524 66904 34536
rect 66858 34496 66904 34524
rect 66858 34493 66870 34496
rect 66812 34487 66870 34493
rect 66898 34484 66904 34496
rect 66956 34484 66962 34536
rect 67818 34524 67824 34536
rect 67779 34496 67824 34524
rect 67818 34484 67824 34496
rect 67876 34484 67882 34536
rect 68649 34527 68707 34533
rect 68649 34493 68661 34527
rect 68695 34524 68707 34527
rect 73430 34524 73436 34536
rect 68695 34496 73436 34524
rect 68695 34493 68707 34496
rect 68649 34487 68707 34493
rect 73430 34484 73436 34496
rect 73488 34484 73494 34536
rect 26510 34416 26516 34468
rect 26568 34456 26574 34468
rect 30374 34456 30380 34468
rect 26568 34428 30380 34456
rect 26568 34416 26574 34428
rect 30374 34416 30380 34428
rect 30432 34416 30438 34468
rect 41598 34416 41604 34468
rect 41656 34456 41662 34468
rect 65426 34456 65432 34468
rect 41656 34428 65432 34456
rect 41656 34416 41662 34428
rect 65426 34416 65432 34428
rect 65484 34416 65490 34468
rect 35250 34348 35256 34400
rect 35308 34388 35314 34400
rect 65610 34388 65616 34400
rect 35308 34360 65616 34388
rect 35308 34348 35314 34360
rect 65610 34348 65616 34360
rect 65668 34348 65674 34400
rect 1104 34298 98808 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 50326 34298
rect 50378 34246 50390 34298
rect 50442 34246 50454 34298
rect 50506 34246 50518 34298
rect 50570 34246 81046 34298
rect 81098 34246 81110 34298
rect 81162 34246 81174 34298
rect 81226 34246 81238 34298
rect 81290 34246 98808 34298
rect 1104 34224 98808 34246
rect 3510 34144 3516 34196
rect 3568 34184 3574 34196
rect 44174 34184 44180 34196
rect 3568 34156 44180 34184
rect 3568 34144 3574 34156
rect 44174 34144 44180 34156
rect 44232 34144 44238 34196
rect 56594 34184 56600 34196
rect 56555 34156 56600 34184
rect 56594 34144 56600 34156
rect 56652 34144 56658 34196
rect 65426 34144 65432 34196
rect 65484 34184 65490 34196
rect 73246 34184 73252 34196
rect 65484 34156 73252 34184
rect 65484 34144 65490 34156
rect 73246 34144 73252 34156
rect 73304 34144 73310 34196
rect 21637 34119 21695 34125
rect 21637 34085 21649 34119
rect 21683 34116 21695 34119
rect 21726 34116 21732 34128
rect 21683 34088 21732 34116
rect 21683 34085 21695 34088
rect 21637 34079 21695 34085
rect 21726 34076 21732 34088
rect 21784 34076 21790 34128
rect 39942 34116 39948 34128
rect 31864 34088 39948 34116
rect 17678 34008 17684 34060
rect 17736 34048 17742 34060
rect 19981 34051 20039 34057
rect 19981 34048 19993 34051
rect 17736 34020 19993 34048
rect 17736 34008 17742 34020
rect 19981 34017 19993 34020
rect 20027 34017 20039 34051
rect 31864 34048 31892 34088
rect 39942 34076 39948 34088
rect 40000 34076 40006 34128
rect 56612 34116 56640 34144
rect 56612 34088 56916 34116
rect 56888 34057 56916 34088
rect 64138 34076 64144 34128
rect 64196 34116 64202 34128
rect 90726 34116 90732 34128
rect 64196 34088 90732 34116
rect 64196 34076 64202 34088
rect 90726 34076 90732 34088
rect 90784 34076 90790 34128
rect 35989 34051 36047 34057
rect 35989 34048 36001 34051
rect 19981 34011 20039 34017
rect 22066 34020 31892 34048
rect 35912 34020 36001 34048
rect 20257 33983 20315 33989
rect 20257 33949 20269 33983
rect 20303 33980 20315 33983
rect 22066 33980 22094 34020
rect 20303 33952 22094 33980
rect 20303 33949 20315 33952
rect 20257 33943 20315 33949
rect 31110 33872 31116 33924
rect 31168 33912 31174 33924
rect 35912 33912 35940 34020
rect 35989 34017 36001 34020
rect 36035 34017 36047 34051
rect 56689 34051 56747 34057
rect 56689 34048 56701 34051
rect 35989 34011 36047 34017
rect 45526 34020 56701 34048
rect 44542 33940 44548 33992
rect 44600 33980 44606 33992
rect 45526 33980 45554 34020
rect 56689 34017 56701 34020
rect 56735 34017 56747 34051
rect 56689 34011 56747 34017
rect 56873 34051 56931 34057
rect 56873 34017 56885 34051
rect 56919 34017 56931 34051
rect 57054 34048 57060 34060
rect 57015 34020 57060 34048
rect 56873 34011 56931 34017
rect 57054 34008 57060 34020
rect 57112 34008 57118 34060
rect 57241 34051 57299 34057
rect 57241 34017 57253 34051
rect 57287 34048 57299 34051
rect 62942 34048 62948 34060
rect 57287 34020 62948 34048
rect 57287 34017 57299 34020
rect 57241 34011 57299 34017
rect 62942 34008 62948 34020
rect 63000 34048 63006 34060
rect 63402 34048 63408 34060
rect 63000 34020 63408 34048
rect 63000 34008 63006 34020
rect 63402 34008 63408 34020
rect 63460 34008 63466 34060
rect 65610 34008 65616 34060
rect 65668 34048 65674 34060
rect 74442 34048 74448 34060
rect 65668 34020 74448 34048
rect 65668 34008 65674 34020
rect 74442 34008 74448 34020
rect 74500 34008 74506 34060
rect 56962 33980 56968 33992
rect 44600 33952 45554 33980
rect 56923 33952 56968 33980
rect 44600 33940 44606 33952
rect 56962 33940 56968 33952
rect 57020 33980 57026 33992
rect 57517 33983 57575 33989
rect 57517 33980 57529 33983
rect 57020 33952 57529 33980
rect 57020 33940 57026 33952
rect 57517 33949 57529 33952
rect 57563 33949 57575 33983
rect 57517 33943 57575 33949
rect 57790 33940 57796 33992
rect 57848 33980 57854 33992
rect 92934 33980 92940 33992
rect 57848 33952 92940 33980
rect 57848 33940 57854 33952
rect 92934 33940 92940 33952
rect 92992 33940 92998 33992
rect 31168 33884 35940 33912
rect 31168 33872 31174 33884
rect 33042 33804 33048 33856
rect 33100 33844 33106 33856
rect 34514 33844 34520 33856
rect 33100 33816 34520 33844
rect 33100 33804 33106 33816
rect 34514 33804 34520 33816
rect 34572 33804 34578 33856
rect 35805 33847 35863 33853
rect 35805 33813 35817 33847
rect 35851 33844 35863 33847
rect 35912 33844 35940 33884
rect 36173 33915 36231 33921
rect 36173 33881 36185 33915
rect 36219 33912 36231 33915
rect 67818 33912 67824 33924
rect 36219 33884 67824 33912
rect 36219 33881 36231 33884
rect 36173 33875 36231 33881
rect 67818 33872 67824 33884
rect 67876 33872 67882 33924
rect 40954 33844 40960 33856
rect 35851 33816 40960 33844
rect 35851 33813 35863 33816
rect 35805 33807 35863 33813
rect 40954 33804 40960 33816
rect 41012 33804 41018 33856
rect 57422 33844 57428 33856
rect 57383 33816 57428 33844
rect 57422 33804 57428 33816
rect 57480 33804 57486 33856
rect 60001 33847 60059 33853
rect 60001 33813 60013 33847
rect 60047 33844 60059 33847
rect 60277 33847 60335 33853
rect 60277 33844 60289 33847
rect 60047 33816 60289 33844
rect 60047 33813 60059 33816
rect 60001 33807 60059 33813
rect 60277 33813 60289 33816
rect 60323 33844 60335 33847
rect 95786 33844 95792 33856
rect 60323 33816 95792 33844
rect 60323 33813 60335 33816
rect 60277 33807 60335 33813
rect 95786 33804 95792 33816
rect 95844 33804 95850 33856
rect 1104 33754 98808 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 65686 33754
rect 65738 33702 65750 33754
rect 65802 33702 65814 33754
rect 65866 33702 65878 33754
rect 65930 33702 96406 33754
rect 96458 33702 96470 33754
rect 96522 33702 96534 33754
rect 96586 33702 96598 33754
rect 96650 33702 98808 33754
rect 1104 33680 98808 33702
rect 10870 33600 10876 33652
rect 10928 33640 10934 33652
rect 90818 33640 90824 33652
rect 10928 33612 90824 33640
rect 10928 33600 10934 33612
rect 90818 33600 90824 33612
rect 90876 33600 90882 33652
rect 65426 33532 65432 33584
rect 65484 33572 65490 33584
rect 66162 33572 66168 33584
rect 65484 33544 66168 33572
rect 65484 33532 65490 33544
rect 66162 33532 66168 33544
rect 66220 33532 66226 33584
rect 9582 33464 9588 33516
rect 9640 33504 9646 33516
rect 56962 33504 56968 33516
rect 9640 33476 56968 33504
rect 9640 33464 9646 33476
rect 56962 33464 56968 33476
rect 57020 33464 57026 33516
rect 31018 33396 31024 33448
rect 31076 33436 31082 33448
rect 33042 33436 33048 33448
rect 31076 33408 33048 33436
rect 31076 33396 31082 33408
rect 33042 33396 33048 33408
rect 33100 33396 33106 33448
rect 33318 33396 33324 33448
rect 33376 33436 33382 33448
rect 40497 33439 40555 33445
rect 33376 33408 33421 33436
rect 33376 33396 33382 33408
rect 40497 33405 40509 33439
rect 40543 33436 40555 33439
rect 40773 33439 40831 33445
rect 40773 33436 40785 33439
rect 40543 33408 40785 33436
rect 40543 33405 40555 33408
rect 40497 33399 40555 33405
rect 40773 33405 40785 33408
rect 40819 33436 40831 33439
rect 97534 33436 97540 33448
rect 40819 33408 97540 33436
rect 40819 33405 40831 33408
rect 40773 33399 40831 33405
rect 97534 33396 97540 33408
rect 97592 33396 97598 33448
rect 34701 33371 34759 33377
rect 34701 33337 34713 33371
rect 34747 33368 34759 33371
rect 34747 33340 45554 33368
rect 34747 33337 34759 33340
rect 34701 33331 34759 33337
rect 31202 33260 31208 33312
rect 31260 33300 31266 33312
rect 34716 33300 34744 33331
rect 31260 33272 34744 33300
rect 45526 33300 45554 33340
rect 66254 33300 66260 33312
rect 45526 33272 66260 33300
rect 31260 33260 31266 33272
rect 66254 33260 66260 33272
rect 66312 33300 66318 33312
rect 66898 33300 66904 33312
rect 66312 33272 66904 33300
rect 66312 33260 66318 33272
rect 66898 33260 66904 33272
rect 66956 33260 66962 33312
rect 1104 33210 98808 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 50326 33210
rect 50378 33158 50390 33210
rect 50442 33158 50454 33210
rect 50506 33158 50518 33210
rect 50570 33158 81046 33210
rect 81098 33158 81110 33210
rect 81162 33158 81174 33210
rect 81226 33158 81238 33210
rect 81290 33158 98808 33210
rect 1104 33136 98808 33158
rect 31938 33056 31944 33108
rect 31996 33096 32002 33108
rect 40770 33096 40776 33108
rect 31996 33068 40776 33096
rect 31996 33056 32002 33068
rect 40770 33056 40776 33068
rect 40828 33056 40834 33108
rect 70946 33056 70952 33108
rect 71004 33096 71010 33108
rect 71314 33096 71320 33108
rect 71004 33068 71320 33096
rect 71004 33056 71010 33068
rect 71314 33056 71320 33068
rect 71372 33056 71378 33108
rect 58894 33028 58900 33040
rect 58855 33000 58900 33028
rect 58894 32988 58900 33000
rect 58952 32988 58958 33040
rect 58066 32960 58072 32972
rect 58027 32932 58072 32960
rect 58066 32920 58072 32932
rect 58124 32920 58130 32972
rect 13998 32784 14004 32836
rect 14056 32824 14062 32836
rect 34146 32824 34152 32836
rect 14056 32796 34152 32824
rect 14056 32784 14062 32796
rect 34146 32784 34152 32796
rect 34204 32784 34210 32836
rect 30377 32759 30435 32765
rect 30377 32725 30389 32759
rect 30423 32756 30435 32759
rect 30653 32759 30711 32765
rect 30653 32756 30665 32759
rect 30423 32728 30665 32756
rect 30423 32725 30435 32728
rect 30377 32719 30435 32725
rect 30653 32725 30665 32728
rect 30699 32756 30711 32759
rect 56042 32756 56048 32768
rect 30699 32728 56048 32756
rect 30699 32725 30711 32728
rect 30653 32719 30711 32725
rect 56042 32716 56048 32728
rect 56100 32716 56106 32768
rect 1104 32666 98808 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 65686 32666
rect 65738 32614 65750 32666
rect 65802 32614 65814 32666
rect 65866 32614 65878 32666
rect 65930 32614 96406 32666
rect 96458 32614 96470 32666
rect 96522 32614 96534 32666
rect 96586 32614 96598 32666
rect 96650 32614 98808 32666
rect 1104 32592 98808 32614
rect 9030 32512 9036 32564
rect 9088 32552 9094 32564
rect 10781 32555 10839 32561
rect 9088 32524 10180 32552
rect 9088 32512 9094 32524
rect 10152 32484 10180 32524
rect 10781 32521 10793 32555
rect 10827 32552 10839 32555
rect 16206 32552 16212 32564
rect 10827 32524 16212 32552
rect 10827 32521 10839 32524
rect 10781 32515 10839 32521
rect 16206 32512 16212 32524
rect 16264 32512 16270 32564
rect 30282 32552 30288 32564
rect 16546 32524 30288 32552
rect 16546 32484 16574 32524
rect 30282 32512 30288 32524
rect 30340 32512 30346 32564
rect 10152 32456 16574 32484
rect 24118 32444 24124 32496
rect 24176 32484 24182 32496
rect 91925 32487 91983 32493
rect 91925 32484 91937 32487
rect 24176 32456 91937 32484
rect 24176 32444 24182 32456
rect 91925 32453 91937 32456
rect 91971 32484 91983 32487
rect 92247 32487 92305 32493
rect 92247 32484 92259 32487
rect 91971 32456 92259 32484
rect 91971 32453 91983 32456
rect 91925 32447 91983 32453
rect 92247 32453 92259 32456
rect 92293 32453 92305 32487
rect 92382 32484 92388 32496
rect 92343 32456 92388 32484
rect 92247 32447 92305 32453
rect 92382 32444 92388 32456
rect 92440 32444 92446 32496
rect 2777 32419 2835 32425
rect 2777 32385 2789 32419
rect 2823 32416 2835 32419
rect 2823 32388 5488 32416
rect 2823 32385 2835 32388
rect 2777 32379 2835 32385
rect 3050 32348 3056 32360
rect 3011 32320 3056 32348
rect 3050 32308 3056 32320
rect 3108 32308 3114 32360
rect 5460 32348 5488 32388
rect 6362 32376 6368 32428
rect 6420 32416 6426 32428
rect 43530 32416 43536 32428
rect 6420 32388 43536 32416
rect 6420 32376 6426 32388
rect 43530 32376 43536 32388
rect 43588 32376 43594 32428
rect 47302 32376 47308 32428
rect 47360 32416 47366 32428
rect 67082 32416 67088 32428
rect 47360 32388 67088 32416
rect 47360 32376 47366 32388
rect 67082 32376 67088 32388
rect 67140 32376 67146 32428
rect 92474 32416 92480 32428
rect 92435 32388 92480 32416
rect 92474 32376 92480 32388
rect 92532 32376 92538 32428
rect 6730 32348 6736 32360
rect 5460 32320 6736 32348
rect 6730 32308 6736 32320
rect 6788 32348 6794 32360
rect 9217 32351 9275 32357
rect 9217 32348 9229 32351
rect 6788 32320 9229 32348
rect 6788 32308 6794 32320
rect 9217 32317 9229 32320
rect 9263 32317 9275 32351
rect 9217 32311 9275 32317
rect 9493 32351 9551 32357
rect 9493 32317 9505 32351
rect 9539 32348 9551 32351
rect 12158 32348 12164 32360
rect 9539 32320 12164 32348
rect 9539 32317 9551 32320
rect 9493 32311 9551 32317
rect 12158 32308 12164 32320
rect 12216 32308 12222 32360
rect 30742 32308 30748 32360
rect 30800 32348 30806 32360
rect 95050 32348 95056 32360
rect 30800 32320 95056 32348
rect 30800 32308 30806 32320
rect 95050 32308 95056 32320
rect 95108 32308 95114 32360
rect 83734 32240 83740 32292
rect 83792 32280 83798 32292
rect 92109 32283 92167 32289
rect 92109 32280 92121 32283
rect 83792 32252 92121 32280
rect 83792 32240 83798 32252
rect 92109 32249 92121 32252
rect 92155 32249 92167 32283
rect 92109 32243 92167 32249
rect 4338 32212 4344 32224
rect 4299 32184 4344 32212
rect 4338 32172 4344 32184
rect 4396 32172 4402 32224
rect 41782 32172 41788 32224
rect 41840 32212 41846 32224
rect 45002 32212 45008 32224
rect 41840 32184 45008 32212
rect 41840 32172 41846 32184
rect 45002 32172 45008 32184
rect 45060 32172 45066 32224
rect 73062 32172 73068 32224
rect 73120 32212 73126 32224
rect 88978 32212 88984 32224
rect 73120 32184 88984 32212
rect 73120 32172 73126 32184
rect 88978 32172 88984 32184
rect 89036 32172 89042 32224
rect 92750 32212 92756 32224
rect 92711 32184 92756 32212
rect 92750 32172 92756 32184
rect 92808 32172 92814 32224
rect 1104 32122 98808 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 50326 32122
rect 50378 32070 50390 32122
rect 50442 32070 50454 32122
rect 50506 32070 50518 32122
rect 50570 32070 81046 32122
rect 81098 32070 81110 32122
rect 81162 32070 81174 32122
rect 81226 32070 81238 32122
rect 81290 32070 98808 32122
rect 1104 32048 98808 32070
rect 4338 31968 4344 32020
rect 4396 32008 4402 32020
rect 12342 32008 12348 32020
rect 4396 31980 12348 32008
rect 4396 31968 4402 31980
rect 12342 31968 12348 31980
rect 12400 31968 12406 32020
rect 85022 32008 85028 32020
rect 32324 31980 85028 32008
rect 32324 31881 32352 31980
rect 85022 31968 85028 31980
rect 85080 31968 85086 32020
rect 95050 32008 95056 32020
rect 88352 31980 94636 32008
rect 95011 31980 95056 32008
rect 69842 31900 69848 31952
rect 69900 31940 69906 31952
rect 70210 31940 70216 31952
rect 69900 31912 70216 31940
rect 69900 31900 69906 31912
rect 70210 31900 70216 31912
rect 70268 31940 70274 31952
rect 88352 31940 88380 31980
rect 70268 31912 88380 31940
rect 88444 31912 93992 31940
rect 70268 31900 70274 31912
rect 32033 31875 32091 31881
rect 32033 31841 32045 31875
rect 32079 31872 32091 31875
rect 32309 31875 32367 31881
rect 32309 31872 32321 31875
rect 32079 31844 32321 31872
rect 32079 31841 32091 31844
rect 32033 31835 32091 31841
rect 32309 31841 32321 31844
rect 32355 31841 32367 31875
rect 32309 31835 32367 31841
rect 40770 31832 40776 31884
rect 40828 31872 40834 31884
rect 88444 31872 88472 31912
rect 40828 31844 88472 31872
rect 40828 31832 40834 31844
rect 88978 31832 88984 31884
rect 89036 31872 89042 31884
rect 93857 31875 93915 31881
rect 93857 31872 93869 31875
rect 89036 31844 93869 31872
rect 89036 31832 89042 31844
rect 93857 31841 93869 31844
rect 93903 31841 93915 31875
rect 93964 31872 93992 31912
rect 94038 31900 94044 31952
rect 94096 31940 94102 31952
rect 94096 31912 94268 31940
rect 94096 31900 94102 31912
rect 94240 31881 94268 31912
rect 94608 31881 94636 31980
rect 95050 31968 95056 31980
rect 95108 31968 95114 32020
rect 94225 31875 94283 31881
rect 93964 31844 94176 31872
rect 93857 31835 93915 31841
rect 39942 31764 39948 31816
rect 40000 31804 40006 31816
rect 41785 31807 41843 31813
rect 41785 31804 41797 31807
rect 40000 31776 41797 31804
rect 40000 31764 40006 31776
rect 41785 31773 41797 31776
rect 41831 31804 41843 31807
rect 41969 31807 42027 31813
rect 41969 31804 41981 31807
rect 41831 31776 41981 31804
rect 41831 31773 41843 31776
rect 41785 31767 41843 31773
rect 41969 31773 41981 31776
rect 42015 31773 42027 31807
rect 43070 31804 43076 31816
rect 43031 31776 43076 31804
rect 41969 31767 42027 31773
rect 43070 31764 43076 31776
rect 43128 31764 43134 31816
rect 43346 31804 43352 31816
rect 43307 31776 43352 31804
rect 43346 31764 43352 31776
rect 43404 31764 43410 31816
rect 44729 31807 44787 31813
rect 44729 31773 44741 31807
rect 44775 31804 44787 31807
rect 71314 31804 71320 31816
rect 44775 31776 69796 31804
rect 44775 31773 44787 31776
rect 44729 31767 44787 31773
rect 69768 31736 69796 31776
rect 70320 31776 71320 31804
rect 70320 31736 70348 31776
rect 71314 31764 71320 31776
rect 71372 31764 71378 31816
rect 92658 31764 92664 31816
rect 92716 31804 92722 31816
rect 94041 31807 94099 31813
rect 94041 31804 94053 31807
rect 92716 31776 94053 31804
rect 92716 31764 92722 31776
rect 94041 31773 94053 31776
rect 94087 31773 94099 31807
rect 94148 31804 94176 31844
rect 94225 31841 94237 31875
rect 94271 31841 94283 31875
rect 94225 31835 94283 31841
rect 94593 31875 94651 31881
rect 94593 31841 94605 31875
rect 94639 31841 94651 31875
rect 94593 31835 94651 31841
rect 94501 31807 94559 31813
rect 94501 31804 94513 31807
rect 94148 31776 94513 31804
rect 94041 31767 94099 31773
rect 94501 31773 94513 31776
rect 94547 31773 94559 31807
rect 94501 31767 94559 31773
rect 69768 31708 70348 31736
rect 63954 31628 63960 31680
rect 64012 31668 64018 31680
rect 69474 31668 69480 31680
rect 64012 31640 69480 31668
rect 64012 31628 64018 31640
rect 69474 31628 69480 31640
rect 69532 31628 69538 31680
rect 1104 31578 98808 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 65686 31578
rect 65738 31526 65750 31578
rect 65802 31526 65814 31578
rect 65866 31526 65878 31578
rect 65930 31526 96406 31578
rect 96458 31526 96470 31578
rect 96522 31526 96534 31578
rect 96586 31526 96598 31578
rect 96650 31526 98808 31578
rect 1104 31504 98808 31526
rect 64598 31464 64604 31476
rect 64559 31436 64604 31464
rect 64598 31424 64604 31436
rect 64656 31424 64662 31476
rect 67818 31424 67824 31476
rect 67876 31464 67882 31476
rect 67876 31436 70164 31464
rect 67876 31424 67882 31436
rect 64138 31356 64144 31408
rect 64196 31396 64202 31408
rect 70026 31396 70032 31408
rect 64196 31368 70032 31396
rect 64196 31356 64202 31368
rect 70026 31356 70032 31368
rect 70084 31356 70090 31408
rect 70136 31396 70164 31436
rect 70136 31368 72832 31396
rect 53834 31288 53840 31340
rect 53892 31328 53898 31340
rect 64322 31328 64328 31340
rect 53892 31300 64328 31328
rect 53892 31288 53898 31300
rect 64322 31288 64328 31300
rect 64380 31288 64386 31340
rect 68646 31288 68652 31340
rect 68704 31328 68710 31340
rect 72804 31337 72832 31368
rect 70581 31331 70639 31337
rect 70581 31328 70593 31331
rect 68704 31300 70593 31328
rect 68704 31288 68710 31300
rect 70581 31297 70593 31300
rect 70627 31297 70639 31331
rect 70581 31291 70639 31297
rect 72789 31331 72847 31337
rect 72789 31297 72801 31331
rect 72835 31297 72847 31331
rect 72789 31291 72847 31297
rect 74353 31331 74411 31337
rect 74353 31297 74365 31331
rect 74399 31328 74411 31331
rect 77846 31328 77852 31340
rect 74399 31300 77852 31328
rect 74399 31297 74411 31300
rect 74353 31291 74411 31297
rect 77846 31288 77852 31300
rect 77904 31288 77910 31340
rect 48130 31220 48136 31272
rect 48188 31260 48194 31272
rect 70305 31263 70363 31269
rect 48188 31232 64368 31260
rect 48188 31220 48194 31232
rect 34790 31152 34796 31204
rect 34848 31192 34854 31204
rect 64138 31192 64144 31204
rect 34848 31164 64144 31192
rect 34848 31152 34854 31164
rect 64138 31152 64144 31164
rect 64196 31152 64202 31204
rect 64340 31192 64368 31232
rect 70305 31229 70317 31263
rect 70351 31229 70363 31263
rect 71590 31260 71596 31272
rect 71551 31232 71596 31260
rect 70305 31223 70363 31229
rect 70320 31192 70348 31223
rect 71590 31220 71596 31232
rect 71648 31220 71654 31272
rect 72513 31263 72571 31269
rect 72513 31229 72525 31263
rect 72559 31260 72571 31263
rect 81526 31260 81532 31272
rect 72559 31232 81532 31260
rect 72559 31229 72571 31232
rect 72513 31223 72571 31229
rect 81526 31220 81532 31232
rect 81584 31220 81590 31272
rect 74353 31195 74411 31201
rect 74353 31192 74365 31195
rect 64340 31164 70348 31192
rect 70412 31164 74365 31192
rect 24210 31084 24216 31136
rect 24268 31124 24274 31136
rect 33410 31124 33416 31136
rect 24268 31096 33416 31124
rect 24268 31084 24274 31096
rect 33410 31084 33416 31096
rect 33468 31124 33474 31136
rect 63954 31124 63960 31136
rect 33468 31096 63960 31124
rect 33468 31084 33474 31096
rect 63954 31084 63960 31096
rect 64012 31084 64018 31136
rect 64046 31084 64052 31136
rect 64104 31124 64110 31136
rect 64417 31127 64475 31133
rect 64417 31124 64429 31127
rect 64104 31096 64429 31124
rect 64104 31084 64110 31096
rect 64417 31093 64429 31096
rect 64463 31124 64475 31127
rect 64598 31124 64604 31136
rect 64463 31096 64604 31124
rect 64463 31093 64475 31096
rect 64417 31087 64475 31093
rect 64598 31084 64604 31096
rect 64656 31084 64662 31136
rect 67082 31084 67088 31136
rect 67140 31124 67146 31136
rect 68738 31124 68744 31136
rect 67140 31096 68744 31124
rect 67140 31084 67146 31096
rect 68738 31084 68744 31096
rect 68796 31124 68802 31136
rect 70412 31124 70440 31164
rect 74353 31161 74365 31164
rect 74399 31161 74411 31195
rect 74353 31155 74411 31161
rect 71406 31124 71412 31136
rect 68796 31096 70440 31124
rect 71367 31096 71412 31124
rect 68796 31084 68802 31096
rect 71406 31084 71412 31096
rect 71464 31084 71470 31136
rect 1104 31034 98808 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 50326 31034
rect 50378 30982 50390 31034
rect 50442 30982 50454 31034
rect 50506 30982 50518 31034
rect 50570 30982 81046 31034
rect 81098 30982 81110 31034
rect 81162 30982 81174 31034
rect 81226 30982 81238 31034
rect 81290 30982 98808 31034
rect 1104 30960 98808 30982
rect 26510 30880 26516 30932
rect 26568 30920 26574 30932
rect 30006 30920 30012 30932
rect 26568 30892 30012 30920
rect 26568 30880 26574 30892
rect 30006 30880 30012 30892
rect 30064 30880 30070 30932
rect 31110 30880 31116 30932
rect 31168 30920 31174 30932
rect 31294 30920 31300 30932
rect 31168 30892 31300 30920
rect 31168 30880 31174 30892
rect 31294 30880 31300 30892
rect 31352 30920 31358 30932
rect 84838 30920 84844 30932
rect 31352 30892 84844 30920
rect 31352 30880 31358 30892
rect 11882 30852 11888 30864
rect 10336 30824 11888 30852
rect 9950 30784 9956 30796
rect 9911 30756 9956 30784
rect 9950 30744 9956 30756
rect 10008 30744 10014 30796
rect 10336 30793 10364 30824
rect 11882 30812 11888 30824
rect 11940 30812 11946 30864
rect 32214 30812 32220 30864
rect 32272 30852 32278 30864
rect 67910 30852 67916 30864
rect 32272 30824 67916 30852
rect 32272 30812 32278 30824
rect 67910 30812 67916 30824
rect 67968 30812 67974 30864
rect 10321 30787 10379 30793
rect 10321 30753 10333 30787
rect 10367 30753 10379 30787
rect 10321 30747 10379 30753
rect 10413 30787 10471 30793
rect 10413 30753 10425 30787
rect 10459 30784 10471 30787
rect 10594 30784 10600 30796
rect 10459 30756 10600 30784
rect 10459 30753 10471 30756
rect 10413 30747 10471 30753
rect 10594 30744 10600 30756
rect 10652 30744 10658 30796
rect 15194 30744 15200 30796
rect 15252 30784 15258 30796
rect 21085 30787 21143 30793
rect 21085 30784 21097 30787
rect 15252 30756 21097 30784
rect 15252 30744 15258 30756
rect 21085 30753 21097 30756
rect 21131 30753 21143 30787
rect 21085 30747 21143 30753
rect 64322 30744 64328 30796
rect 64380 30784 64386 30796
rect 67637 30787 67695 30793
rect 67637 30784 67649 30787
rect 64380 30756 67649 30784
rect 64380 30744 64386 30756
rect 67637 30753 67649 30756
rect 67683 30753 67695 30787
rect 67637 30747 67695 30753
rect 67818 30744 67824 30796
rect 67876 30784 67882 30796
rect 68204 30793 68232 30892
rect 84838 30880 84844 30892
rect 84896 30880 84902 30932
rect 69474 30852 69480 30864
rect 69435 30824 69480 30852
rect 69474 30812 69480 30824
rect 69532 30852 69538 30864
rect 69532 30824 70164 30852
rect 69532 30812 69538 30824
rect 68189 30787 68247 30793
rect 67876 30756 67921 30784
rect 67876 30744 67882 30756
rect 68189 30753 68201 30787
rect 68235 30753 68247 30787
rect 68189 30747 68247 30753
rect 68557 30787 68615 30793
rect 68557 30753 68569 30787
rect 68603 30784 68615 30787
rect 68646 30784 68652 30796
rect 68603 30756 68652 30784
rect 68603 30753 68615 30756
rect 68557 30747 68615 30753
rect 68646 30744 68652 30756
rect 68704 30744 68710 30796
rect 69658 30784 69664 30796
rect 69619 30756 69664 30784
rect 69658 30744 69664 30756
rect 69716 30744 69722 30796
rect 70026 30784 70032 30796
rect 69987 30756 70032 30784
rect 70026 30744 70032 30756
rect 70084 30744 70090 30796
rect 70136 30784 70164 30824
rect 70305 30787 70363 30793
rect 70305 30784 70317 30787
rect 70136 30756 70317 30784
rect 70305 30753 70317 30756
rect 70351 30753 70363 30787
rect 70305 30747 70363 30753
rect 70397 30787 70455 30793
rect 70397 30753 70409 30787
rect 70443 30784 70455 30787
rect 70486 30784 70492 30796
rect 70443 30756 70492 30784
rect 70443 30753 70455 30756
rect 70397 30747 70455 30753
rect 21358 30676 21364 30728
rect 21416 30716 21422 30728
rect 21453 30719 21511 30725
rect 21453 30716 21465 30719
rect 21416 30688 21465 30716
rect 21416 30676 21422 30688
rect 21453 30685 21465 30688
rect 21499 30685 21511 30719
rect 21453 30679 21511 30685
rect 22278 30676 22284 30728
rect 22336 30716 22342 30728
rect 68373 30719 68431 30725
rect 22336 30688 67496 30716
rect 22336 30676 22342 30688
rect 2866 30608 2872 30660
rect 2924 30648 2930 30660
rect 9766 30648 9772 30660
rect 2924 30620 6914 30648
rect 9727 30620 9772 30648
rect 2924 30608 2930 30620
rect 6886 30580 6914 30620
rect 9766 30608 9772 30620
rect 9824 30608 9830 30660
rect 67361 30651 67419 30657
rect 67361 30648 67373 30651
rect 16546 30620 67373 30648
rect 16546 30580 16574 30620
rect 67361 30617 67373 30620
rect 67407 30617 67419 30651
rect 67468 30648 67496 30688
rect 68373 30685 68385 30719
rect 68419 30716 68431 30719
rect 68738 30716 68744 30728
rect 68419 30688 68744 30716
rect 68419 30685 68431 30688
rect 68373 30679 68431 30685
rect 68738 30676 68744 30688
rect 68796 30676 68802 30728
rect 69845 30719 69903 30725
rect 69845 30716 69857 30719
rect 69584 30688 69857 30716
rect 69584 30648 69612 30688
rect 69845 30685 69857 30688
rect 69891 30685 69903 30719
rect 70320 30716 70348 30747
rect 70486 30744 70492 30756
rect 70544 30744 70550 30796
rect 92382 30716 92388 30728
rect 70320 30688 92388 30716
rect 69845 30679 69903 30685
rect 92382 30676 92388 30688
rect 92440 30676 92446 30728
rect 67468 30620 69612 30648
rect 67361 30611 67419 30617
rect 6886 30552 16574 30580
rect 67082 30540 67088 30592
rect 67140 30580 67146 30592
rect 67140 30552 67185 30580
rect 67140 30540 67146 30552
rect 70026 30540 70032 30592
rect 70084 30580 70090 30592
rect 70857 30583 70915 30589
rect 70857 30580 70869 30583
rect 70084 30552 70869 30580
rect 70084 30540 70090 30552
rect 70857 30549 70869 30552
rect 70903 30549 70915 30583
rect 70857 30543 70915 30549
rect 1104 30490 98808 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 65686 30490
rect 65738 30438 65750 30490
rect 65802 30438 65814 30490
rect 65866 30438 65878 30490
rect 65930 30438 96406 30490
rect 96458 30438 96470 30490
rect 96522 30438 96534 30490
rect 96586 30438 96598 30490
rect 96650 30438 98808 30490
rect 1104 30416 98808 30438
rect 20070 30336 20076 30388
rect 20128 30376 20134 30388
rect 67818 30376 67824 30388
rect 20128 30348 67824 30376
rect 20128 30336 20134 30348
rect 67818 30336 67824 30348
rect 67876 30336 67882 30388
rect 67910 30336 67916 30388
rect 67968 30376 67974 30388
rect 70026 30376 70032 30388
rect 67968 30348 70032 30376
rect 67968 30336 67974 30348
rect 70026 30336 70032 30348
rect 70084 30336 70090 30388
rect 81526 30336 81532 30388
rect 81584 30376 81590 30388
rect 82354 30376 82360 30388
rect 81584 30348 82360 30376
rect 81584 30336 81590 30348
rect 82354 30336 82360 30348
rect 82412 30336 82418 30388
rect 84562 30336 84568 30388
rect 84620 30376 84626 30388
rect 84838 30376 84844 30388
rect 84620 30348 84844 30376
rect 84620 30336 84626 30348
rect 84838 30336 84844 30348
rect 84896 30336 84902 30388
rect 34514 30268 34520 30320
rect 34572 30308 34578 30320
rect 43070 30308 43076 30320
rect 34572 30280 43076 30308
rect 34572 30268 34578 30280
rect 43070 30268 43076 30280
rect 43128 30308 43134 30320
rect 43714 30308 43720 30320
rect 43128 30280 43720 30308
rect 43128 30268 43134 30280
rect 43714 30268 43720 30280
rect 43772 30268 43778 30320
rect 25774 30200 25780 30252
rect 25832 30240 25838 30252
rect 77754 30240 77760 30252
rect 25832 30212 77760 30240
rect 25832 30200 25838 30212
rect 77754 30200 77760 30212
rect 77812 30200 77818 30252
rect 78490 30240 78496 30252
rect 78451 30212 78496 30240
rect 78490 30200 78496 30212
rect 78548 30200 78554 30252
rect 26050 30132 26056 30184
rect 26108 30172 26114 30184
rect 41230 30172 41236 30184
rect 26108 30144 26234 30172
rect 41191 30144 41236 30172
rect 26108 30132 26114 30144
rect 26206 30104 26234 30144
rect 41230 30132 41236 30144
rect 41288 30132 41294 30184
rect 58069 30175 58127 30181
rect 41386 30144 51074 30172
rect 41386 30104 41414 30144
rect 26206 30076 41414 30104
rect 41601 30107 41659 30113
rect 41601 30073 41613 30107
rect 41647 30073 41659 30107
rect 51046 30104 51074 30144
rect 58069 30141 58081 30175
rect 58115 30172 58127 30175
rect 58158 30172 58164 30184
rect 58115 30144 58164 30172
rect 58115 30141 58127 30144
rect 58069 30135 58127 30141
rect 58158 30132 58164 30144
rect 58216 30132 58222 30184
rect 77849 30175 77907 30181
rect 77849 30172 77861 30175
rect 74506 30144 77861 30172
rect 69750 30104 69756 30116
rect 51046 30076 69756 30104
rect 41601 30067 41659 30073
rect 26694 29996 26700 30048
rect 26752 30036 26758 30048
rect 36538 30036 36544 30048
rect 26752 30008 36544 30036
rect 26752 29996 26758 30008
rect 36538 29996 36544 30008
rect 36596 29996 36602 30048
rect 41046 29996 41052 30048
rect 41104 30036 41110 30048
rect 41616 30036 41644 30067
rect 69750 30064 69756 30076
rect 69808 30064 69814 30116
rect 41104 30008 41644 30036
rect 58253 30039 58311 30045
rect 41104 29996 41110 30008
rect 58253 30005 58265 30039
rect 58299 30036 58311 30039
rect 74506 30036 74534 30144
rect 77849 30141 77861 30144
rect 77895 30172 77907 30175
rect 86218 30172 86224 30184
rect 77895 30144 86224 30172
rect 77895 30141 77907 30144
rect 77849 30135 77907 30141
rect 86218 30132 86224 30144
rect 86276 30132 86282 30184
rect 58299 30008 74534 30036
rect 58299 30005 58311 30008
rect 58253 29999 58311 30005
rect 1104 29946 98808 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 50326 29946
rect 50378 29894 50390 29946
rect 50442 29894 50454 29946
rect 50506 29894 50518 29946
rect 50570 29894 81046 29946
rect 81098 29894 81110 29946
rect 81162 29894 81174 29946
rect 81226 29894 81238 29946
rect 81290 29894 98808 29946
rect 1104 29872 98808 29894
rect 27341 29835 27399 29841
rect 27341 29801 27353 29835
rect 27387 29832 27399 29835
rect 40034 29832 40040 29844
rect 27387 29804 40040 29832
rect 27387 29801 27399 29804
rect 27341 29795 27399 29801
rect 40034 29792 40040 29804
rect 40092 29832 40098 29844
rect 40494 29832 40500 29844
rect 40092 29804 40500 29832
rect 40092 29792 40098 29804
rect 40494 29792 40500 29804
rect 40552 29792 40558 29844
rect 46290 29792 46296 29844
rect 46348 29832 46354 29844
rect 87506 29832 87512 29844
rect 46348 29804 87512 29832
rect 46348 29792 46354 29804
rect 87506 29792 87512 29804
rect 87564 29832 87570 29844
rect 88058 29832 88064 29844
rect 87564 29804 88064 29832
rect 87564 29792 87570 29804
rect 88058 29792 88064 29804
rect 88116 29792 88122 29844
rect 88720 29804 89576 29832
rect 21266 29764 21272 29776
rect 21227 29736 21272 29764
rect 21266 29724 21272 29736
rect 21324 29724 21330 29776
rect 26142 29724 26148 29776
rect 26200 29764 26206 29776
rect 26605 29767 26663 29773
rect 26605 29764 26617 29767
rect 26200 29736 26617 29764
rect 26200 29724 26206 29736
rect 26605 29733 26617 29736
rect 26651 29733 26663 29767
rect 26605 29727 26663 29733
rect 26973 29767 27031 29773
rect 26973 29733 26985 29767
rect 27019 29764 27031 29767
rect 27249 29767 27307 29773
rect 27249 29764 27261 29767
rect 27019 29736 27261 29764
rect 27019 29733 27031 29736
rect 26973 29727 27031 29733
rect 27249 29733 27261 29736
rect 27295 29764 27307 29767
rect 48314 29764 48320 29776
rect 27295 29736 48320 29764
rect 27295 29733 27307 29736
rect 27249 29727 27307 29733
rect 48314 29724 48320 29736
rect 48372 29724 48378 29776
rect 84930 29724 84936 29776
rect 84988 29764 84994 29776
rect 88720 29764 88748 29804
rect 84988 29736 88748 29764
rect 88812 29736 89207 29764
rect 84988 29724 84994 29736
rect 16206 29656 16212 29708
rect 16264 29696 16270 29708
rect 20717 29699 20775 29705
rect 20717 29696 20729 29699
rect 16264 29668 20729 29696
rect 16264 29656 16270 29668
rect 20717 29665 20729 29668
rect 20763 29665 20775 29699
rect 21910 29696 21916 29708
rect 21871 29668 21916 29696
rect 20717 29659 20775 29665
rect 21910 29656 21916 29668
rect 21968 29656 21974 29708
rect 26421 29699 26479 29705
rect 26421 29665 26433 29699
rect 26467 29696 26479 29699
rect 26786 29696 26792 29708
rect 26467 29668 26792 29696
rect 26467 29665 26479 29668
rect 26421 29659 26479 29665
rect 26786 29656 26792 29668
rect 26844 29656 26850 29708
rect 27065 29699 27123 29705
rect 27065 29665 27077 29699
rect 27111 29696 27123 29699
rect 27341 29699 27399 29705
rect 27341 29696 27353 29699
rect 27111 29668 27353 29696
rect 27111 29665 27123 29668
rect 27065 29659 27123 29665
rect 27341 29665 27353 29668
rect 27387 29665 27399 29699
rect 27341 29659 27399 29665
rect 27709 29699 27767 29705
rect 27709 29665 27721 29699
rect 27755 29696 27767 29699
rect 27798 29696 27804 29708
rect 27755 29668 27804 29696
rect 27755 29665 27767 29668
rect 27709 29659 27767 29665
rect 26237 29631 26295 29637
rect 26237 29597 26249 29631
rect 26283 29628 26295 29631
rect 27080 29628 27108 29659
rect 27798 29656 27804 29668
rect 27856 29656 27862 29708
rect 27982 29656 27988 29708
rect 28040 29696 28046 29708
rect 88812 29705 88840 29736
rect 89179 29705 89207 29736
rect 89548 29705 89576 29804
rect 88797 29699 88855 29705
rect 88797 29696 88809 29699
rect 28040 29668 88809 29696
rect 28040 29656 28046 29668
rect 88797 29665 88809 29668
rect 88843 29665 88855 29699
rect 88797 29659 88855 29665
rect 88981 29699 89039 29705
rect 88981 29665 88993 29699
rect 89027 29665 89039 29699
rect 88981 29659 89039 29665
rect 89146 29699 89207 29705
rect 89146 29665 89158 29699
rect 89192 29668 89207 29699
rect 89533 29699 89591 29705
rect 89192 29665 89204 29668
rect 89146 29659 89204 29665
rect 89533 29665 89545 29699
rect 89579 29665 89591 29699
rect 89533 29659 89591 29665
rect 26283 29600 27108 29628
rect 27433 29631 27491 29637
rect 26283 29597 26295 29600
rect 26237 29591 26295 29597
rect 27433 29597 27445 29631
rect 27479 29628 27491 29631
rect 34698 29628 34704 29640
rect 27479 29600 34704 29628
rect 27479 29597 27491 29600
rect 27433 29591 27491 29597
rect 34698 29588 34704 29600
rect 34756 29588 34762 29640
rect 34790 29588 34796 29640
rect 34848 29628 34854 29640
rect 46658 29628 46664 29640
rect 34848 29600 46664 29628
rect 34848 29588 34854 29600
rect 46658 29588 46664 29600
rect 46716 29628 46722 29640
rect 46716 29600 80054 29628
rect 46716 29588 46722 29600
rect 26418 29520 26424 29572
rect 26476 29560 26482 29572
rect 26476 29532 28994 29560
rect 26476 29520 26482 29532
rect 22186 29492 22192 29504
rect 22147 29464 22192 29492
rect 22186 29452 22192 29464
rect 22244 29452 22250 29504
rect 22278 29452 22284 29504
rect 22336 29492 22342 29504
rect 27433 29495 27491 29501
rect 27433 29492 27445 29495
rect 22336 29464 27445 29492
rect 22336 29452 22342 29464
rect 27433 29461 27445 29464
rect 27479 29492 27491 29495
rect 27525 29495 27583 29501
rect 27525 29492 27537 29495
rect 27479 29464 27537 29492
rect 27479 29461 27491 29464
rect 27433 29455 27491 29461
rect 27525 29461 27537 29464
rect 27571 29461 27583 29495
rect 28966 29492 28994 29532
rect 45002 29520 45008 29572
rect 45060 29560 45066 29572
rect 46290 29560 46296 29572
rect 45060 29532 46296 29560
rect 45060 29520 45066 29532
rect 46290 29520 46296 29532
rect 46348 29520 46354 29572
rect 80026 29560 80054 29600
rect 88058 29588 88064 29640
rect 88116 29628 88122 29640
rect 88996 29628 89024 29659
rect 89254 29628 89260 29640
rect 88116 29600 89024 29628
rect 89215 29600 89260 29628
rect 88116 29588 88122 29600
rect 89254 29588 89260 29600
rect 89312 29588 89318 29640
rect 89349 29631 89407 29637
rect 89349 29597 89361 29631
rect 89395 29628 89407 29631
rect 96154 29628 96160 29640
rect 89395 29600 96160 29628
rect 89395 29597 89407 29600
rect 89349 29591 89407 29597
rect 89364 29560 89392 29591
rect 96154 29588 96160 29600
rect 96212 29588 96218 29640
rect 80026 29532 89392 29560
rect 46566 29492 46572 29504
rect 28966 29464 46572 29492
rect 27525 29455 27583 29461
rect 46566 29452 46572 29464
rect 46624 29452 46630 29504
rect 84102 29452 84108 29504
rect 84160 29492 84166 29504
rect 89625 29495 89683 29501
rect 89625 29492 89637 29495
rect 84160 29464 89637 29492
rect 84160 29452 84166 29464
rect 89625 29461 89637 29464
rect 89671 29461 89683 29495
rect 89625 29455 89683 29461
rect 1104 29402 98808 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 65686 29402
rect 65738 29350 65750 29402
rect 65802 29350 65814 29402
rect 65866 29350 65878 29402
rect 65930 29350 96406 29402
rect 96458 29350 96470 29402
rect 96522 29350 96534 29402
rect 96586 29350 96598 29402
rect 96650 29350 98808 29402
rect 1104 29328 98808 29350
rect 17313 29291 17371 29297
rect 17313 29257 17325 29291
rect 17359 29288 17371 29291
rect 17678 29288 17684 29300
rect 17359 29260 17684 29288
rect 17359 29257 17371 29260
rect 17313 29251 17371 29257
rect 17678 29248 17684 29260
rect 17736 29248 17742 29300
rect 25501 29291 25559 29297
rect 25501 29257 25513 29291
rect 25547 29288 25559 29291
rect 25774 29288 25780 29300
rect 25547 29260 25780 29288
rect 25547 29257 25559 29260
rect 25501 29251 25559 29257
rect 25774 29248 25780 29260
rect 25832 29248 25838 29300
rect 26234 29248 26240 29300
rect 26292 29288 26298 29300
rect 26418 29288 26424 29300
rect 26292 29260 26424 29288
rect 26292 29248 26298 29260
rect 26418 29248 26424 29260
rect 26476 29248 26482 29300
rect 26786 29248 26792 29300
rect 26844 29288 26850 29300
rect 26844 29260 36492 29288
rect 26844 29248 26850 29260
rect 22186 29180 22192 29232
rect 22244 29220 22250 29232
rect 36464 29220 36492 29260
rect 36538 29248 36544 29300
rect 36596 29288 36602 29300
rect 45002 29288 45008 29300
rect 36596 29260 45008 29288
rect 36596 29248 36602 29260
rect 45002 29248 45008 29260
rect 45060 29248 45066 29300
rect 45094 29248 45100 29300
rect 45152 29288 45158 29300
rect 45281 29291 45339 29297
rect 45281 29288 45293 29291
rect 45152 29260 45293 29288
rect 45152 29248 45158 29260
rect 45281 29257 45293 29260
rect 45327 29288 45339 29291
rect 46842 29288 46848 29300
rect 45327 29260 46848 29288
rect 45327 29257 45339 29260
rect 45281 29251 45339 29257
rect 46842 29248 46848 29260
rect 46900 29248 46906 29300
rect 78766 29288 78772 29300
rect 48286 29260 78772 29288
rect 40126 29220 40132 29232
rect 22244 29192 36400 29220
rect 36464 29192 40132 29220
rect 22244 29180 22250 29192
rect 35342 29152 35348 29164
rect 16546 29124 35348 29152
rect 14461 29087 14519 29093
rect 14461 29053 14473 29087
rect 14507 29084 14519 29087
rect 16546 29084 16574 29124
rect 35342 29112 35348 29124
rect 35400 29112 35406 29164
rect 36372 29152 36400 29192
rect 40126 29180 40132 29192
rect 40184 29180 40190 29232
rect 41230 29152 41236 29164
rect 36372 29124 41236 29152
rect 41230 29112 41236 29124
rect 41288 29112 41294 29164
rect 44913 29155 44971 29161
rect 44913 29121 44925 29155
rect 44959 29152 44971 29155
rect 46385 29155 46443 29161
rect 46385 29152 46397 29155
rect 44959 29124 46397 29152
rect 44959 29121 44971 29124
rect 44913 29115 44971 29121
rect 46385 29121 46397 29124
rect 46431 29152 46443 29155
rect 48286 29152 48314 29260
rect 78766 29248 78772 29260
rect 78824 29248 78830 29300
rect 89254 29248 89260 29300
rect 89312 29288 89318 29300
rect 90634 29288 90640 29300
rect 89312 29260 90640 29288
rect 89312 29248 89318 29260
rect 90634 29248 90640 29260
rect 90692 29248 90698 29300
rect 66990 29180 66996 29232
rect 67048 29220 67054 29232
rect 75089 29223 75147 29229
rect 75089 29220 75101 29223
rect 67048 29192 75101 29220
rect 67048 29180 67054 29192
rect 75089 29189 75101 29192
rect 75135 29189 75147 29223
rect 75089 29183 75147 29189
rect 78214 29152 78220 29164
rect 46431 29124 48314 29152
rect 55186 29124 78220 29152
rect 46431 29121 46443 29124
rect 46385 29115 46443 29121
rect 14507 29056 16574 29084
rect 17497 29087 17555 29093
rect 14507 29053 14519 29056
rect 14461 29047 14519 29053
rect 17497 29053 17509 29087
rect 17543 29084 17555 29087
rect 22278 29084 22284 29096
rect 17543 29056 22284 29084
rect 17543 29053 17555 29056
rect 17497 29047 17555 29053
rect 22278 29044 22284 29056
rect 22336 29044 22342 29096
rect 25225 29087 25283 29093
rect 25225 29053 25237 29087
rect 25271 29084 25283 29087
rect 25961 29087 26019 29093
rect 25271 29056 25912 29084
rect 25271 29053 25283 29056
rect 25225 29047 25283 29053
rect 14829 29019 14887 29025
rect 14829 28985 14841 29019
rect 14875 29016 14887 29019
rect 16206 29016 16212 29028
rect 14875 28988 16212 29016
rect 14875 28985 14887 28988
rect 14829 28979 14887 28985
rect 16206 28976 16212 28988
rect 16264 28976 16270 29028
rect 16482 28976 16488 29028
rect 16540 29016 16546 29028
rect 25682 29016 25688 29028
rect 16540 28988 25688 29016
rect 16540 28976 16546 28988
rect 25682 28976 25688 28988
rect 25740 28976 25746 29028
rect 25884 28948 25912 29056
rect 25961 29053 25973 29087
rect 26007 29053 26019 29087
rect 25961 29047 26019 29053
rect 25976 29016 26004 29047
rect 26050 29044 26056 29096
rect 26108 29084 26114 29096
rect 26108 29056 26153 29084
rect 26108 29044 26114 29056
rect 26234 29044 26240 29096
rect 26292 29084 26298 29096
rect 26329 29087 26387 29093
rect 26329 29084 26341 29087
rect 26292 29056 26341 29084
rect 26292 29044 26298 29056
rect 26329 29053 26341 29056
rect 26375 29053 26387 29087
rect 26510 29084 26516 29096
rect 26471 29056 26516 29084
rect 26329 29047 26387 29053
rect 26510 29044 26516 29056
rect 26568 29044 26574 29096
rect 26694 29084 26700 29096
rect 26655 29056 26700 29084
rect 26694 29044 26700 29056
rect 26752 29044 26758 29096
rect 43714 29044 43720 29096
rect 43772 29084 43778 29096
rect 46661 29087 46719 29093
rect 46661 29084 46673 29087
rect 43772 29056 46673 29084
rect 43772 29044 43778 29056
rect 46661 29053 46673 29056
rect 46707 29053 46719 29087
rect 46661 29047 46719 29053
rect 46842 29044 46848 29096
rect 46900 29084 46906 29096
rect 55186 29084 55214 29124
rect 78214 29112 78220 29124
rect 78272 29112 78278 29164
rect 75086 29084 75092 29096
rect 46900 29056 55214 29084
rect 75047 29056 75092 29084
rect 46900 29044 46906 29056
rect 75086 29044 75092 29056
rect 75144 29044 75150 29096
rect 34790 29016 34796 29028
rect 25976 28988 34796 29016
rect 34790 28976 34796 28988
rect 34848 28976 34854 29028
rect 44744 28988 45232 29016
rect 26050 28948 26056 28960
rect 25884 28920 26056 28948
rect 26050 28908 26056 28920
rect 26108 28908 26114 28960
rect 40034 28908 40040 28960
rect 40092 28948 40098 28960
rect 44744 28948 44772 28988
rect 40092 28920 44772 28948
rect 45204 28948 45232 28988
rect 63954 28948 63960 28960
rect 45204 28920 63960 28948
rect 40092 28908 40098 28920
rect 63954 28908 63960 28920
rect 64012 28908 64018 28960
rect 1104 28858 98808 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 50326 28858
rect 50378 28806 50390 28858
rect 50442 28806 50454 28858
rect 50506 28806 50518 28858
rect 50570 28806 81046 28858
rect 81098 28806 81110 28858
rect 81162 28806 81174 28858
rect 81226 28806 81238 28858
rect 81290 28806 98808 28858
rect 1104 28784 98808 28806
rect 53466 28704 53472 28756
rect 53524 28744 53530 28756
rect 53524 28716 63908 28744
rect 53524 28704 53530 28716
rect 15565 28679 15623 28685
rect 15565 28645 15577 28679
rect 15611 28676 15623 28679
rect 23198 28676 23204 28688
rect 15611 28648 23204 28676
rect 15611 28645 15623 28648
rect 15565 28639 15623 28645
rect 23198 28636 23204 28648
rect 23256 28636 23262 28688
rect 40126 28636 40132 28688
rect 40184 28676 40190 28688
rect 63494 28676 63500 28688
rect 40184 28648 63356 28676
rect 63455 28648 63500 28676
rect 40184 28636 40190 28648
rect 15381 28611 15439 28617
rect 15381 28577 15393 28611
rect 15427 28608 15439 28611
rect 15470 28608 15476 28620
rect 15427 28580 15476 28608
rect 15427 28577 15439 28580
rect 15381 28571 15439 28577
rect 15470 28568 15476 28580
rect 15528 28568 15534 28620
rect 15654 28608 15660 28620
rect 15615 28580 15660 28608
rect 15654 28568 15660 28580
rect 15712 28568 15718 28620
rect 60369 28611 60427 28617
rect 60369 28577 60381 28611
rect 60415 28608 60427 28611
rect 60734 28608 60740 28620
rect 60415 28580 60740 28608
rect 60415 28577 60427 28580
rect 60369 28571 60427 28577
rect 60734 28568 60740 28580
rect 60792 28608 60798 28620
rect 61286 28608 61292 28620
rect 60792 28580 61292 28608
rect 60792 28568 60798 28580
rect 61286 28568 61292 28580
rect 61344 28568 61350 28620
rect 63328 28608 63356 28648
rect 63494 28636 63500 28648
rect 63552 28636 63558 28688
rect 63880 28617 63908 28716
rect 63954 28636 63960 28688
rect 64012 28676 64018 28688
rect 91922 28676 91928 28688
rect 64012 28648 91928 28676
rect 64012 28636 64018 28648
rect 91922 28636 91928 28648
rect 91980 28636 91986 28688
rect 63681 28611 63739 28617
rect 63681 28608 63693 28611
rect 63328 28580 63693 28608
rect 63681 28577 63693 28580
rect 63727 28577 63739 28611
rect 63681 28571 63739 28577
rect 63865 28611 63923 28617
rect 63865 28577 63877 28611
rect 63911 28577 63923 28611
rect 77662 28608 77668 28620
rect 77623 28580 77668 28608
rect 63865 28571 63923 28577
rect 60642 28540 60648 28552
rect 60603 28512 60648 28540
rect 60642 28500 60648 28512
rect 60700 28500 60706 28552
rect 63696 28472 63724 28571
rect 63880 28540 63908 28571
rect 77662 28568 77668 28580
rect 77720 28568 77726 28620
rect 77938 28540 77944 28552
rect 63880 28512 76052 28540
rect 77899 28512 77944 28540
rect 76024 28472 76052 28512
rect 77938 28500 77944 28512
rect 77996 28500 78002 28552
rect 84930 28472 84936 28484
rect 63696 28444 70394 28472
rect 76024 28444 84936 28472
rect 15197 28407 15255 28413
rect 15197 28373 15209 28407
rect 15243 28404 15255 28407
rect 17862 28404 17868 28416
rect 15243 28376 17868 28404
rect 15243 28373 15255 28376
rect 15197 28367 15255 28373
rect 17862 28364 17868 28376
rect 17920 28364 17926 28416
rect 21358 28364 21364 28416
rect 21416 28404 21422 28416
rect 44634 28404 44640 28416
rect 21416 28376 44640 28404
rect 21416 28364 21422 28376
rect 44634 28364 44640 28376
rect 44692 28364 44698 28416
rect 70366 28404 70394 28444
rect 84930 28432 84936 28444
rect 84988 28432 84994 28484
rect 77662 28404 77668 28416
rect 70366 28376 77668 28404
rect 77662 28364 77668 28376
rect 77720 28364 77726 28416
rect 1104 28314 98808 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 65686 28314
rect 65738 28262 65750 28314
rect 65802 28262 65814 28314
rect 65866 28262 65878 28314
rect 65930 28262 96406 28314
rect 96458 28262 96470 28314
rect 96522 28262 96534 28314
rect 96586 28262 96598 28314
rect 96650 28262 98808 28314
rect 1104 28240 98808 28262
rect 44174 28200 44180 28212
rect 26206 28172 44180 28200
rect 8202 27956 8208 28008
rect 8260 27996 8266 28008
rect 26206 27996 26234 28172
rect 44174 28160 44180 28172
rect 44232 28200 44238 28212
rect 44232 28172 45600 28200
rect 44232 28160 44238 28172
rect 43809 28135 43867 28141
rect 43809 28132 43821 28135
rect 8260 27968 26234 27996
rect 38626 28104 43821 28132
rect 8260 27956 8266 27968
rect 9398 27888 9404 27940
rect 9456 27928 9462 27940
rect 38626 27928 38654 28104
rect 43809 28101 43821 28104
rect 43855 28101 43867 28135
rect 43809 28095 43867 28101
rect 44269 28067 44327 28073
rect 44269 28064 44281 28067
rect 43732 28036 44281 28064
rect 43732 28008 43760 28036
rect 44269 28033 44281 28036
rect 44315 28033 44327 28067
rect 44269 28027 44327 28033
rect 43533 27999 43591 28005
rect 43533 27965 43545 27999
rect 43579 27996 43591 27999
rect 43714 27996 43720 28008
rect 43579 27968 43720 27996
rect 43579 27965 43591 27968
rect 43533 27959 43591 27965
rect 43714 27956 43720 27968
rect 43772 27956 43778 28008
rect 43990 27996 43996 28008
rect 43951 27968 43996 27996
rect 43990 27956 43996 27968
rect 44048 27956 44054 28008
rect 44174 27996 44180 28008
rect 44135 27968 44180 27996
rect 44174 27956 44180 27968
rect 44232 27956 44238 28008
rect 44379 27999 44437 28005
rect 44379 27996 44391 27999
rect 44376 27965 44391 27996
rect 44425 27965 44437 27999
rect 44542 27996 44548 28008
rect 44503 27968 44548 27996
rect 44376 27959 44437 27965
rect 9456 27900 38654 27928
rect 9456 27888 9462 27900
rect 44266 27888 44272 27940
rect 44324 27928 44330 27940
rect 44376 27928 44404 27959
rect 44542 27956 44548 27968
rect 44600 27956 44606 28008
rect 44637 27931 44695 27937
rect 44637 27928 44649 27931
rect 44324 27900 44649 27928
rect 44324 27888 44330 27900
rect 44637 27897 44649 27900
rect 44683 27897 44695 27931
rect 45572 27928 45600 28172
rect 77938 28160 77944 28212
rect 77996 28200 78002 28212
rect 91646 28200 91652 28212
rect 77996 28172 91652 28200
rect 77996 28160 78002 28172
rect 91646 28160 91652 28172
rect 91704 28200 91710 28212
rect 95970 28200 95976 28212
rect 91704 28172 95976 28200
rect 91704 28160 91710 28172
rect 95970 28160 95976 28172
rect 96028 28160 96034 28212
rect 48133 28135 48191 28141
rect 48133 28101 48145 28135
rect 48179 28132 48191 28135
rect 83182 28132 83188 28144
rect 48179 28104 83188 28132
rect 48179 28101 48191 28104
rect 48133 28095 48191 28101
rect 83182 28092 83188 28104
rect 83240 28092 83246 28144
rect 55950 28064 55956 28076
rect 55911 28036 55956 28064
rect 55950 28024 55956 28036
rect 56008 28024 56014 28076
rect 74626 28064 74632 28076
rect 56060 28036 74632 28064
rect 49418 27956 49424 28008
rect 49476 27996 49482 28008
rect 55585 27999 55643 28005
rect 55585 27996 55597 27999
rect 49476 27968 55597 27996
rect 49476 27956 49482 27968
rect 55585 27965 55597 27968
rect 55631 27965 55643 27999
rect 55766 27996 55772 28008
rect 55727 27968 55772 27996
rect 55585 27959 55643 27965
rect 55766 27956 55772 27968
rect 55824 27956 55830 28008
rect 55861 27999 55919 28005
rect 55861 27965 55873 27999
rect 55907 27996 55919 27999
rect 56060 27996 56088 28036
rect 74626 28024 74632 28036
rect 74684 28024 74690 28076
rect 55907 27968 56088 27996
rect 56137 27999 56195 28005
rect 55907 27965 55919 27968
rect 55861 27959 55919 27965
rect 56137 27965 56149 27999
rect 56183 27996 56195 27999
rect 56226 27996 56232 28008
rect 56183 27968 56232 27996
rect 56183 27965 56195 27968
rect 56137 27959 56195 27965
rect 56226 27956 56232 27968
rect 56284 27956 56290 28008
rect 82081 27999 82139 28005
rect 82081 27965 82093 27999
rect 82127 27996 82139 27999
rect 82357 27999 82415 28005
rect 82357 27996 82369 27999
rect 82127 27968 82369 27996
rect 82127 27965 82139 27968
rect 82081 27959 82139 27965
rect 82357 27965 82369 27968
rect 82403 27996 82415 27999
rect 83458 27996 83464 28008
rect 82403 27968 83464 27996
rect 82403 27965 82415 27968
rect 82357 27959 82415 27965
rect 83458 27956 83464 27968
rect 83516 27956 83522 28008
rect 60642 27928 60648 27940
rect 45572 27900 60648 27928
rect 44637 27891 44695 27897
rect 8110 27820 8116 27872
rect 8168 27860 8174 27872
rect 43717 27863 43775 27869
rect 43717 27860 43729 27863
rect 8168 27832 43729 27860
rect 8168 27820 8174 27832
rect 43717 27829 43729 27832
rect 43763 27860 43775 27863
rect 44542 27860 44548 27872
rect 43763 27832 44548 27860
rect 43763 27829 43775 27832
rect 43717 27823 43775 27829
rect 44542 27820 44548 27832
rect 44600 27820 44606 27872
rect 44652 27860 44680 27891
rect 60642 27888 60648 27900
rect 60700 27888 60706 27940
rect 48133 27863 48191 27869
rect 48133 27860 48145 27863
rect 44652 27832 48145 27860
rect 48133 27829 48145 27832
rect 48179 27829 48191 27863
rect 56226 27860 56232 27872
rect 56187 27832 56232 27860
rect 48133 27823 48191 27829
rect 56226 27820 56232 27832
rect 56284 27820 56290 27872
rect 1104 27770 98808 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 50326 27770
rect 50378 27718 50390 27770
rect 50442 27718 50454 27770
rect 50506 27718 50518 27770
rect 50570 27718 81046 27770
rect 81098 27718 81110 27770
rect 81162 27718 81174 27770
rect 81226 27718 81238 27770
rect 81290 27718 98808 27770
rect 1104 27696 98808 27718
rect 2406 27616 2412 27668
rect 2464 27656 2470 27668
rect 7466 27656 7472 27668
rect 2464 27628 7472 27656
rect 2464 27616 2470 27628
rect 7466 27616 7472 27628
rect 7524 27656 7530 27668
rect 8202 27656 8208 27668
rect 7524 27628 8208 27656
rect 7524 27616 7530 27628
rect 8202 27616 8208 27628
rect 8260 27616 8266 27668
rect 28626 27616 28632 27668
rect 28684 27656 28690 27668
rect 28902 27656 28908 27668
rect 28684 27628 28908 27656
rect 28684 27616 28690 27628
rect 28902 27616 28908 27628
rect 28960 27656 28966 27668
rect 43714 27656 43720 27668
rect 28960 27628 43720 27656
rect 28960 27616 28966 27628
rect 43714 27616 43720 27628
rect 43772 27616 43778 27668
rect 56226 27616 56232 27668
rect 56284 27656 56290 27668
rect 88794 27656 88800 27668
rect 56284 27628 88800 27656
rect 56284 27616 56290 27628
rect 88794 27616 88800 27628
rect 88852 27616 88858 27668
rect 16022 27548 16028 27600
rect 16080 27588 16086 27600
rect 90174 27588 90180 27600
rect 16080 27560 90180 27588
rect 16080 27548 16086 27560
rect 90174 27548 90180 27560
rect 90232 27548 90238 27600
rect 12802 27520 12808 27532
rect 12763 27492 12808 27520
rect 12802 27480 12808 27492
rect 12860 27480 12866 27532
rect 13633 27523 13691 27529
rect 13633 27489 13645 27523
rect 13679 27520 13691 27523
rect 15470 27520 15476 27532
rect 13679 27492 15476 27520
rect 13679 27489 13691 27492
rect 13633 27483 13691 27489
rect 15470 27480 15476 27492
rect 15528 27480 15534 27532
rect 17126 27480 17132 27532
rect 17184 27520 17190 27532
rect 21726 27520 21732 27532
rect 17184 27492 21732 27520
rect 17184 27480 17190 27492
rect 21726 27480 21732 27492
rect 21784 27480 21790 27532
rect 42058 27480 42064 27532
rect 42116 27520 42122 27532
rect 42429 27523 42487 27529
rect 42429 27520 42441 27523
rect 42116 27492 42441 27520
rect 42116 27480 42122 27492
rect 42429 27489 42441 27492
rect 42475 27489 42487 27523
rect 42794 27520 42800 27532
rect 42707 27492 42800 27520
rect 42429 27483 42487 27489
rect 42794 27480 42800 27492
rect 42852 27480 42858 27532
rect 42886 27480 42892 27532
rect 42944 27520 42950 27532
rect 43073 27523 43131 27529
rect 43073 27520 43085 27523
rect 42944 27492 43085 27520
rect 42944 27480 42950 27492
rect 43073 27489 43085 27492
rect 43119 27489 43131 27523
rect 43073 27483 43131 27489
rect 43165 27523 43223 27529
rect 43165 27489 43177 27523
rect 43211 27520 43223 27523
rect 51902 27520 51908 27532
rect 43211 27492 51908 27520
rect 43211 27489 43223 27492
rect 43165 27483 43223 27489
rect 51902 27480 51908 27492
rect 51960 27480 51966 27532
rect 73338 27480 73344 27532
rect 73396 27520 73402 27532
rect 73433 27523 73491 27529
rect 73433 27520 73445 27523
rect 73396 27492 73445 27520
rect 73396 27480 73402 27492
rect 73433 27489 73445 27492
rect 73479 27489 73491 27523
rect 73433 27483 73491 27489
rect 74261 27523 74319 27529
rect 74261 27489 74273 27523
rect 74307 27520 74319 27523
rect 74442 27520 74448 27532
rect 74307 27492 74448 27520
rect 74307 27489 74319 27492
rect 74261 27483 74319 27489
rect 74442 27480 74448 27492
rect 74500 27480 74506 27532
rect 77113 27523 77171 27529
rect 77113 27489 77125 27523
rect 77159 27520 77171 27523
rect 77849 27523 77907 27529
rect 77849 27520 77861 27523
rect 77159 27492 77861 27520
rect 77159 27489 77171 27492
rect 77113 27483 77171 27489
rect 77849 27489 77861 27492
rect 77895 27489 77907 27523
rect 77849 27483 77907 27489
rect 85393 27523 85451 27529
rect 85393 27489 85405 27523
rect 85439 27520 85451 27523
rect 89622 27520 89628 27532
rect 85439 27492 89628 27520
rect 85439 27489 85451 27492
rect 85393 27483 85451 27489
rect 89622 27480 89628 27492
rect 89680 27480 89686 27532
rect 14918 27452 14924 27464
rect 14879 27424 14924 27452
rect 14918 27412 14924 27424
rect 14976 27412 14982 27464
rect 15197 27455 15255 27461
rect 15197 27421 15209 27455
rect 15243 27452 15255 27455
rect 25406 27452 25412 27464
rect 15243 27424 16574 27452
rect 25367 27424 25412 27452
rect 15243 27421 15255 27424
rect 15197 27415 15255 27421
rect 16546 27384 16574 27424
rect 25406 27412 25412 27424
rect 25464 27412 25470 27464
rect 42702 27452 42708 27464
rect 42663 27424 42708 27452
rect 42702 27412 42708 27424
rect 42760 27412 42766 27464
rect 42812 27452 42840 27480
rect 42978 27452 42984 27464
rect 42812 27424 42984 27452
rect 42978 27412 42984 27424
rect 43036 27412 43042 27464
rect 43530 27452 43536 27464
rect 43491 27424 43536 27452
rect 43530 27412 43536 27424
rect 43588 27412 43594 27464
rect 46106 27412 46112 27464
rect 46164 27452 46170 27464
rect 60182 27452 60188 27464
rect 46164 27424 60188 27452
rect 46164 27412 46170 27424
rect 60182 27412 60188 27424
rect 60240 27412 60246 27464
rect 85577 27455 85635 27461
rect 85577 27452 85589 27455
rect 74368 27424 85589 27452
rect 60274 27384 60280 27396
rect 16546 27356 60280 27384
rect 60274 27344 60280 27356
rect 60332 27344 60338 27396
rect 64690 27344 64696 27396
rect 64748 27384 64754 27396
rect 74368 27384 74396 27424
rect 85577 27421 85589 27424
rect 85623 27421 85635 27455
rect 85577 27415 85635 27421
rect 77113 27387 77171 27393
rect 77113 27384 77125 27387
rect 64748 27356 74396 27384
rect 74506 27356 77125 27384
rect 64748 27344 64754 27356
rect 16485 27319 16543 27325
rect 16485 27285 16497 27319
rect 16531 27316 16543 27319
rect 42610 27316 42616 27328
rect 16531 27288 42616 27316
rect 16531 27285 16543 27288
rect 16485 27279 16543 27285
rect 42610 27276 42616 27288
rect 42668 27276 42674 27328
rect 56594 27316 56600 27328
rect 56555 27288 56600 27316
rect 56594 27276 56600 27288
rect 56652 27316 56658 27328
rect 56689 27319 56747 27325
rect 56689 27316 56701 27319
rect 56652 27288 56701 27316
rect 56652 27276 56658 27288
rect 56689 27285 56701 27288
rect 56735 27285 56747 27319
rect 56689 27279 56747 27285
rect 70394 27276 70400 27328
rect 70452 27316 70458 27328
rect 71406 27316 71412 27328
rect 70452 27288 71412 27316
rect 70452 27276 70458 27288
rect 71406 27276 71412 27288
rect 71464 27316 71470 27328
rect 74506 27316 74534 27356
rect 77113 27353 77125 27356
rect 77159 27353 77171 27387
rect 77113 27347 77171 27353
rect 77570 27344 77576 27396
rect 77628 27384 77634 27396
rect 77665 27387 77723 27393
rect 77665 27384 77677 27387
rect 77628 27356 77677 27384
rect 77628 27344 77634 27356
rect 77665 27353 77677 27356
rect 77711 27384 77723 27387
rect 78214 27384 78220 27396
rect 77711 27356 78220 27384
rect 77711 27353 77723 27356
rect 77665 27347 77723 27353
rect 78214 27344 78220 27356
rect 78272 27344 78278 27396
rect 71464 27288 74534 27316
rect 71464 27276 71470 27288
rect 84838 27276 84844 27328
rect 84896 27316 84902 27328
rect 95234 27316 95240 27328
rect 84896 27288 95240 27316
rect 84896 27276 84902 27288
rect 95234 27276 95240 27288
rect 95292 27276 95298 27328
rect 1104 27226 98808 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 65686 27226
rect 65738 27174 65750 27226
rect 65802 27174 65814 27226
rect 65866 27174 65878 27226
rect 65930 27174 96406 27226
rect 96458 27174 96470 27226
rect 96522 27174 96534 27226
rect 96586 27174 96598 27226
rect 96650 27174 98808 27226
rect 1104 27152 98808 27174
rect 7009 27115 7067 27121
rect 7009 27081 7021 27115
rect 7055 27112 7067 27115
rect 16022 27112 16028 27124
rect 7055 27084 16028 27112
rect 7055 27081 7067 27084
rect 7009 27075 7067 27081
rect 16022 27072 16028 27084
rect 16080 27072 16086 27124
rect 84838 27112 84844 27124
rect 16132 27084 84844 27112
rect 11698 27044 11704 27056
rect 7576 27016 11704 27044
rect 7576 26985 7604 27016
rect 11698 27004 11704 27016
rect 11756 27004 11762 27056
rect 12618 27004 12624 27056
rect 12676 27044 12682 27056
rect 16132 27044 16160 27084
rect 84838 27072 84844 27084
rect 84896 27072 84902 27124
rect 86052 27084 88012 27112
rect 28902 27044 28908 27056
rect 12676 27016 16160 27044
rect 16546 27016 28908 27044
rect 12676 27004 12682 27016
rect 7561 26979 7619 26985
rect 7561 26945 7573 26979
rect 7607 26945 7619 26979
rect 16546 26976 16574 27016
rect 28902 27004 28908 27016
rect 28960 27004 28966 27056
rect 42610 27004 42616 27056
rect 42668 27044 42674 27056
rect 46106 27044 46112 27056
rect 42668 27016 46112 27044
rect 42668 27004 42674 27016
rect 46106 27004 46112 27016
rect 46164 27004 46170 27056
rect 86052 27044 86080 27084
rect 87984 27053 88012 27084
rect 87858 27047 87916 27053
rect 87858 27044 87870 27047
rect 46216 27016 86080 27044
rect 86144 27016 87870 27044
rect 7561 26939 7619 26945
rect 7852 26948 16574 26976
rect 7466 26908 7472 26920
rect 7427 26880 7472 26908
rect 7466 26868 7472 26880
rect 7524 26868 7530 26920
rect 7852 26917 7880 26948
rect 17862 26936 17868 26988
rect 17920 26976 17926 26988
rect 20349 26979 20407 26985
rect 20349 26976 20361 26979
rect 17920 26948 20361 26976
rect 17920 26936 17926 26948
rect 20349 26945 20361 26948
rect 20395 26945 20407 26979
rect 20349 26939 20407 26945
rect 20916 26948 26234 26976
rect 7837 26911 7895 26917
rect 7837 26877 7849 26911
rect 7883 26877 7895 26911
rect 7837 26871 7895 26877
rect 8021 26911 8079 26917
rect 8021 26877 8033 26911
rect 8067 26877 8079 26911
rect 8021 26871 8079 26877
rect 6733 26843 6791 26849
rect 6733 26809 6745 26843
rect 6779 26840 6791 26843
rect 8036 26840 8064 26871
rect 8110 26868 8116 26920
rect 8168 26908 8174 26920
rect 8205 26911 8263 26917
rect 8205 26908 8217 26911
rect 8168 26880 8217 26908
rect 8168 26868 8174 26880
rect 8205 26877 8217 26880
rect 8251 26877 8263 26911
rect 8205 26871 8263 26877
rect 20165 26911 20223 26917
rect 20165 26877 20177 26911
rect 20211 26877 20223 26911
rect 20530 26908 20536 26920
rect 20491 26880 20536 26908
rect 20165 26871 20223 26877
rect 12618 26840 12624 26852
rect 6779 26812 12624 26840
rect 6779 26809 6791 26812
rect 6733 26803 6791 26809
rect 12618 26800 12624 26812
rect 12676 26800 12682 26852
rect 20180 26840 20208 26871
rect 20530 26868 20536 26880
rect 20588 26868 20594 26920
rect 20916 26917 20944 26948
rect 20901 26911 20959 26917
rect 20901 26877 20913 26911
rect 20947 26877 20959 26911
rect 21082 26908 21088 26920
rect 21043 26880 21088 26908
rect 20901 26871 20959 26877
rect 21082 26868 21088 26880
rect 21140 26868 21146 26920
rect 26206 26908 26234 26948
rect 41414 26936 41420 26988
rect 41472 26976 41478 26988
rect 46216 26976 46244 27016
rect 41472 26948 46244 26976
rect 41472 26936 41478 26948
rect 46290 26936 46296 26988
rect 46348 26976 46354 26988
rect 86144 26976 86172 27016
rect 87858 27013 87870 27016
rect 87904 27044 87916 27047
rect 87969 27047 88027 27053
rect 87904 27013 87920 27044
rect 87858 27007 87920 27013
rect 87969 27013 87981 27047
rect 88015 27044 88027 27047
rect 88705 27047 88763 27053
rect 88705 27044 88717 27047
rect 88015 27016 88717 27044
rect 88015 27013 88027 27016
rect 87969 27007 88027 27013
rect 88705 27013 88717 27016
rect 88751 27013 88763 27047
rect 88705 27007 88763 27013
rect 46348 26948 86172 26976
rect 46348 26936 46354 26948
rect 87046 26936 87052 26988
rect 87104 26976 87110 26988
rect 87417 26979 87475 26985
rect 87417 26976 87429 26979
rect 87104 26948 87429 26976
rect 87104 26936 87110 26948
rect 87417 26945 87429 26948
rect 87463 26976 87475 26979
rect 87892 26976 87920 27007
rect 88521 26979 88579 26985
rect 88521 26976 88533 26979
rect 87463 26948 87828 26976
rect 87892 26948 88533 26976
rect 87463 26945 87475 26948
rect 87417 26939 87475 26945
rect 45002 26908 45008 26920
rect 26206 26880 45008 26908
rect 45002 26868 45008 26880
rect 45060 26908 45066 26920
rect 57054 26908 57060 26920
rect 45060 26880 57060 26908
rect 45060 26868 45066 26880
rect 57054 26868 57060 26880
rect 57112 26868 57118 26920
rect 65337 26911 65395 26917
rect 65337 26877 65349 26911
rect 65383 26908 65395 26911
rect 70394 26908 70400 26920
rect 65383 26880 70400 26908
rect 65383 26877 65395 26880
rect 65337 26871 65395 26877
rect 70394 26868 70400 26880
rect 70452 26868 70458 26920
rect 87509 26911 87567 26917
rect 87509 26908 87521 26911
rect 86926 26880 87521 26908
rect 21358 26840 21364 26852
rect 20180 26812 21364 26840
rect 21358 26800 21364 26812
rect 21416 26800 21422 26852
rect 21453 26843 21511 26849
rect 21453 26809 21465 26843
rect 21499 26840 21511 26843
rect 23014 26840 23020 26852
rect 21499 26812 23020 26840
rect 21499 26809 21511 26812
rect 21453 26803 21511 26809
rect 23014 26800 23020 26812
rect 23072 26800 23078 26852
rect 35342 26800 35348 26852
rect 35400 26840 35406 26852
rect 86926 26840 86954 26880
rect 87509 26877 87521 26880
rect 87555 26908 87567 26911
rect 87693 26911 87751 26917
rect 87693 26908 87705 26911
rect 87555 26880 87705 26908
rect 87555 26877 87567 26880
rect 87509 26871 87567 26877
rect 87693 26877 87705 26880
rect 87739 26877 87751 26911
rect 87800 26908 87828 26948
rect 88521 26945 88533 26948
rect 88567 26945 88579 26979
rect 88521 26939 88579 26945
rect 88032 26911 88090 26917
rect 88032 26908 88044 26911
rect 87800 26880 88044 26908
rect 87693 26871 87751 26877
rect 88032 26877 88044 26880
rect 88078 26877 88090 26911
rect 88032 26871 88090 26877
rect 35400 26812 86954 26840
rect 35400 26800 35406 26812
rect 41690 26732 41696 26784
rect 41748 26772 41754 26784
rect 46290 26772 46296 26784
rect 41748 26744 46296 26772
rect 41748 26732 41754 26744
rect 46290 26732 46296 26744
rect 46348 26732 46354 26784
rect 61562 26732 61568 26784
rect 61620 26772 61626 26784
rect 62022 26772 62028 26784
rect 61620 26744 62028 26772
rect 61620 26732 61626 26744
rect 62022 26732 62028 26744
rect 62080 26772 62086 26784
rect 65153 26775 65211 26781
rect 65153 26772 65165 26775
rect 62080 26744 65165 26772
rect 62080 26732 62086 26744
rect 65153 26741 65165 26744
rect 65199 26741 65211 26775
rect 65153 26735 65211 26741
rect 69014 26732 69020 26784
rect 69072 26772 69078 26784
rect 69750 26772 69756 26784
rect 69072 26744 69756 26772
rect 69072 26732 69078 26744
rect 69750 26732 69756 26744
rect 69808 26772 69814 26784
rect 87046 26772 87052 26784
rect 69808 26744 87052 26772
rect 69808 26732 69814 26744
rect 87046 26732 87052 26744
rect 87104 26732 87110 26784
rect 87414 26732 87420 26784
rect 87472 26772 87478 26784
rect 88337 26775 88395 26781
rect 88337 26772 88349 26775
rect 87472 26744 88349 26772
rect 87472 26732 87478 26744
rect 88337 26741 88349 26744
rect 88383 26741 88395 26775
rect 88337 26735 88395 26741
rect 1104 26682 98808 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 50326 26682
rect 50378 26630 50390 26682
rect 50442 26630 50454 26682
rect 50506 26630 50518 26682
rect 50570 26630 81046 26682
rect 81098 26630 81110 26682
rect 81162 26630 81174 26682
rect 81226 26630 81238 26682
rect 81290 26630 98808 26682
rect 1104 26608 98808 26630
rect 21726 26528 21732 26580
rect 21784 26568 21790 26580
rect 21821 26571 21879 26577
rect 21821 26568 21833 26571
rect 21784 26540 21833 26568
rect 21784 26528 21790 26540
rect 21821 26537 21833 26540
rect 21867 26537 21879 26571
rect 21821 26531 21879 26537
rect 32950 26528 32956 26580
rect 33008 26568 33014 26580
rect 40034 26568 40040 26580
rect 33008 26540 40040 26568
rect 33008 26528 33014 26540
rect 40034 26528 40040 26540
rect 40092 26568 40098 26580
rect 87414 26568 87420 26580
rect 40092 26540 87420 26568
rect 40092 26528 40098 26540
rect 87414 26528 87420 26540
rect 87472 26528 87478 26580
rect 17218 26392 17224 26444
rect 17276 26432 17282 26444
rect 20717 26435 20775 26441
rect 20717 26432 20729 26435
rect 17276 26404 20729 26432
rect 17276 26392 17282 26404
rect 20717 26401 20729 26404
rect 20763 26401 20775 26435
rect 34698 26432 34704 26444
rect 34659 26404 34704 26432
rect 20717 26395 20775 26401
rect 34698 26392 34704 26404
rect 34756 26392 34762 26444
rect 20441 26367 20499 26373
rect 20441 26333 20453 26367
rect 20487 26333 20499 26367
rect 20441 26327 20499 26333
rect 17678 26256 17684 26308
rect 17736 26296 17742 26308
rect 19426 26296 19432 26308
rect 17736 26268 19432 26296
rect 17736 26256 17742 26268
rect 19426 26256 19432 26268
rect 19484 26296 19490 26308
rect 20456 26296 20484 26327
rect 21082 26324 21088 26376
rect 21140 26364 21146 26376
rect 21140 26336 21956 26364
rect 21140 26324 21146 26336
rect 19484 26268 20484 26296
rect 19484 26256 19490 26268
rect 21928 26228 21956 26336
rect 34440 26268 34744 26296
rect 34440 26228 34468 26268
rect 21928 26200 34468 26228
rect 34514 26188 34520 26240
rect 34572 26228 34578 26240
rect 34716 26228 34744 26268
rect 42794 26256 42800 26308
rect 42852 26296 42858 26308
rect 43254 26296 43260 26308
rect 42852 26268 43260 26296
rect 42852 26256 42858 26268
rect 43254 26256 43260 26268
rect 43312 26256 43318 26308
rect 84378 26256 84384 26308
rect 84436 26296 84442 26308
rect 84749 26299 84807 26305
rect 84749 26296 84761 26299
rect 84436 26268 84761 26296
rect 84436 26256 84442 26268
rect 84749 26265 84761 26268
rect 84795 26265 84807 26299
rect 84749 26259 84807 26265
rect 95970 26256 95976 26308
rect 96028 26296 96034 26308
rect 96617 26299 96675 26305
rect 96617 26296 96629 26299
rect 96028 26268 96629 26296
rect 96028 26256 96034 26268
rect 96617 26265 96629 26268
rect 96663 26296 96675 26299
rect 96709 26299 96767 26305
rect 96709 26296 96721 26299
rect 96663 26268 96721 26296
rect 96663 26265 96675 26268
rect 96617 26259 96675 26265
rect 96709 26265 96721 26268
rect 96755 26265 96767 26299
rect 96709 26259 96767 26265
rect 72326 26228 72332 26240
rect 34572 26200 34617 26228
rect 34716 26200 72332 26228
rect 34572 26188 34578 26200
rect 72326 26188 72332 26200
rect 72384 26188 72390 26240
rect 1104 26138 98808 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 65686 26138
rect 65738 26086 65750 26138
rect 65802 26086 65814 26138
rect 65866 26086 65878 26138
rect 65930 26086 96406 26138
rect 96458 26086 96470 26138
rect 96522 26086 96534 26138
rect 96586 26086 96598 26138
rect 96650 26086 98808 26138
rect 1104 26064 98808 26086
rect 10594 25984 10600 26036
rect 10652 26024 10658 26036
rect 21082 26024 21088 26036
rect 10652 25996 21088 26024
rect 10652 25984 10658 25996
rect 21082 25984 21088 25996
rect 21140 25984 21146 26036
rect 22646 25984 22652 26036
rect 22704 26024 22710 26036
rect 43806 26024 43812 26036
rect 22704 25996 43812 26024
rect 22704 25984 22710 25996
rect 43806 25984 43812 25996
rect 43864 26024 43870 26036
rect 44082 26024 44088 26036
rect 43864 25996 44088 26024
rect 43864 25984 43870 25996
rect 44082 25984 44088 25996
rect 44140 25984 44146 26036
rect 44450 25984 44456 26036
rect 44508 26024 44514 26036
rect 69474 26024 69480 26036
rect 44508 25996 69480 26024
rect 44508 25984 44514 25996
rect 69474 25984 69480 25996
rect 69532 25984 69538 26036
rect 13262 25916 13268 25968
rect 13320 25956 13326 25968
rect 44266 25956 44272 25968
rect 13320 25928 44272 25956
rect 13320 25916 13326 25928
rect 44266 25916 44272 25928
rect 44324 25916 44330 25968
rect 57330 25956 57336 25968
rect 51046 25928 57336 25956
rect 7742 25848 7748 25900
rect 7800 25888 7806 25900
rect 51046 25888 51074 25928
rect 57330 25916 57336 25928
rect 57388 25916 57394 25968
rect 7800 25860 51074 25888
rect 7800 25848 7806 25860
rect 72786 25848 72792 25900
rect 72844 25888 72850 25900
rect 80146 25888 80152 25900
rect 72844 25860 80152 25888
rect 72844 25848 72850 25860
rect 80146 25848 80152 25860
rect 80204 25848 80210 25900
rect 2869 25823 2927 25829
rect 2869 25789 2881 25823
rect 2915 25820 2927 25823
rect 42242 25820 42248 25832
rect 2915 25792 42248 25820
rect 2915 25789 2927 25792
rect 2869 25783 2927 25789
rect 42242 25780 42248 25792
rect 42300 25780 42306 25832
rect 49145 25823 49203 25829
rect 49145 25789 49157 25823
rect 49191 25789 49203 25823
rect 49145 25783 49203 25789
rect 5902 25712 5908 25764
rect 5960 25752 5966 25764
rect 45094 25752 45100 25764
rect 5960 25724 45100 25752
rect 5960 25712 5966 25724
rect 45094 25712 45100 25724
rect 45152 25712 45158 25764
rect 49160 25752 49188 25783
rect 49602 25780 49608 25832
rect 49660 25820 49666 25832
rect 49789 25823 49847 25829
rect 49789 25820 49801 25823
rect 49660 25792 49801 25820
rect 49660 25780 49666 25792
rect 49789 25789 49801 25792
rect 49835 25789 49847 25823
rect 74994 25820 75000 25832
rect 74955 25792 75000 25820
rect 49789 25783 49847 25789
rect 74994 25780 75000 25792
rect 75052 25780 75058 25832
rect 49694 25752 49700 25764
rect 49160 25724 49700 25752
rect 49694 25712 49700 25724
rect 49752 25712 49758 25764
rect 56778 25712 56784 25764
rect 56836 25752 56842 25764
rect 73890 25752 73896 25764
rect 56836 25724 73896 25752
rect 56836 25712 56842 25724
rect 73890 25712 73896 25724
rect 73948 25712 73954 25764
rect 75825 25755 75883 25761
rect 75825 25721 75837 25755
rect 75871 25752 75883 25755
rect 75914 25752 75920 25764
rect 75871 25724 75920 25752
rect 75871 25721 75883 25724
rect 75825 25715 75883 25721
rect 75914 25712 75920 25724
rect 75972 25712 75978 25764
rect 10502 25644 10508 25696
rect 10560 25684 10566 25696
rect 66070 25684 66076 25696
rect 10560 25656 66076 25684
rect 10560 25644 10566 25656
rect 66070 25644 66076 25656
rect 66128 25644 66134 25696
rect 66254 25644 66260 25696
rect 66312 25684 66318 25696
rect 67082 25684 67088 25696
rect 66312 25656 67088 25684
rect 66312 25644 66318 25656
rect 67082 25644 67088 25656
rect 67140 25684 67146 25696
rect 92474 25684 92480 25696
rect 67140 25656 92480 25684
rect 67140 25644 67146 25656
rect 92474 25644 92480 25656
rect 92532 25644 92538 25696
rect 1104 25594 98808 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 50326 25594
rect 50378 25542 50390 25594
rect 50442 25542 50454 25594
rect 50506 25542 50518 25594
rect 50570 25542 81046 25594
rect 81098 25542 81110 25594
rect 81162 25542 81174 25594
rect 81226 25542 81238 25594
rect 81290 25542 98808 25594
rect 1104 25520 98808 25542
rect 27798 25440 27804 25492
rect 27856 25480 27862 25492
rect 39390 25480 39396 25492
rect 27856 25452 39396 25480
rect 27856 25440 27862 25452
rect 39390 25440 39396 25452
rect 39448 25440 39454 25492
rect 44082 25440 44088 25492
rect 44140 25480 44146 25492
rect 66254 25480 66260 25492
rect 44140 25452 66260 25480
rect 44140 25440 44146 25452
rect 66254 25440 66260 25452
rect 66312 25440 66318 25492
rect 71314 25440 71320 25492
rect 71372 25480 71378 25492
rect 71372 25452 80928 25480
rect 71372 25440 71378 25452
rect 35526 25372 35532 25424
rect 35584 25412 35590 25424
rect 80146 25412 80152 25424
rect 35584 25384 41414 25412
rect 80107 25384 80152 25412
rect 35584 25372 35590 25384
rect 41386 25276 41414 25384
rect 80146 25372 80152 25384
rect 80204 25412 80210 25424
rect 80204 25384 80560 25412
rect 80204 25372 80210 25384
rect 47765 25347 47823 25353
rect 47765 25313 47777 25347
rect 47811 25344 47823 25347
rect 65150 25344 65156 25356
rect 47811 25316 65156 25344
rect 47811 25313 47823 25316
rect 47765 25307 47823 25313
rect 65150 25304 65156 25316
rect 65208 25344 65214 25356
rect 80532 25353 80560 25384
rect 80900 25353 80928 25452
rect 80333 25347 80391 25353
rect 80333 25344 80345 25347
rect 65208 25316 80345 25344
rect 65208 25304 65214 25316
rect 80333 25313 80345 25316
rect 80379 25313 80391 25347
rect 80333 25307 80391 25313
rect 80516 25347 80574 25353
rect 80516 25313 80528 25347
rect 80562 25313 80574 25347
rect 80516 25307 80574 25313
rect 80885 25347 80943 25353
rect 80885 25313 80897 25347
rect 80931 25313 80943 25347
rect 80885 25307 80943 25313
rect 44358 25276 44364 25288
rect 41386 25248 44364 25276
rect 44358 25236 44364 25248
rect 44416 25276 44422 25288
rect 47949 25279 48007 25285
rect 47949 25276 47961 25279
rect 44416 25248 47961 25276
rect 44416 25236 44422 25248
rect 47949 25245 47961 25248
rect 47995 25245 48007 25279
rect 78214 25276 78220 25288
rect 78175 25248 78220 25276
rect 47949 25239 48007 25245
rect 78214 25236 78220 25248
rect 78272 25236 78278 25288
rect 78490 25276 78496 25288
rect 78451 25248 78496 25276
rect 78490 25236 78496 25248
rect 78548 25236 78554 25288
rect 80238 25236 80244 25288
rect 80296 25276 80302 25288
rect 80609 25279 80667 25285
rect 80609 25276 80621 25279
rect 80296 25248 80621 25276
rect 80296 25236 80302 25248
rect 80609 25245 80621 25248
rect 80655 25245 80667 25279
rect 80609 25239 80667 25245
rect 80701 25279 80759 25285
rect 80701 25245 80713 25279
rect 80747 25245 80759 25279
rect 80701 25239 80759 25245
rect 72326 25168 72332 25220
rect 72384 25208 72390 25220
rect 72694 25208 72700 25220
rect 72384 25180 72700 25208
rect 72384 25168 72390 25180
rect 72694 25168 72700 25180
rect 72752 25168 72758 25220
rect 80716 25208 80744 25239
rect 79152 25180 80744 25208
rect 37829 25143 37887 25149
rect 37829 25109 37841 25143
rect 37875 25140 37887 25143
rect 46842 25140 46848 25152
rect 37875 25112 46848 25140
rect 37875 25109 37887 25112
rect 37829 25103 37887 25109
rect 46842 25100 46848 25112
rect 46900 25100 46906 25152
rect 72605 25143 72663 25149
rect 72605 25109 72617 25143
rect 72651 25140 72663 25143
rect 73798 25140 73804 25152
rect 72651 25112 73804 25140
rect 72651 25109 72663 25112
rect 72605 25103 72663 25109
rect 73798 25100 73804 25112
rect 73856 25100 73862 25152
rect 75914 25100 75920 25152
rect 75972 25140 75978 25152
rect 76650 25140 76656 25152
rect 75972 25112 76656 25140
rect 75972 25100 75978 25112
rect 76650 25100 76656 25112
rect 76708 25140 76714 25152
rect 79152 25140 79180 25180
rect 79594 25140 79600 25152
rect 76708 25112 79180 25140
rect 79555 25112 79600 25140
rect 76708 25100 76714 25112
rect 79594 25100 79600 25112
rect 79652 25100 79658 25152
rect 80974 25140 80980 25152
rect 80935 25112 80980 25140
rect 80974 25100 80980 25112
rect 81032 25100 81038 25152
rect 1104 25050 98808 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 65686 25050
rect 65738 24998 65750 25050
rect 65802 24998 65814 25050
rect 65866 24998 65878 25050
rect 65930 24998 96406 25050
rect 96458 24998 96470 25050
rect 96522 24998 96534 25050
rect 96586 24998 96598 25050
rect 96650 24998 98808 25050
rect 1104 24976 98808 24998
rect 9861 24939 9919 24945
rect 9861 24905 9873 24939
rect 9907 24936 9919 24939
rect 9907 24908 10180 24936
rect 9907 24905 9919 24908
rect 9861 24899 9919 24905
rect 9950 24828 9956 24880
rect 10008 24868 10014 24880
rect 10008 24840 10053 24868
rect 10008 24828 10014 24840
rect 9401 24803 9459 24809
rect 9401 24769 9413 24803
rect 9447 24800 9459 24803
rect 10042 24800 10048 24812
rect 9447 24772 10048 24800
rect 9447 24769 9459 24772
rect 9401 24763 9459 24769
rect 10042 24760 10048 24772
rect 10100 24760 10106 24812
rect 9493 24735 9551 24741
rect 9493 24701 9505 24735
rect 9539 24701 9551 24735
rect 10152 24732 10180 24908
rect 71406 24896 71412 24948
rect 71464 24936 71470 24948
rect 72786 24936 72792 24948
rect 71464 24908 72792 24936
rect 71464 24896 71470 24908
rect 72786 24896 72792 24908
rect 72844 24896 72850 24948
rect 77018 24896 77024 24948
rect 77076 24936 77082 24948
rect 80238 24936 80244 24948
rect 77076 24908 80244 24936
rect 77076 24896 77082 24908
rect 80238 24896 80244 24908
rect 80296 24896 80302 24948
rect 16022 24828 16028 24880
rect 16080 24868 16086 24880
rect 18782 24868 18788 24880
rect 16080 24840 18788 24868
rect 16080 24828 16086 24840
rect 18782 24828 18788 24840
rect 18840 24828 18846 24880
rect 43346 24828 43352 24880
rect 43404 24868 43410 24880
rect 80974 24868 80980 24880
rect 43404 24840 80980 24868
rect 43404 24828 43410 24840
rect 80974 24828 80980 24840
rect 81032 24828 81038 24880
rect 10413 24803 10471 24809
rect 10413 24769 10425 24803
rect 10459 24800 10471 24803
rect 10502 24800 10508 24812
rect 10459 24772 10508 24800
rect 10459 24769 10471 24772
rect 10413 24763 10471 24769
rect 10502 24760 10508 24772
rect 10560 24760 10566 24812
rect 19613 24803 19671 24809
rect 19613 24769 19625 24803
rect 19659 24800 19671 24803
rect 19659 24772 20024 24800
rect 19659 24769 19671 24772
rect 19613 24763 19671 24769
rect 10152 24704 10640 24732
rect 9493 24695 9551 24701
rect 9122 24596 9128 24608
rect 9083 24568 9128 24596
rect 9122 24556 9128 24568
rect 9180 24596 9186 24608
rect 9508 24596 9536 24695
rect 10612 24608 10640 24704
rect 12710 24692 12716 24744
rect 12768 24732 12774 24744
rect 14918 24732 14924 24744
rect 12768 24704 14924 24732
rect 12768 24692 12774 24704
rect 14918 24692 14924 24704
rect 14976 24732 14982 24744
rect 19150 24732 19156 24744
rect 14976 24704 19156 24732
rect 14976 24692 14982 24704
rect 19150 24692 19156 24704
rect 19208 24732 19214 24744
rect 19426 24732 19432 24744
rect 19208 24704 19432 24732
rect 19208 24692 19214 24704
rect 19426 24692 19432 24704
rect 19484 24732 19490 24744
rect 19996 24741 20024 24772
rect 30558 24760 30564 24812
rect 30616 24800 30622 24812
rect 36078 24800 36084 24812
rect 30616 24772 36084 24800
rect 30616 24760 30622 24772
rect 36078 24760 36084 24772
rect 36136 24760 36142 24812
rect 54202 24760 54208 24812
rect 54260 24800 54266 24812
rect 54260 24772 85896 24800
rect 54260 24760 54266 24772
rect 19705 24735 19763 24741
rect 19705 24732 19717 24735
rect 19484 24704 19717 24732
rect 19484 24692 19490 24704
rect 19705 24701 19717 24704
rect 19751 24701 19763 24735
rect 19705 24695 19763 24701
rect 19981 24735 20039 24741
rect 19981 24701 19993 24735
rect 20027 24732 20039 24735
rect 20070 24732 20076 24744
rect 20027 24704 20076 24732
rect 20027 24701 20039 24704
rect 19981 24695 20039 24701
rect 20070 24692 20076 24704
rect 20128 24692 20134 24744
rect 34514 24692 34520 24744
rect 34572 24732 34578 24744
rect 35802 24732 35808 24744
rect 34572 24704 35808 24732
rect 34572 24692 34578 24704
rect 35802 24692 35808 24704
rect 35860 24732 35866 24744
rect 37093 24735 37151 24741
rect 37093 24732 37105 24735
rect 35860 24704 37105 24732
rect 35860 24692 35866 24704
rect 37093 24701 37105 24704
rect 37139 24701 37151 24735
rect 37093 24695 37151 24701
rect 59354 24692 59360 24744
rect 59412 24732 59418 24744
rect 59449 24735 59507 24741
rect 59449 24732 59461 24735
rect 59412 24704 59461 24732
rect 59412 24692 59418 24704
rect 59449 24701 59461 24704
rect 59495 24701 59507 24735
rect 59449 24695 59507 24701
rect 80790 24692 80796 24744
rect 80848 24732 80854 24744
rect 85485 24735 85543 24741
rect 85485 24732 85497 24735
rect 80848 24704 85497 24732
rect 80848 24692 80854 24704
rect 85485 24701 85497 24704
rect 85531 24701 85543 24735
rect 85485 24695 85543 24701
rect 85574 24692 85580 24744
rect 85632 24732 85638 24744
rect 85868 24741 85896 24772
rect 85669 24735 85727 24741
rect 85669 24732 85681 24735
rect 85632 24704 85681 24732
rect 85632 24692 85638 24704
rect 85669 24701 85681 24704
rect 85715 24701 85727 24735
rect 85669 24695 85727 24701
rect 85853 24735 85911 24741
rect 85853 24701 85865 24735
rect 85899 24701 85911 24735
rect 86218 24732 86224 24744
rect 86179 24704 86224 24732
rect 85853 24695 85911 24701
rect 86218 24692 86224 24704
rect 86276 24692 86282 24744
rect 86402 24732 86408 24744
rect 86363 24704 86408 24732
rect 86402 24692 86408 24704
rect 86460 24692 86466 24744
rect 36826 24667 36884 24673
rect 36826 24664 36838 24667
rect 35452 24636 36838 24664
rect 35452 24608 35480 24636
rect 36826 24633 36838 24636
rect 36872 24633 36884 24667
rect 36826 24627 36884 24633
rect 41386 24636 85528 24664
rect 10594 24596 10600 24608
rect 9180 24568 9536 24596
rect 10555 24568 10600 24596
rect 9180 24556 9186 24568
rect 10594 24556 10600 24568
rect 10652 24556 10658 24608
rect 21266 24596 21272 24608
rect 21227 24568 21272 24596
rect 21266 24556 21272 24568
rect 21324 24556 21330 24608
rect 35434 24596 35440 24608
rect 35395 24568 35440 24596
rect 35434 24556 35440 24568
rect 35492 24556 35498 24608
rect 35710 24596 35716 24608
rect 35671 24568 35716 24596
rect 35710 24556 35716 24568
rect 35768 24556 35774 24608
rect 36078 24556 36084 24608
rect 36136 24596 36142 24608
rect 41386 24596 41414 24636
rect 36136 24568 41414 24596
rect 36136 24556 36142 24568
rect 85206 24556 85212 24608
rect 85264 24596 85270 24608
rect 85301 24599 85359 24605
rect 85301 24596 85313 24599
rect 85264 24568 85313 24596
rect 85264 24556 85270 24568
rect 85301 24565 85313 24568
rect 85347 24596 85359 24599
rect 85390 24596 85396 24608
rect 85347 24568 85396 24596
rect 85347 24565 85359 24568
rect 85301 24559 85359 24565
rect 85390 24556 85396 24568
rect 85448 24556 85454 24608
rect 85500 24596 85528 24636
rect 86681 24599 86739 24605
rect 86681 24596 86693 24599
rect 85500 24568 86693 24596
rect 86681 24565 86693 24568
rect 86727 24565 86739 24599
rect 86681 24559 86739 24565
rect 1104 24506 98808 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 50326 24506
rect 50378 24454 50390 24506
rect 50442 24454 50454 24506
rect 50506 24454 50518 24506
rect 50570 24454 81046 24506
rect 81098 24454 81110 24506
rect 81162 24454 81174 24506
rect 81226 24454 81238 24506
rect 81290 24454 98808 24506
rect 1104 24432 98808 24454
rect 9122 24352 9128 24404
rect 9180 24392 9186 24404
rect 41414 24392 41420 24404
rect 9180 24364 41420 24392
rect 9180 24352 9186 24364
rect 41414 24352 41420 24364
rect 41472 24352 41478 24404
rect 21266 24284 21272 24336
rect 21324 24324 21330 24336
rect 36630 24324 36636 24336
rect 21324 24296 36636 24324
rect 21324 24284 21330 24296
rect 36630 24284 36636 24296
rect 36688 24284 36694 24336
rect 9950 24216 9956 24268
rect 10008 24256 10014 24268
rect 35342 24256 35348 24268
rect 10008 24228 35348 24256
rect 10008 24216 10014 24228
rect 35342 24216 35348 24228
rect 35400 24216 35406 24268
rect 36630 24148 36636 24200
rect 36688 24188 36694 24200
rect 52270 24188 52276 24200
rect 36688 24160 52276 24188
rect 36688 24148 36694 24160
rect 52270 24148 52276 24160
rect 52328 24148 52334 24200
rect 11054 24080 11060 24132
rect 11112 24120 11118 24132
rect 11790 24120 11796 24132
rect 11112 24092 11796 24120
rect 11112 24080 11118 24092
rect 11790 24080 11796 24092
rect 11848 24120 11854 24132
rect 31386 24120 31392 24132
rect 11848 24092 31392 24120
rect 11848 24080 11854 24092
rect 31386 24080 31392 24092
rect 31444 24080 31450 24132
rect 40954 24080 40960 24132
rect 41012 24120 41018 24132
rect 64966 24120 64972 24132
rect 41012 24092 64972 24120
rect 41012 24080 41018 24092
rect 64966 24080 64972 24092
rect 65024 24080 65030 24132
rect 20070 24012 20076 24064
rect 20128 24052 20134 24064
rect 80054 24052 80060 24064
rect 20128 24024 80060 24052
rect 20128 24012 20134 24024
rect 80054 24012 80060 24024
rect 80112 24012 80118 24064
rect 1104 23962 98808 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 65686 23962
rect 65738 23910 65750 23962
rect 65802 23910 65814 23962
rect 65866 23910 65878 23962
rect 65930 23910 96406 23962
rect 96458 23910 96470 23962
rect 96522 23910 96534 23962
rect 96586 23910 96598 23962
rect 96650 23910 98808 23962
rect 1104 23888 98808 23910
rect 9766 23808 9772 23860
rect 9824 23848 9830 23860
rect 85206 23848 85212 23860
rect 9824 23820 85212 23848
rect 9824 23808 9830 23820
rect 85206 23808 85212 23820
rect 85264 23808 85270 23860
rect 10594 23740 10600 23792
rect 10652 23780 10658 23792
rect 41690 23780 41696 23792
rect 10652 23752 41696 23780
rect 10652 23740 10658 23752
rect 41690 23740 41696 23752
rect 41748 23740 41754 23792
rect 42242 23740 42248 23792
rect 42300 23780 42306 23792
rect 49418 23780 49424 23792
rect 42300 23752 49424 23780
rect 42300 23740 42306 23752
rect 49418 23740 49424 23752
rect 49476 23740 49482 23792
rect 5718 23672 5724 23724
rect 5776 23712 5782 23724
rect 6825 23715 6883 23721
rect 6825 23712 6837 23715
rect 5776 23684 6837 23712
rect 5776 23672 5782 23684
rect 6825 23681 6837 23684
rect 6871 23712 6883 23715
rect 12710 23712 12716 23724
rect 6871 23684 12716 23712
rect 6871 23681 6883 23684
rect 6825 23675 6883 23681
rect 12710 23672 12716 23684
rect 12768 23672 12774 23724
rect 40310 23672 40316 23724
rect 40368 23712 40374 23724
rect 40773 23715 40831 23721
rect 40773 23712 40785 23715
rect 40368 23684 40785 23712
rect 40368 23672 40374 23684
rect 40773 23681 40785 23684
rect 40819 23681 40831 23715
rect 40773 23675 40831 23681
rect 66898 23672 66904 23724
rect 66956 23712 66962 23724
rect 66956 23684 77616 23712
rect 66956 23672 66962 23684
rect 7101 23647 7159 23653
rect 7101 23613 7113 23647
rect 7147 23644 7159 23647
rect 31662 23644 31668 23656
rect 7147 23616 31668 23644
rect 7147 23613 7159 23616
rect 7101 23607 7159 23613
rect 31662 23604 31668 23616
rect 31720 23604 31726 23656
rect 40034 23644 40040 23656
rect 39995 23616 40040 23644
rect 40034 23604 40040 23616
rect 40092 23604 40098 23656
rect 77588 23653 77616 23684
rect 77389 23647 77447 23653
rect 77389 23613 77401 23647
rect 77435 23613 77447 23647
rect 77389 23607 77447 23613
rect 77573 23647 77631 23653
rect 77573 23613 77585 23647
rect 77619 23613 77631 23647
rect 77573 23607 77631 23613
rect 77665 23647 77723 23653
rect 77665 23613 77677 23647
rect 77711 23644 77723 23647
rect 77846 23644 77852 23656
rect 77711 23616 77852 23644
rect 77711 23613 77723 23616
rect 77665 23607 77723 23613
rect 8481 23579 8539 23585
rect 8481 23545 8493 23579
rect 8527 23576 8539 23579
rect 11054 23576 11060 23588
rect 8527 23548 11060 23576
rect 8527 23545 8539 23548
rect 8481 23539 8539 23545
rect 11054 23536 11060 23548
rect 11112 23536 11118 23588
rect 49234 23536 49240 23588
rect 49292 23576 49298 23588
rect 77205 23579 77263 23585
rect 77205 23576 77217 23579
rect 49292 23548 77217 23576
rect 49292 23536 49298 23548
rect 77205 23545 77217 23548
rect 77251 23545 77263 23579
rect 77205 23539 77263 23545
rect 48958 23468 48964 23520
rect 49016 23508 49022 23520
rect 49510 23508 49516 23520
rect 49016 23480 49516 23508
rect 49016 23468 49022 23480
rect 49510 23468 49516 23480
rect 49568 23508 49574 23520
rect 72878 23508 72884 23520
rect 49568 23480 72884 23508
rect 49568 23468 49574 23480
rect 72878 23468 72884 23480
rect 72936 23508 72942 23520
rect 76929 23511 76987 23517
rect 76929 23508 76941 23511
rect 72936 23480 76941 23508
rect 72936 23468 72942 23480
rect 76929 23477 76941 23480
rect 76975 23508 76987 23511
rect 77404 23508 77432 23607
rect 77846 23604 77852 23616
rect 77904 23604 77910 23656
rect 76975 23480 77432 23508
rect 76975 23477 76987 23480
rect 76929 23471 76987 23477
rect 1104 23418 98808 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 50326 23418
rect 50378 23366 50390 23418
rect 50442 23366 50454 23418
rect 50506 23366 50518 23418
rect 50570 23366 81046 23418
rect 81098 23366 81110 23418
rect 81162 23366 81174 23418
rect 81226 23366 81238 23418
rect 81290 23366 98808 23418
rect 1104 23344 98808 23366
rect 16114 23264 16120 23316
rect 16172 23304 16178 23316
rect 78766 23304 78772 23316
rect 16172 23276 78772 23304
rect 16172 23264 16178 23276
rect 78766 23264 78772 23276
rect 78824 23264 78830 23316
rect 44542 23196 44548 23248
rect 44600 23236 44606 23248
rect 59357 23239 59415 23245
rect 44600 23208 59308 23236
rect 44600 23196 44606 23208
rect 16390 23128 16396 23180
rect 16448 23168 16454 23180
rect 59280 23168 59308 23208
rect 59357 23205 59369 23239
rect 59403 23236 59415 23239
rect 59541 23239 59599 23245
rect 59541 23236 59553 23239
rect 59403 23208 59553 23236
rect 59403 23205 59415 23208
rect 59357 23199 59415 23205
rect 59541 23205 59553 23208
rect 59587 23236 59599 23239
rect 59587 23208 60136 23236
rect 59587 23205 59599 23208
rect 59541 23199 59599 23205
rect 59722 23168 59728 23180
rect 16448 23140 55214 23168
rect 59280 23140 59728 23168
rect 16448 23128 16454 23140
rect 29546 23060 29552 23112
rect 29604 23100 29610 23112
rect 46014 23100 46020 23112
rect 29604 23072 46020 23100
rect 29604 23060 29610 23072
rect 46014 23060 46020 23072
rect 46072 23060 46078 23112
rect 55186 23100 55214 23140
rect 59722 23128 59728 23140
rect 59780 23168 59786 23180
rect 59817 23171 59875 23177
rect 59817 23168 59829 23171
rect 59780 23140 59829 23168
rect 59780 23128 59786 23140
rect 59817 23137 59829 23140
rect 59863 23137 59875 23171
rect 59817 23131 59875 23137
rect 60001 23171 60059 23177
rect 60001 23137 60013 23171
rect 60047 23137 60059 23171
rect 60001 23131 60059 23137
rect 60016 23100 60044 23131
rect 60108 23112 60136 23208
rect 60200 23208 60504 23236
rect 60200 23177 60228 23208
rect 60185 23171 60243 23177
rect 60185 23137 60197 23171
rect 60231 23137 60243 23171
rect 60366 23168 60372 23180
rect 60327 23140 60372 23168
rect 60185 23131 60243 23137
rect 60366 23128 60372 23140
rect 60424 23128 60430 23180
rect 60476 23168 60504 23208
rect 60734 23168 60740 23180
rect 60476 23140 60740 23168
rect 60734 23128 60740 23140
rect 60792 23168 60798 23180
rect 61562 23168 61568 23180
rect 60792 23140 61568 23168
rect 60792 23128 60798 23140
rect 61562 23128 61568 23140
rect 61620 23128 61626 23180
rect 77665 23171 77723 23177
rect 77665 23137 77677 23171
rect 77711 23168 77723 23171
rect 78214 23168 78220 23180
rect 77711 23140 78220 23168
rect 77711 23137 77723 23140
rect 77665 23131 77723 23137
rect 78214 23128 78220 23140
rect 78272 23168 78278 23180
rect 90174 23168 90180 23180
rect 78272 23140 90180 23168
rect 78272 23128 78278 23140
rect 90174 23128 90180 23140
rect 90232 23128 90238 23180
rect 55186 23072 60044 23100
rect 60090 23060 60096 23112
rect 60148 23100 60154 23112
rect 61381 23103 61439 23109
rect 61381 23100 61393 23103
rect 60148 23072 60193 23100
rect 60292 23072 61393 23100
rect 60148 23060 60154 23072
rect 3418 22992 3424 23044
rect 3476 23032 3482 23044
rect 35434 23032 35440 23044
rect 3476 23004 35440 23032
rect 3476 22992 3482 23004
rect 35434 22992 35440 23004
rect 35492 22992 35498 23044
rect 43714 22992 43720 23044
rect 43772 23032 43778 23044
rect 59265 23035 59323 23041
rect 59265 23032 59277 23035
rect 43772 23004 59277 23032
rect 43772 22992 43778 23004
rect 59265 23001 59277 23004
rect 59311 23001 59323 23035
rect 60292 23032 60320 23072
rect 61381 23069 61393 23072
rect 61427 23069 61439 23103
rect 77938 23100 77944 23112
rect 77899 23072 77944 23100
rect 61381 23063 61439 23069
rect 77938 23060 77944 23072
rect 77996 23060 78002 23112
rect 59265 22995 59323 23001
rect 59372 23004 60320 23032
rect 60553 23035 60611 23041
rect 20073 22967 20131 22973
rect 20073 22933 20085 22967
rect 20119 22964 20131 22967
rect 20349 22967 20407 22973
rect 20349 22964 20361 22967
rect 20119 22936 20361 22964
rect 20119 22933 20131 22936
rect 20073 22927 20131 22933
rect 20349 22933 20361 22936
rect 20395 22964 20407 22967
rect 59372 22964 59400 23004
rect 60553 23001 60565 23035
rect 60599 23032 60611 23035
rect 72050 23032 72056 23044
rect 60599 23004 72056 23032
rect 60599 23001 60611 23004
rect 60553 22995 60611 23001
rect 72050 22992 72056 23004
rect 72108 22992 72114 23044
rect 78968 23004 93854 23032
rect 59722 22964 59728 22976
rect 20395 22936 59400 22964
rect 59683 22936 59728 22964
rect 20395 22933 20407 22936
rect 20349 22927 20407 22933
rect 59722 22924 59728 22936
rect 59780 22924 59786 22976
rect 61381 22967 61439 22973
rect 61381 22933 61393 22967
rect 61427 22964 61439 22967
rect 78968 22964 78996 23004
rect 61427 22936 78996 22964
rect 79229 22967 79287 22973
rect 61427 22933 61439 22936
rect 61381 22927 61439 22933
rect 79229 22933 79241 22967
rect 79275 22964 79287 22967
rect 79410 22964 79416 22976
rect 79275 22936 79416 22964
rect 79275 22933 79287 22936
rect 79229 22927 79287 22933
rect 79410 22924 79416 22936
rect 79468 22924 79474 22976
rect 84933 22967 84991 22973
rect 84933 22933 84945 22967
rect 84979 22964 84991 22967
rect 85114 22964 85120 22976
rect 84979 22936 85120 22964
rect 84979 22933 84991 22936
rect 84933 22927 84991 22933
rect 85114 22924 85120 22936
rect 85172 22924 85178 22976
rect 93826 22964 93854 23004
rect 95878 22964 95884 22976
rect 93826 22936 95884 22964
rect 95878 22924 95884 22936
rect 95936 22924 95942 22976
rect 1104 22874 98808 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 65686 22874
rect 65738 22822 65750 22874
rect 65802 22822 65814 22874
rect 65866 22822 65878 22874
rect 65930 22822 96406 22874
rect 96458 22822 96470 22874
rect 96522 22822 96534 22874
rect 96586 22822 96598 22874
rect 96650 22822 98808 22874
rect 1104 22800 98808 22822
rect 6362 22720 6368 22772
rect 6420 22760 6426 22772
rect 66990 22760 66996 22772
rect 6420 22732 66996 22760
rect 6420 22720 6426 22732
rect 66990 22720 66996 22732
rect 67048 22720 67054 22772
rect 49510 22652 49516 22704
rect 49568 22692 49574 22704
rect 79502 22692 79508 22704
rect 49568 22664 79508 22692
rect 49568 22652 49574 22664
rect 79502 22652 79508 22664
rect 79560 22652 79566 22704
rect 15102 22584 15108 22636
rect 15160 22624 15166 22636
rect 57514 22624 57520 22636
rect 15160 22596 57520 22624
rect 15160 22584 15166 22596
rect 57514 22584 57520 22596
rect 57572 22584 57578 22636
rect 19150 22556 19156 22568
rect 19111 22528 19156 22556
rect 19150 22516 19156 22528
rect 19208 22516 19214 22568
rect 19426 22556 19432 22568
rect 19387 22528 19432 22556
rect 19426 22516 19432 22528
rect 19484 22516 19490 22568
rect 38473 22559 38531 22565
rect 38473 22525 38485 22559
rect 38519 22556 38531 22559
rect 45465 22559 45523 22565
rect 38519 22528 41414 22556
rect 38519 22525 38531 22528
rect 38473 22519 38531 22525
rect 20809 22491 20867 22497
rect 20809 22457 20821 22491
rect 20855 22488 20867 22491
rect 22094 22488 22100 22500
rect 20855 22460 22100 22488
rect 20855 22457 20867 22460
rect 20809 22451 20867 22457
rect 22094 22448 22100 22460
rect 22152 22488 22158 22500
rect 23106 22488 23112 22500
rect 22152 22460 23112 22488
rect 22152 22448 22158 22460
rect 23106 22448 23112 22460
rect 23164 22448 23170 22500
rect 41386 22488 41414 22528
rect 45465 22525 45477 22559
rect 45511 22556 45523 22559
rect 48866 22556 48872 22568
rect 45511 22528 48872 22556
rect 45511 22525 45523 22528
rect 45465 22519 45523 22525
rect 48866 22516 48872 22528
rect 48924 22516 48930 22568
rect 47578 22488 47584 22500
rect 41386 22460 47584 22488
rect 47578 22448 47584 22460
rect 47636 22448 47642 22500
rect 48314 22448 48320 22500
rect 48372 22488 48378 22500
rect 79410 22488 79416 22500
rect 48372 22460 79416 22488
rect 48372 22448 48378 22460
rect 79410 22448 79416 22460
rect 79468 22448 79474 22500
rect 1104 22330 98808 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 50326 22330
rect 50378 22278 50390 22330
rect 50442 22278 50454 22330
rect 50506 22278 50518 22330
rect 50570 22278 81046 22330
rect 81098 22278 81110 22330
rect 81162 22278 81174 22330
rect 81226 22278 81238 22330
rect 81290 22278 98808 22330
rect 1104 22256 98808 22278
rect 19426 22176 19432 22228
rect 19484 22216 19490 22228
rect 61838 22216 61844 22228
rect 19484 22188 61844 22216
rect 19484 22176 19490 22188
rect 61838 22176 61844 22188
rect 61896 22176 61902 22228
rect 36170 22148 36176 22160
rect 36131 22120 36176 22148
rect 36170 22108 36176 22120
rect 36228 22108 36234 22160
rect 65518 22108 65524 22160
rect 65576 22148 65582 22160
rect 72234 22148 72240 22160
rect 65576 22120 72240 22148
rect 65576 22108 65582 22120
rect 72234 22108 72240 22120
rect 72292 22108 72298 22160
rect 76558 22108 76564 22160
rect 76616 22148 76622 22160
rect 83001 22151 83059 22157
rect 83001 22148 83013 22151
rect 76616 22120 83013 22148
rect 76616 22108 76622 22120
rect 83001 22117 83013 22120
rect 83047 22117 83059 22151
rect 83001 22111 83059 22117
rect 36906 22080 36912 22092
rect 36867 22052 36912 22080
rect 36906 22040 36912 22052
rect 36964 22040 36970 22092
rect 47489 22083 47547 22089
rect 47489 22049 47501 22083
rect 47535 22080 47547 22083
rect 47535 22052 47716 22080
rect 47535 22049 47547 22052
rect 47489 22043 47547 22049
rect 36078 21972 36084 22024
rect 36136 22012 36142 22024
rect 43070 22012 43076 22024
rect 36136 21984 43076 22012
rect 36136 21972 36142 21984
rect 43070 21972 43076 21984
rect 43128 21972 43134 22024
rect 47394 21972 47400 22024
rect 47452 22012 47458 22024
rect 47581 22015 47639 22021
rect 47581 22012 47593 22015
rect 47452 21984 47593 22012
rect 47452 21972 47458 21984
rect 47581 21981 47593 21984
rect 47627 21981 47639 22015
rect 47688 22012 47716 22052
rect 47946 22040 47952 22092
rect 48004 22080 48010 22092
rect 71130 22080 71136 22092
rect 48004 22052 71136 22080
rect 48004 22040 48010 22052
rect 71130 22040 71136 22052
rect 71188 22040 71194 22092
rect 47857 22015 47915 22021
rect 47857 22012 47869 22015
rect 47688 21984 47869 22012
rect 47581 21975 47639 21981
rect 47857 21981 47869 21984
rect 47903 22012 47915 22015
rect 88150 22012 88156 22024
rect 47903 21984 88156 22012
rect 47903 21981 47915 21984
rect 47857 21975 47915 21981
rect 88150 21972 88156 21984
rect 88208 21972 88214 22024
rect 33778 21904 33784 21956
rect 33836 21944 33842 21956
rect 34330 21944 34336 21956
rect 33836 21916 34336 21944
rect 33836 21904 33842 21916
rect 34330 21904 34336 21916
rect 34388 21944 34394 21956
rect 34388 21916 41414 21944
rect 34388 21904 34394 21916
rect 26786 21836 26792 21888
rect 26844 21876 26850 21888
rect 35618 21876 35624 21888
rect 26844 21848 35624 21876
rect 26844 21836 26850 21848
rect 35618 21836 35624 21848
rect 35676 21836 35682 21888
rect 41386 21876 41414 21916
rect 50062 21904 50068 21956
rect 50120 21944 50126 21956
rect 64414 21944 64420 21956
rect 50120 21916 64420 21944
rect 50120 21904 50126 21916
rect 64414 21904 64420 21916
rect 64472 21904 64478 21956
rect 48961 21879 49019 21885
rect 48961 21876 48973 21879
rect 41386 21848 48973 21876
rect 48961 21845 48973 21848
rect 49007 21845 49019 21879
rect 48961 21839 49019 21845
rect 63034 21836 63040 21888
rect 63092 21876 63098 21888
rect 83093 21879 83151 21885
rect 83093 21876 83105 21879
rect 63092 21848 83105 21876
rect 63092 21836 63098 21848
rect 83093 21845 83105 21848
rect 83139 21845 83151 21879
rect 83093 21839 83151 21845
rect 1104 21786 98808 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 65686 21786
rect 65738 21734 65750 21786
rect 65802 21734 65814 21786
rect 65866 21734 65878 21786
rect 65930 21734 96406 21786
rect 96458 21734 96470 21786
rect 96522 21734 96534 21786
rect 96586 21734 96598 21786
rect 96650 21734 98808 21786
rect 1104 21712 98808 21734
rect 11974 21632 11980 21684
rect 12032 21672 12038 21684
rect 28810 21672 28816 21684
rect 12032 21644 28816 21672
rect 12032 21632 12038 21644
rect 28810 21632 28816 21644
rect 28868 21632 28874 21684
rect 35342 21632 35348 21684
rect 35400 21672 35406 21684
rect 35710 21672 35716 21684
rect 35400 21644 35716 21672
rect 35400 21632 35406 21644
rect 35710 21632 35716 21644
rect 35768 21672 35774 21684
rect 36008 21675 36066 21681
rect 36008 21672 36020 21675
rect 35768 21644 36020 21672
rect 35768 21632 35774 21644
rect 36008 21641 36020 21644
rect 36054 21641 36066 21675
rect 36008 21635 36066 21641
rect 43714 21632 43720 21684
rect 43772 21672 43778 21684
rect 69566 21672 69572 21684
rect 43772 21644 69572 21672
rect 43772 21632 43778 21644
rect 69566 21632 69572 21644
rect 69624 21632 69630 21684
rect 22370 21564 22376 21616
rect 22428 21604 22434 21616
rect 22830 21604 22836 21616
rect 22428 21576 22836 21604
rect 22428 21564 22434 21576
rect 22830 21564 22836 21576
rect 22888 21604 22894 21616
rect 35897 21607 35955 21613
rect 35897 21604 35909 21607
rect 22888 21576 35909 21604
rect 22888 21564 22894 21576
rect 35897 21573 35909 21576
rect 35943 21573 35955 21607
rect 35897 21567 35955 21573
rect 48866 21564 48872 21616
rect 48924 21604 48930 21616
rect 76558 21604 76564 21616
rect 48924 21576 76564 21604
rect 48924 21564 48930 21576
rect 76558 21564 76564 21576
rect 76616 21564 76622 21616
rect 76926 21564 76932 21616
rect 76984 21604 76990 21616
rect 76984 21576 81388 21604
rect 76984 21564 76990 21576
rect 15378 21496 15384 21548
rect 15436 21536 15442 21548
rect 28258 21536 28264 21548
rect 15436 21508 28264 21536
rect 15436 21496 15442 21508
rect 28258 21496 28264 21508
rect 28316 21496 28322 21548
rect 28350 21496 28356 21548
rect 28408 21536 28414 21548
rect 35805 21539 35863 21545
rect 35805 21536 35817 21539
rect 28408 21508 35817 21536
rect 28408 21496 28414 21508
rect 35805 21505 35817 21508
rect 35851 21536 35863 21539
rect 64506 21536 64512 21548
rect 35851 21508 64512 21536
rect 35851 21505 35863 21508
rect 35805 21499 35863 21505
rect 64506 21496 64512 21508
rect 64564 21496 64570 21548
rect 76742 21496 76748 21548
rect 76800 21536 76806 21548
rect 76800 21508 81020 21536
rect 76800 21496 76806 21508
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 26786 21468 26792 21480
rect 12768 21440 26792 21468
rect 12768 21428 12774 21440
rect 26786 21428 26792 21440
rect 26844 21428 26850 21480
rect 26970 21428 26976 21480
rect 27028 21468 27034 21480
rect 33870 21468 33876 21480
rect 27028 21440 33876 21468
rect 27028 21428 27034 21440
rect 33870 21428 33876 21440
rect 33928 21428 33934 21480
rect 80606 21468 80612 21480
rect 80567 21440 80612 21468
rect 80606 21428 80612 21440
rect 80664 21428 80670 21480
rect 80790 21468 80796 21480
rect 80751 21440 80796 21468
rect 80790 21428 80796 21440
rect 80848 21428 80854 21480
rect 80992 21477 81020 21508
rect 81360 21477 81388 21576
rect 80977 21471 81035 21477
rect 80977 21437 80989 21471
rect 81023 21437 81035 21471
rect 80977 21431 81035 21437
rect 81253 21471 81311 21477
rect 81253 21437 81265 21471
rect 81299 21437 81311 21471
rect 81253 21431 81311 21437
rect 81345 21471 81403 21477
rect 81345 21437 81357 21471
rect 81391 21437 81403 21471
rect 81345 21431 81403 21437
rect 1670 21360 1676 21412
rect 1728 21400 1734 21412
rect 28626 21400 28632 21412
rect 1728 21372 28632 21400
rect 1728 21360 1734 21372
rect 28626 21360 28632 21372
rect 28684 21360 28690 21412
rect 33962 21360 33968 21412
rect 34020 21400 34026 21412
rect 35437 21403 35495 21409
rect 35437 21400 35449 21403
rect 34020 21372 35449 21400
rect 34020 21360 34026 21372
rect 35437 21369 35449 21372
rect 35483 21369 35495 21403
rect 36173 21403 36231 21409
rect 36173 21400 36185 21403
rect 35437 21363 35495 21369
rect 35866 21372 36185 21400
rect 35345 21335 35403 21341
rect 35345 21301 35357 21335
rect 35391 21332 35403 21335
rect 35618 21332 35624 21344
rect 35391 21304 35624 21332
rect 35391 21301 35403 21304
rect 35345 21295 35403 21301
rect 35618 21292 35624 21304
rect 35676 21332 35682 21344
rect 35866 21332 35894 21372
rect 36173 21369 36185 21372
rect 36219 21400 36231 21403
rect 56134 21400 56140 21412
rect 36219 21372 56140 21400
rect 36219 21369 36231 21372
rect 36173 21363 36231 21369
rect 56134 21360 56140 21372
rect 56192 21360 56198 21412
rect 58986 21360 58992 21412
rect 59044 21400 59050 21412
rect 81268 21400 81296 21431
rect 59044 21372 81296 21400
rect 59044 21360 59050 21372
rect 35676 21304 35894 21332
rect 35676 21292 35682 21304
rect 57146 21292 57152 21344
rect 57204 21332 57210 21344
rect 81805 21335 81863 21341
rect 81805 21332 81817 21335
rect 57204 21304 81817 21332
rect 57204 21292 57210 21304
rect 81805 21301 81817 21304
rect 81851 21301 81863 21335
rect 81805 21295 81863 21301
rect 1104 21242 98808 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 50326 21242
rect 50378 21190 50390 21242
rect 50442 21190 50454 21242
rect 50506 21190 50518 21242
rect 50570 21190 81046 21242
rect 81098 21190 81110 21242
rect 81162 21190 81174 21242
rect 81226 21190 81238 21242
rect 81290 21190 98808 21242
rect 1104 21168 98808 21190
rect 77662 21088 77668 21140
rect 77720 21088 77726 21140
rect 97166 21128 97172 21140
rect 80026 21100 97172 21128
rect 77680 21060 77708 21088
rect 77941 21063 77999 21069
rect 77941 21060 77953 21063
rect 77680 21032 77953 21060
rect 77941 21029 77953 21032
rect 77987 21029 77999 21063
rect 77941 21023 77999 21029
rect 77662 20992 77668 21004
rect 77623 20964 77668 20992
rect 77662 20952 77668 20964
rect 77720 20992 77726 21004
rect 80026 20992 80054 21100
rect 97166 21088 97172 21100
rect 97224 21088 97230 21140
rect 77720 20964 80054 20992
rect 77720 20952 77726 20964
rect 90174 20952 90180 21004
rect 90232 20992 90238 21004
rect 94317 20995 94375 21001
rect 94317 20992 94329 20995
rect 90232 20964 94329 20992
rect 90232 20952 90238 20964
rect 94317 20961 94329 20964
rect 94363 20961 94375 20995
rect 94317 20955 94375 20961
rect 94593 20927 94651 20933
rect 94593 20924 94605 20927
rect 94332 20896 94605 20924
rect 94332 20856 94360 20896
rect 94593 20893 94605 20896
rect 94639 20893 94651 20927
rect 94593 20887 94651 20893
rect 94148 20828 94360 20856
rect 20714 20748 20720 20800
rect 20772 20788 20778 20800
rect 21910 20788 21916 20800
rect 20772 20760 21916 20788
rect 20772 20748 20778 20760
rect 21910 20748 21916 20760
rect 21968 20788 21974 20800
rect 50062 20788 50068 20800
rect 21968 20760 50068 20788
rect 21968 20748 21974 20760
rect 50062 20748 50068 20760
rect 50120 20748 50126 20800
rect 71314 20748 71320 20800
rect 71372 20788 71378 20800
rect 94148 20797 94176 20828
rect 94133 20791 94191 20797
rect 94133 20788 94145 20791
rect 71372 20760 94145 20788
rect 71372 20748 71378 20760
rect 94133 20757 94145 20760
rect 94179 20757 94191 20791
rect 94133 20751 94191 20757
rect 95234 20748 95240 20800
rect 95292 20788 95298 20800
rect 95697 20791 95755 20797
rect 95697 20788 95709 20791
rect 95292 20760 95709 20788
rect 95292 20748 95298 20760
rect 95697 20757 95709 20760
rect 95743 20757 95755 20791
rect 95697 20751 95755 20757
rect 1104 20698 98808 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 65686 20698
rect 65738 20646 65750 20698
rect 65802 20646 65814 20698
rect 65866 20646 65878 20698
rect 65930 20646 96406 20698
rect 96458 20646 96470 20698
rect 96522 20646 96534 20698
rect 96586 20646 96598 20698
rect 96650 20646 98808 20698
rect 1104 20624 98808 20646
rect 21910 20544 21916 20596
rect 21968 20584 21974 20596
rect 24210 20584 24216 20596
rect 21968 20556 24216 20584
rect 21968 20544 21974 20556
rect 24210 20544 24216 20556
rect 24268 20544 24274 20596
rect 64230 20544 64236 20596
rect 64288 20584 64294 20596
rect 66254 20584 66260 20596
rect 64288 20556 66260 20584
rect 64288 20544 64294 20556
rect 66254 20544 66260 20556
rect 66312 20544 66318 20596
rect 10778 20476 10784 20528
rect 10836 20516 10842 20528
rect 10836 20488 24164 20516
rect 10836 20476 10842 20488
rect 3605 20383 3663 20389
rect 3605 20349 3617 20383
rect 3651 20380 3663 20383
rect 4798 20380 4804 20392
rect 3651 20352 4804 20380
rect 3651 20349 3663 20352
rect 3605 20343 3663 20349
rect 4798 20340 4804 20352
rect 4856 20380 4862 20392
rect 5258 20380 5264 20392
rect 4856 20352 5264 20380
rect 4856 20340 4862 20352
rect 5258 20340 5264 20352
rect 5316 20340 5322 20392
rect 15838 20340 15844 20392
rect 15896 20380 15902 20392
rect 19426 20380 19432 20392
rect 15896 20352 19432 20380
rect 15896 20340 15902 20352
rect 19426 20340 19432 20352
rect 19484 20380 19490 20392
rect 19521 20383 19579 20389
rect 19521 20380 19533 20383
rect 19484 20352 19533 20380
rect 19484 20340 19490 20352
rect 19521 20349 19533 20352
rect 19567 20349 19579 20383
rect 23934 20380 23940 20392
rect 23895 20352 23940 20380
rect 19521 20343 19579 20349
rect 23934 20340 23940 20352
rect 23992 20340 23998 20392
rect 24136 20389 24164 20488
rect 24302 20448 24308 20460
rect 24263 20420 24308 20448
rect 24302 20408 24308 20420
rect 24360 20408 24366 20460
rect 30190 20448 30196 20460
rect 24412 20420 30196 20448
rect 24120 20383 24178 20389
rect 24120 20349 24132 20383
rect 24166 20349 24178 20383
rect 24120 20343 24178 20349
rect 24210 20340 24216 20392
rect 24268 20380 24274 20392
rect 24412 20380 24440 20420
rect 30190 20408 30196 20420
rect 30248 20408 30254 20460
rect 51261 20451 51319 20457
rect 51261 20417 51273 20451
rect 51307 20448 51319 20451
rect 88426 20448 88432 20460
rect 51307 20420 88432 20448
rect 51307 20417 51319 20420
rect 51261 20411 51319 20417
rect 88426 20408 88432 20420
rect 88484 20408 88490 20460
rect 24268 20352 24440 20380
rect 24268 20340 24274 20352
rect 24486 20340 24492 20392
rect 24544 20380 24550 20392
rect 24854 20380 24860 20392
rect 24544 20352 24860 20380
rect 24544 20340 24550 20352
rect 24854 20340 24860 20352
rect 24912 20340 24918 20392
rect 50985 20383 51043 20389
rect 50985 20349 50997 20383
rect 51031 20380 51043 20383
rect 55030 20380 55036 20392
rect 51031 20352 55036 20380
rect 51031 20349 51043 20352
rect 50985 20343 51043 20349
rect 55030 20340 55036 20352
rect 55088 20340 55094 20392
rect 78122 20380 78128 20392
rect 78083 20352 78128 20380
rect 78122 20340 78128 20352
rect 78180 20340 78186 20392
rect 19797 20315 19855 20321
rect 19797 20281 19809 20315
rect 19843 20312 19855 20315
rect 45278 20312 45284 20324
rect 19843 20284 45284 20312
rect 19843 20281 19855 20284
rect 19797 20275 19855 20281
rect 45278 20272 45284 20284
rect 45336 20272 45342 20324
rect 3789 20247 3847 20253
rect 3789 20213 3801 20247
rect 3835 20244 3847 20247
rect 12802 20244 12808 20256
rect 3835 20216 12808 20244
rect 3835 20213 3847 20216
rect 3789 20207 3847 20213
rect 12802 20204 12808 20216
rect 12860 20204 12866 20256
rect 23845 20247 23903 20253
rect 23845 20213 23857 20247
rect 23891 20244 23903 20247
rect 24486 20244 24492 20256
rect 23891 20216 24492 20244
rect 23891 20213 23903 20216
rect 23845 20207 23903 20213
rect 24486 20204 24492 20216
rect 24544 20204 24550 20256
rect 24581 20247 24639 20253
rect 24581 20213 24593 20247
rect 24627 20244 24639 20247
rect 28166 20244 28172 20256
rect 24627 20216 28172 20244
rect 24627 20213 24639 20216
rect 24581 20207 24639 20213
rect 28166 20204 28172 20216
rect 28224 20204 28230 20256
rect 43622 20204 43628 20256
rect 43680 20244 43686 20256
rect 52365 20247 52423 20253
rect 52365 20244 52377 20247
rect 43680 20216 52377 20244
rect 43680 20204 43686 20216
rect 52365 20213 52377 20216
rect 52411 20213 52423 20247
rect 52365 20207 52423 20213
rect 62850 20204 62856 20256
rect 62908 20244 62914 20256
rect 74166 20244 74172 20256
rect 62908 20216 74172 20244
rect 62908 20204 62914 20216
rect 74166 20204 74172 20216
rect 74224 20204 74230 20256
rect 1104 20154 98808 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 50326 20154
rect 50378 20102 50390 20154
rect 50442 20102 50454 20154
rect 50506 20102 50518 20154
rect 50570 20102 81046 20154
rect 81098 20102 81110 20154
rect 81162 20102 81174 20154
rect 81226 20102 81238 20154
rect 81290 20102 98808 20154
rect 1104 20080 98808 20102
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 24302 20040 24308 20052
rect 16172 20012 24308 20040
rect 16172 20000 16178 20012
rect 24302 20000 24308 20012
rect 24360 20000 24366 20052
rect 65150 20040 65156 20052
rect 65111 20012 65156 20040
rect 65150 20000 65156 20012
rect 65208 20000 65214 20052
rect 71682 20000 71688 20052
rect 71740 20040 71746 20052
rect 95234 20040 95240 20052
rect 71740 20012 95240 20040
rect 71740 20000 71746 20012
rect 95234 20000 95240 20012
rect 95292 20000 95298 20052
rect 19058 19932 19064 19984
rect 19116 19972 19122 19984
rect 24210 19972 24216 19984
rect 19116 19944 24216 19972
rect 19116 19932 19122 19944
rect 24210 19932 24216 19944
rect 24268 19932 24274 19984
rect 24854 19932 24860 19984
rect 24912 19972 24918 19984
rect 25866 19972 25872 19984
rect 24912 19944 25872 19972
rect 24912 19932 24918 19944
rect 25866 19932 25872 19944
rect 25924 19972 25930 19984
rect 62206 19972 62212 19984
rect 25924 19944 62212 19972
rect 25924 19932 25930 19944
rect 62206 19932 62212 19944
rect 62264 19932 62270 19984
rect 64690 19932 64696 19984
rect 64748 19972 64754 19984
rect 83642 19972 83648 19984
rect 64748 19944 83648 19972
rect 64748 19932 64754 19944
rect 83642 19932 83648 19944
rect 83700 19932 83706 19984
rect 88794 19972 88800 19984
rect 88755 19944 88800 19972
rect 88794 19932 88800 19944
rect 88852 19972 88858 19984
rect 88852 19944 89714 19972
rect 88852 19932 88858 19944
rect 28166 19864 28172 19916
rect 28224 19904 28230 19916
rect 61746 19904 61752 19916
rect 28224 19876 61752 19904
rect 28224 19864 28230 19876
rect 61746 19864 61752 19876
rect 61804 19864 61810 19916
rect 64966 19904 64972 19916
rect 64927 19876 64972 19904
rect 64966 19864 64972 19876
rect 65024 19864 65030 19916
rect 68370 19864 68376 19916
rect 68428 19904 68434 19916
rect 72421 19907 72479 19913
rect 72421 19904 72433 19907
rect 68428 19876 72433 19904
rect 68428 19864 68434 19876
rect 72421 19873 72433 19876
rect 72467 19873 72479 19907
rect 72878 19904 72884 19916
rect 72839 19876 72884 19904
rect 72421 19867 72479 19873
rect 72878 19864 72884 19876
rect 72936 19864 72942 19916
rect 73065 19907 73123 19913
rect 73065 19873 73077 19907
rect 73111 19873 73123 19907
rect 73246 19904 73252 19916
rect 73207 19876 73252 19904
rect 73065 19867 73123 19873
rect 45278 19796 45284 19848
rect 45336 19836 45342 19848
rect 50890 19836 50896 19848
rect 45336 19808 50896 19836
rect 45336 19796 45342 19808
rect 50890 19796 50896 19808
rect 50948 19836 50954 19848
rect 73080 19836 73108 19867
rect 73246 19864 73252 19876
rect 73304 19864 73310 19916
rect 82630 19864 82636 19916
rect 82688 19904 82694 19916
rect 85850 19904 85856 19916
rect 82688 19876 85856 19904
rect 82688 19864 82694 19876
rect 85850 19864 85856 19876
rect 85908 19864 85914 19916
rect 89686 19904 89714 19944
rect 90361 19907 90419 19913
rect 90361 19904 90373 19907
rect 89686 19876 90373 19904
rect 90361 19873 90373 19876
rect 90407 19873 90419 19907
rect 90361 19867 90419 19873
rect 90542 19864 90548 19916
rect 90600 19904 90606 19916
rect 91097 19907 91155 19913
rect 91097 19904 91109 19907
rect 90600 19876 91109 19904
rect 90600 19864 90606 19876
rect 91097 19873 91109 19876
rect 91143 19873 91155 19907
rect 91097 19867 91155 19873
rect 50948 19808 73108 19836
rect 50948 19796 50954 19808
rect 90174 19796 90180 19848
rect 90232 19836 90238 19848
rect 90450 19836 90456 19848
rect 90232 19808 90456 19836
rect 90232 19796 90238 19808
rect 90450 19796 90456 19808
rect 90508 19836 90514 19848
rect 90637 19839 90695 19845
rect 90637 19836 90649 19839
rect 90508 19808 90649 19836
rect 90508 19796 90514 19808
rect 90637 19805 90649 19808
rect 90683 19805 90695 19839
rect 90637 19799 90695 19805
rect 56134 19728 56140 19780
rect 56192 19768 56198 19780
rect 89073 19771 89131 19777
rect 89073 19768 89085 19771
rect 56192 19740 69520 19768
rect 56192 19728 56198 19740
rect 43070 19660 43076 19712
rect 43128 19700 43134 19712
rect 46106 19700 46112 19712
rect 43128 19672 46112 19700
rect 43128 19660 43134 19672
rect 46106 19660 46112 19672
rect 46164 19660 46170 19712
rect 69492 19700 69520 19740
rect 80026 19740 89085 19768
rect 80026 19700 80054 19740
rect 89073 19737 89085 19740
rect 89119 19737 89131 19771
rect 89073 19731 89131 19737
rect 69492 19672 80054 19700
rect 89622 19660 89628 19712
rect 89680 19700 89686 19712
rect 91281 19703 91339 19709
rect 91281 19700 91293 19703
rect 89680 19672 91293 19700
rect 89680 19660 89686 19672
rect 91281 19669 91293 19672
rect 91327 19669 91339 19703
rect 91281 19663 91339 19669
rect 1104 19610 98808 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 65686 19610
rect 65738 19558 65750 19610
rect 65802 19558 65814 19610
rect 65866 19558 65878 19610
rect 65930 19558 96406 19610
rect 96458 19558 96470 19610
rect 96522 19558 96534 19610
rect 96586 19558 96598 19610
rect 96650 19558 98808 19610
rect 1104 19536 98808 19558
rect 43070 19496 43076 19508
rect 22066 19468 43076 19496
rect 8938 19320 8944 19372
rect 8996 19360 9002 19372
rect 22066 19360 22094 19468
rect 43070 19456 43076 19468
rect 43128 19456 43134 19508
rect 44542 19388 44548 19440
rect 44600 19428 44606 19440
rect 44600 19400 44863 19428
rect 44600 19388 44606 19400
rect 8996 19332 22094 19360
rect 8996 19320 9002 19332
rect 44450 19320 44456 19372
rect 44508 19360 44514 19372
rect 44835 19360 44863 19400
rect 44913 19363 44971 19369
rect 44508 19332 44588 19360
rect 44835 19332 44864 19360
rect 44508 19320 44514 19332
rect 4985 19295 5043 19301
rect 4985 19261 4997 19295
rect 5031 19292 5043 19295
rect 12250 19292 12256 19304
rect 5031 19264 12256 19292
rect 5031 19261 5043 19264
rect 4985 19255 5043 19261
rect 12250 19252 12256 19264
rect 12308 19252 12314 19304
rect 20990 19252 20996 19304
rect 21048 19292 21054 19304
rect 24118 19292 24124 19304
rect 21048 19264 24124 19292
rect 21048 19252 21054 19264
rect 24118 19252 24124 19264
rect 24176 19252 24182 19304
rect 43162 19252 43168 19304
rect 43220 19292 43226 19304
rect 44560 19292 44588 19332
rect 43220 19264 44588 19292
rect 43220 19252 43226 19264
rect 44634 19252 44640 19304
rect 44692 19292 44698 19304
rect 44836 19301 44864 19332
rect 44913 19329 44925 19363
rect 44959 19360 44971 19363
rect 45094 19360 45100 19372
rect 44959 19332 45100 19360
rect 44959 19329 44971 19332
rect 44913 19323 44971 19329
rect 45094 19320 45100 19332
rect 45152 19320 45158 19372
rect 45370 19320 45376 19372
rect 45428 19320 45434 19372
rect 46106 19320 46112 19372
rect 46164 19360 46170 19372
rect 71682 19360 71688 19372
rect 46164 19332 71688 19360
rect 46164 19320 46170 19332
rect 71682 19320 71688 19332
rect 71740 19320 71746 19372
rect 44820 19295 44878 19301
rect 44820 19292 44832 19295
rect 44692 19264 44737 19292
rect 44799 19264 44832 19292
rect 44692 19252 44698 19264
rect 44820 19261 44832 19264
rect 44866 19261 44878 19295
rect 44820 19255 44878 19261
rect 45002 19252 45008 19304
rect 45060 19292 45066 19304
rect 45060 19264 45105 19292
rect 45060 19252 45066 19264
rect 45186 19252 45192 19304
rect 45244 19292 45250 19304
rect 45388 19292 45416 19320
rect 48225 19295 48283 19301
rect 48225 19292 48237 19295
rect 45244 19264 45289 19292
rect 45388 19264 48237 19292
rect 45244 19252 45250 19264
rect 48225 19261 48237 19264
rect 48271 19261 48283 19295
rect 48225 19255 48283 19261
rect 50065 19295 50123 19301
rect 50065 19261 50077 19295
rect 50111 19261 50123 19295
rect 50614 19292 50620 19304
rect 50575 19264 50620 19292
rect 50065 19255 50123 19261
rect 5537 19227 5595 19233
rect 5537 19193 5549 19227
rect 5583 19224 5595 19227
rect 50080 19224 50108 19255
rect 50614 19252 50620 19264
rect 50672 19252 50678 19304
rect 67634 19292 67640 19304
rect 57946 19264 67640 19292
rect 57946 19224 57974 19264
rect 67634 19252 67640 19264
rect 67692 19252 67698 19304
rect 5583 19196 45416 19224
rect 5583 19193 5595 19196
rect 5537 19187 5595 19193
rect 28534 19116 28540 19168
rect 28592 19156 28598 19168
rect 45281 19159 45339 19165
rect 45281 19156 45293 19159
rect 28592 19128 45293 19156
rect 28592 19116 28598 19128
rect 45281 19125 45293 19128
rect 45327 19125 45339 19159
rect 45388 19156 45416 19196
rect 46860 19196 57974 19224
rect 46860 19156 46888 19196
rect 62114 19184 62120 19236
rect 62172 19224 62178 19236
rect 62758 19224 62764 19236
rect 62172 19196 62764 19224
rect 62172 19184 62178 19196
rect 62758 19184 62764 19196
rect 62816 19224 62822 19236
rect 86862 19224 86868 19236
rect 62816 19196 86868 19224
rect 62816 19184 62822 19196
rect 86862 19184 86868 19196
rect 86920 19184 86926 19236
rect 95234 19224 95240 19236
rect 89686 19196 95240 19224
rect 45388 19128 46888 19156
rect 48225 19159 48283 19165
rect 45281 19119 45339 19125
rect 48225 19125 48237 19159
rect 48271 19156 48283 19159
rect 50154 19156 50160 19168
rect 48271 19128 50160 19156
rect 48271 19125 48283 19128
rect 48225 19119 48283 19125
rect 50154 19116 50160 19128
rect 50212 19116 50218 19168
rect 50614 19116 50620 19168
rect 50672 19156 50678 19168
rect 54110 19156 54116 19168
rect 50672 19128 54116 19156
rect 50672 19116 50678 19128
rect 54110 19116 54116 19128
rect 54168 19116 54174 19168
rect 73430 19116 73436 19168
rect 73488 19156 73494 19168
rect 89686 19156 89714 19196
rect 95234 19184 95240 19196
rect 95292 19184 95298 19236
rect 73488 19128 89714 19156
rect 73488 19116 73494 19128
rect 90634 19116 90640 19168
rect 90692 19156 90698 19168
rect 97258 19156 97264 19168
rect 90692 19128 97264 19156
rect 90692 19116 90698 19128
rect 97258 19116 97264 19128
rect 97316 19116 97322 19168
rect 1104 19066 98808 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 50326 19066
rect 50378 19014 50390 19066
rect 50442 19014 50454 19066
rect 50506 19014 50518 19066
rect 50570 19014 81046 19066
rect 81098 19014 81110 19066
rect 81162 19014 81174 19066
rect 81226 19014 81238 19066
rect 81290 19014 98808 19066
rect 1104 18992 98808 19014
rect 3970 18912 3976 18964
rect 4028 18952 4034 18964
rect 65153 18955 65211 18961
rect 4028 18924 64828 18952
rect 4028 18912 4034 18924
rect 28994 18844 29000 18896
rect 29052 18884 29058 18896
rect 29730 18884 29736 18896
rect 29052 18856 29736 18884
rect 29052 18844 29058 18856
rect 29730 18844 29736 18856
rect 29788 18884 29794 18896
rect 45186 18884 45192 18896
rect 29788 18856 45192 18884
rect 29788 18844 29794 18856
rect 45186 18844 45192 18856
rect 45244 18844 45250 18896
rect 49053 18887 49111 18893
rect 49053 18853 49065 18887
rect 49099 18884 49111 18887
rect 53374 18884 53380 18896
rect 49099 18856 53380 18884
rect 49099 18853 49111 18856
rect 49053 18847 49111 18853
rect 53374 18844 53380 18856
rect 53432 18844 53438 18896
rect 62942 18844 62948 18896
rect 63000 18884 63006 18896
rect 63402 18884 63408 18896
rect 63000 18856 63408 18884
rect 63000 18844 63006 18856
rect 63402 18844 63408 18856
rect 63460 18884 63466 18896
rect 64800 18893 64828 18924
rect 65153 18921 65165 18955
rect 65199 18952 65211 18955
rect 65426 18952 65432 18964
rect 65199 18924 65432 18952
rect 65199 18921 65211 18924
rect 65153 18915 65211 18921
rect 65426 18912 65432 18924
rect 65484 18912 65490 18964
rect 96154 18912 96160 18964
rect 96212 18952 96218 18964
rect 96212 18924 97672 18952
rect 96212 18912 96218 18924
rect 63589 18887 63647 18893
rect 63589 18884 63601 18887
rect 63460 18856 63601 18884
rect 63460 18844 63466 18856
rect 63589 18853 63601 18856
rect 63635 18853 63647 18887
rect 63589 18847 63647 18853
rect 64785 18887 64843 18893
rect 64785 18853 64797 18887
rect 64831 18853 64843 18887
rect 64785 18847 64843 18853
rect 64874 18844 64880 18896
rect 64932 18884 64938 18896
rect 65245 18887 65303 18893
rect 65245 18884 65257 18887
rect 64932 18856 65257 18884
rect 64932 18844 64938 18856
rect 65245 18853 65257 18856
rect 65291 18853 65303 18887
rect 65245 18847 65303 18853
rect 70578 18844 70584 18896
rect 70636 18884 70642 18896
rect 73430 18884 73436 18896
rect 70636 18856 73436 18884
rect 70636 18844 70642 18856
rect 73430 18844 73436 18856
rect 73488 18844 73494 18896
rect 79410 18844 79416 18896
rect 79468 18884 79474 18896
rect 79468 18856 97580 18884
rect 79468 18844 79474 18856
rect 39482 18776 39488 18828
rect 39540 18816 39546 18828
rect 47213 18819 47271 18825
rect 47213 18816 47225 18819
rect 39540 18788 47225 18816
rect 39540 18776 39546 18788
rect 47213 18785 47225 18788
rect 47259 18816 47271 18819
rect 47673 18819 47731 18825
rect 47673 18816 47685 18819
rect 47259 18788 47685 18816
rect 47259 18785 47271 18788
rect 47213 18779 47271 18785
rect 47673 18785 47685 18788
rect 47719 18785 47731 18819
rect 47673 18779 47731 18785
rect 57422 18776 57428 18828
rect 57480 18816 57486 18828
rect 62209 18819 62267 18825
rect 62209 18816 62221 18819
rect 57480 18788 62221 18816
rect 57480 18776 57486 18788
rect 62209 18785 62221 18788
rect 62255 18785 62267 18819
rect 62209 18779 62267 18785
rect 64969 18819 65027 18825
rect 64969 18785 64981 18819
rect 65015 18816 65027 18819
rect 65334 18816 65340 18828
rect 65015 18788 65340 18816
rect 65015 18785 65027 18788
rect 64969 18779 65027 18785
rect 65334 18776 65340 18788
rect 65392 18776 65398 18828
rect 96982 18816 96988 18828
rect 96943 18788 96988 18816
rect 96982 18776 96988 18788
rect 97040 18776 97046 18828
rect 97169 18819 97227 18825
rect 97169 18785 97181 18819
rect 97215 18785 97227 18819
rect 97169 18779 97227 18785
rect 42794 18708 42800 18760
rect 42852 18748 42858 18760
rect 47394 18748 47400 18760
rect 42852 18720 47400 18748
rect 42852 18708 42858 18720
rect 47394 18708 47400 18720
rect 47452 18708 47458 18760
rect 55030 18708 55036 18760
rect 55088 18748 55094 18760
rect 61930 18748 61936 18760
rect 55088 18720 61936 18748
rect 55088 18708 55094 18720
rect 61930 18708 61936 18720
rect 61988 18748 61994 18760
rect 62666 18748 62672 18760
rect 61988 18720 62672 18748
rect 61988 18708 61994 18720
rect 62666 18708 62672 18720
rect 62724 18708 62730 18760
rect 96709 18751 96767 18757
rect 96709 18717 96721 18751
rect 96755 18748 96767 18751
rect 97184 18748 97212 18779
rect 97258 18776 97264 18828
rect 97316 18816 97322 18828
rect 97552 18825 97580 18856
rect 97537 18819 97595 18825
rect 97316 18788 97361 18816
rect 97316 18776 97322 18788
rect 97537 18785 97549 18819
rect 97583 18785 97595 18819
rect 97537 18779 97595 18785
rect 96755 18720 97212 18748
rect 97353 18751 97411 18757
rect 96755 18717 96767 18720
rect 96709 18711 96767 18717
rect 97353 18717 97365 18751
rect 97399 18748 97411 18751
rect 97644 18748 97672 18924
rect 97399 18720 97672 18748
rect 97399 18717 97411 18720
rect 97353 18711 97411 18717
rect 12250 18640 12256 18692
rect 12308 18680 12314 18692
rect 20714 18680 20720 18692
rect 12308 18652 20720 18680
rect 12308 18640 12314 18652
rect 20714 18640 20720 18652
rect 20772 18640 20778 18692
rect 34514 18640 34520 18692
rect 34572 18680 34578 18692
rect 35802 18680 35808 18692
rect 34572 18652 35808 18680
rect 34572 18640 34578 18652
rect 35802 18640 35808 18652
rect 35860 18680 35866 18692
rect 38102 18680 38108 18692
rect 35860 18652 38108 18680
rect 35860 18640 35866 18652
rect 38102 18640 38108 18652
rect 38160 18640 38166 18692
rect 50614 18680 50620 18692
rect 48332 18652 50620 18680
rect 46842 18572 46848 18624
rect 46900 18612 46906 18624
rect 48332 18612 48360 18652
rect 50614 18640 50620 18652
rect 50672 18640 50678 18692
rect 59446 18640 59452 18692
rect 59504 18680 59510 18692
rect 59504 18652 61332 18680
rect 59504 18640 59510 18652
rect 46900 18584 48360 18612
rect 46900 18572 46906 18584
rect 49970 18572 49976 18624
rect 50028 18612 50034 18624
rect 55950 18612 55956 18624
rect 50028 18584 55956 18612
rect 50028 18572 50034 18584
rect 55950 18572 55956 18584
rect 56008 18572 56014 18624
rect 61304 18612 61332 18652
rect 77938 18640 77944 18692
rect 77996 18680 78002 18692
rect 97721 18683 97779 18689
rect 97721 18680 97733 18683
rect 77996 18652 97733 18680
rect 77996 18640 78002 18652
rect 97721 18649 97733 18652
rect 97767 18649 97779 18683
rect 97721 18643 97779 18649
rect 96709 18615 96767 18621
rect 96709 18612 96721 18615
rect 61304 18584 96721 18612
rect 96709 18581 96721 18584
rect 96755 18612 96767 18615
rect 96801 18615 96859 18621
rect 96801 18612 96813 18615
rect 96755 18584 96813 18612
rect 96755 18581 96767 18584
rect 96709 18575 96767 18581
rect 96801 18581 96813 18584
rect 96847 18581 96859 18615
rect 96801 18575 96859 18581
rect 1104 18522 98808 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 65686 18522
rect 65738 18470 65750 18522
rect 65802 18470 65814 18522
rect 65866 18470 65878 18522
rect 65930 18470 96406 18522
rect 96458 18470 96470 18522
rect 96522 18470 96534 18522
rect 96586 18470 96598 18522
rect 96650 18470 98808 18522
rect 1104 18448 98808 18470
rect 56597 18411 56655 18417
rect 56597 18377 56609 18411
rect 56643 18408 56655 18411
rect 62114 18408 62120 18420
rect 56643 18380 62120 18408
rect 56643 18377 56655 18380
rect 56597 18371 56655 18377
rect 62114 18368 62120 18380
rect 62172 18368 62178 18420
rect 73338 18408 73344 18420
rect 64846 18380 73200 18408
rect 73299 18380 73344 18408
rect 58250 18300 58256 18352
rect 58308 18340 58314 18352
rect 64846 18340 64874 18380
rect 58308 18312 64874 18340
rect 58308 18300 58314 18312
rect 67634 18300 67640 18352
rect 67692 18340 67698 18352
rect 71130 18340 71136 18352
rect 67692 18312 70903 18340
rect 67692 18300 67698 18312
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 19484 18244 19533 18272
rect 19484 18232 19490 18244
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 19886 18232 19892 18284
rect 19944 18272 19950 18284
rect 28350 18272 28356 18284
rect 19944 18244 28356 18272
rect 19944 18232 19950 18244
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 29917 18275 29975 18281
rect 29917 18241 29929 18275
rect 29963 18272 29975 18275
rect 34514 18272 34520 18284
rect 29963 18244 34520 18272
rect 29963 18241 29975 18244
rect 29917 18235 29975 18241
rect 34514 18232 34520 18244
rect 34572 18232 34578 18284
rect 41386 18244 55904 18272
rect 19334 18204 19340 18216
rect 19295 18176 19340 18204
rect 19334 18164 19340 18176
rect 19392 18164 19398 18216
rect 30190 18204 30196 18216
rect 30151 18176 30196 18204
rect 30190 18164 30196 18176
rect 30248 18164 30254 18216
rect 31573 18207 31631 18213
rect 31573 18173 31585 18207
rect 31619 18204 31631 18207
rect 31662 18204 31668 18216
rect 31619 18176 31668 18204
rect 31619 18173 31631 18176
rect 31573 18167 31631 18173
rect 31662 18164 31668 18176
rect 31720 18164 31726 18216
rect 41386 18204 41414 18244
rect 55030 18204 55036 18216
rect 35866 18176 41414 18204
rect 54991 18176 55036 18204
rect 18598 18096 18604 18148
rect 18656 18136 18662 18148
rect 18656 18108 22094 18136
rect 18656 18096 18662 18108
rect 22066 18068 22094 18108
rect 30852 18108 31754 18136
rect 30852 18068 30880 18108
rect 22066 18040 30880 18068
rect 31726 18068 31754 18108
rect 35866 18068 35894 18176
rect 55030 18164 55036 18176
rect 55088 18164 55094 18216
rect 55306 18204 55312 18216
rect 55267 18176 55312 18204
rect 55306 18164 55312 18176
rect 55364 18164 55370 18216
rect 55876 18204 55904 18244
rect 55950 18232 55956 18284
rect 56008 18272 56014 18284
rect 67726 18272 67732 18284
rect 56008 18244 67732 18272
rect 56008 18232 56014 18244
rect 67726 18232 67732 18244
rect 67784 18232 67790 18284
rect 70875 18281 70903 18312
rect 70964 18312 71136 18340
rect 70964 18281 70992 18312
rect 71130 18300 71136 18312
rect 71188 18300 71194 18352
rect 71314 18340 71320 18352
rect 71275 18312 71320 18340
rect 71314 18300 71320 18312
rect 71372 18300 71378 18352
rect 70857 18275 70915 18281
rect 70412 18244 70780 18272
rect 70412 18213 70440 18244
rect 70397 18207 70455 18213
rect 70397 18204 70409 18207
rect 55876 18176 70409 18204
rect 70397 18173 70409 18176
rect 70443 18173 70455 18207
rect 70578 18204 70584 18216
rect 70539 18176 70584 18204
rect 70397 18167 70455 18173
rect 70578 18164 70584 18176
rect 70636 18164 70642 18216
rect 70752 18213 70780 18244
rect 70857 18241 70869 18275
rect 70903 18241 70915 18275
rect 70857 18235 70915 18241
rect 70949 18275 71007 18281
rect 70949 18241 70961 18275
rect 70995 18241 71007 18275
rect 70949 18235 71007 18241
rect 70752 18207 70811 18213
rect 70752 18176 70765 18207
rect 70753 18173 70765 18176
rect 70799 18173 70811 18207
rect 70753 18167 70811 18173
rect 71133 18207 71191 18213
rect 71133 18173 71145 18207
rect 71179 18204 71191 18207
rect 71682 18204 71688 18216
rect 71179 18176 71688 18204
rect 71179 18173 71191 18176
rect 71133 18167 71191 18173
rect 71682 18164 71688 18176
rect 71740 18164 71746 18216
rect 73172 18213 73200 18380
rect 73338 18368 73344 18380
rect 73396 18368 73402 18420
rect 73157 18207 73215 18213
rect 73157 18173 73169 18207
rect 73203 18173 73215 18207
rect 73157 18167 73215 18173
rect 59722 18096 59728 18148
rect 59780 18136 59786 18148
rect 70486 18136 70492 18148
rect 59780 18108 70492 18136
rect 59780 18096 59786 18108
rect 70486 18096 70492 18108
rect 70544 18096 70550 18148
rect 71314 18096 71320 18148
rect 71372 18136 71378 18148
rect 96706 18136 96712 18148
rect 71372 18108 96712 18136
rect 71372 18096 71378 18108
rect 96706 18096 96712 18108
rect 96764 18136 96770 18148
rect 96982 18136 96988 18148
rect 96764 18108 96988 18136
rect 96764 18096 96770 18108
rect 96982 18096 96988 18108
rect 97040 18096 97046 18148
rect 31726 18040 35894 18068
rect 38102 18028 38108 18080
rect 38160 18068 38166 18080
rect 42794 18068 42800 18080
rect 38160 18040 42800 18068
rect 38160 18028 38166 18040
rect 42794 18028 42800 18040
rect 42852 18028 42858 18080
rect 51258 18028 51264 18080
rect 51316 18068 51322 18080
rect 53282 18068 53288 18080
rect 51316 18040 53288 18068
rect 51316 18028 51322 18040
rect 53282 18028 53288 18040
rect 53340 18028 53346 18080
rect 1104 17978 98808 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 50326 17978
rect 50378 17926 50390 17978
rect 50442 17926 50454 17978
rect 50506 17926 50518 17978
rect 50570 17926 81046 17978
rect 81098 17926 81110 17978
rect 81162 17926 81174 17978
rect 81226 17926 81238 17978
rect 81290 17926 98808 17978
rect 1104 17904 98808 17926
rect 60274 17824 60280 17876
rect 60332 17864 60338 17876
rect 61102 17864 61108 17876
rect 60332 17836 61108 17864
rect 60332 17824 60338 17836
rect 61102 17824 61108 17836
rect 61160 17824 61166 17876
rect 66990 17824 66996 17876
rect 67048 17864 67054 17876
rect 69842 17864 69848 17876
rect 67048 17836 69848 17864
rect 67048 17824 67054 17836
rect 69842 17824 69848 17836
rect 69900 17824 69906 17876
rect 34054 17620 34060 17672
rect 34112 17660 34118 17672
rect 39850 17660 39856 17672
rect 34112 17632 39856 17660
rect 34112 17620 34118 17632
rect 39850 17620 39856 17632
rect 39908 17620 39914 17672
rect 44450 17620 44456 17672
rect 44508 17660 44514 17672
rect 48314 17660 48320 17672
rect 44508 17632 48320 17660
rect 44508 17620 44514 17632
rect 48314 17620 48320 17632
rect 48372 17660 48378 17672
rect 73706 17660 73712 17672
rect 48372 17632 73712 17660
rect 48372 17620 48378 17632
rect 73706 17620 73712 17632
rect 73764 17620 73770 17672
rect 24762 17552 24768 17604
rect 24820 17592 24826 17604
rect 77662 17592 77668 17604
rect 24820 17564 77668 17592
rect 24820 17552 24826 17564
rect 77662 17552 77668 17564
rect 77720 17552 77726 17604
rect 17126 17524 17132 17536
rect 17087 17496 17132 17524
rect 17126 17484 17132 17496
rect 17184 17484 17190 17536
rect 20441 17527 20499 17533
rect 20441 17493 20453 17527
rect 20487 17524 20499 17527
rect 25958 17524 25964 17536
rect 20487 17496 25964 17524
rect 20487 17493 20499 17496
rect 20441 17487 20499 17493
rect 25958 17484 25964 17496
rect 26016 17484 26022 17536
rect 31110 17484 31116 17536
rect 31168 17524 31174 17536
rect 32585 17527 32643 17533
rect 32585 17524 32597 17527
rect 31168 17496 32597 17524
rect 31168 17484 31174 17496
rect 32585 17493 32597 17496
rect 32631 17493 32643 17527
rect 32585 17487 32643 17493
rect 34238 17484 34244 17536
rect 34296 17524 34302 17536
rect 43806 17524 43812 17536
rect 34296 17496 43812 17524
rect 34296 17484 34302 17496
rect 43806 17484 43812 17496
rect 43864 17484 43870 17536
rect 62117 17527 62175 17533
rect 62117 17493 62129 17527
rect 62163 17524 62175 17527
rect 62390 17524 62396 17536
rect 62163 17496 62396 17524
rect 62163 17493 62175 17496
rect 62117 17487 62175 17493
rect 62390 17484 62396 17496
rect 62448 17484 62454 17536
rect 1104 17434 98808 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 65686 17434
rect 65738 17382 65750 17434
rect 65802 17382 65814 17434
rect 65866 17382 65878 17434
rect 65930 17382 96406 17434
rect 96458 17382 96470 17434
rect 96522 17382 96534 17434
rect 96586 17382 96598 17434
rect 96650 17382 98808 17434
rect 1104 17360 98808 17382
rect 26326 17280 26332 17332
rect 26384 17320 26390 17332
rect 72602 17320 72608 17332
rect 26384 17292 72608 17320
rect 26384 17280 26390 17292
rect 72602 17280 72608 17292
rect 72660 17280 72666 17332
rect 81526 17280 81532 17332
rect 81584 17320 81590 17332
rect 81584 17292 87184 17320
rect 81584 17280 81590 17292
rect 4982 17212 4988 17264
rect 5040 17252 5046 17264
rect 71222 17252 71228 17264
rect 5040 17224 71228 17252
rect 5040 17212 5046 17224
rect 71222 17212 71228 17224
rect 71280 17212 71286 17264
rect 72418 17212 72424 17264
rect 72476 17252 72482 17264
rect 79870 17252 79876 17264
rect 72476 17224 79876 17252
rect 72476 17212 72482 17224
rect 79870 17212 79876 17224
rect 79928 17212 79934 17264
rect 80146 17212 80152 17264
rect 80204 17252 80210 17264
rect 80204 17224 87092 17252
rect 80204 17212 80210 17224
rect 17126 17144 17132 17196
rect 17184 17184 17190 17196
rect 33686 17184 33692 17196
rect 17184 17156 33692 17184
rect 17184 17144 17190 17156
rect 33686 17144 33692 17156
rect 33744 17144 33750 17196
rect 44634 17144 44640 17196
rect 44692 17184 44698 17196
rect 66990 17184 66996 17196
rect 44692 17156 66996 17184
rect 44692 17144 44698 17156
rect 66990 17144 66996 17156
rect 67048 17144 67054 17196
rect 72510 17144 72516 17196
rect 72568 17184 72574 17196
rect 81526 17184 81532 17196
rect 72568 17156 81532 17184
rect 72568 17144 72574 17156
rect 81526 17144 81532 17156
rect 81584 17144 81590 17196
rect 87064 17193 87092 17224
rect 87156 17193 87184 17292
rect 87049 17187 87107 17193
rect 87049 17153 87061 17187
rect 87095 17153 87107 17187
rect 87049 17147 87107 17153
rect 87141 17187 87199 17193
rect 87141 17153 87153 17187
rect 87187 17153 87199 17187
rect 87141 17147 87199 17153
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17116 14979 17119
rect 44545 17119 44603 17125
rect 14967 17088 22094 17116
rect 14967 17085 14979 17088
rect 14921 17079 14979 17085
rect 22066 17048 22094 17088
rect 44545 17085 44557 17119
rect 44591 17116 44603 17119
rect 46474 17116 46480 17128
rect 44591 17088 46480 17116
rect 44591 17085 44603 17088
rect 44545 17079 44603 17085
rect 46474 17076 46480 17088
rect 46532 17076 46538 17128
rect 86681 17119 86739 17125
rect 86681 17116 86693 17119
rect 64846 17088 86693 17116
rect 49050 17048 49056 17060
rect 22066 17020 49056 17048
rect 49050 17008 49056 17020
rect 49108 17008 49114 17060
rect 55306 17008 55312 17060
rect 55364 17048 55370 17060
rect 64846 17048 64874 17088
rect 86681 17085 86693 17088
rect 86727 17085 86739 17119
rect 86862 17116 86868 17128
rect 86823 17088 86868 17116
rect 86681 17079 86739 17085
rect 86862 17076 86868 17088
rect 86920 17076 86926 17128
rect 87234 17119 87292 17125
rect 87234 17116 87246 17119
rect 87156 17088 87246 17116
rect 87156 17048 87184 17088
rect 87234 17085 87246 17088
rect 87280 17085 87292 17119
rect 87414 17116 87420 17128
rect 87375 17088 87420 17116
rect 87234 17079 87292 17085
rect 87414 17076 87420 17088
rect 87472 17076 87478 17128
rect 97166 17116 97172 17128
rect 97127 17088 97172 17116
rect 97166 17076 97172 17088
rect 97224 17076 97230 17128
rect 55364 17020 64874 17048
rect 86512 17020 87184 17048
rect 55364 17008 55370 17020
rect 21174 16940 21180 16992
rect 21232 16980 21238 16992
rect 21358 16980 21364 16992
rect 21232 16952 21364 16980
rect 21232 16940 21238 16952
rect 21358 16940 21364 16952
rect 21416 16980 21422 16992
rect 86512 16989 86540 17020
rect 86497 16983 86555 16989
rect 86497 16980 86509 16983
rect 21416 16952 86509 16980
rect 21416 16940 21422 16952
rect 86497 16949 86509 16952
rect 86543 16949 86555 16983
rect 86497 16943 86555 16949
rect 1104 16890 98808 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 50326 16890
rect 50378 16838 50390 16890
rect 50442 16838 50454 16890
rect 50506 16838 50518 16890
rect 50570 16838 81046 16890
rect 81098 16838 81110 16890
rect 81162 16838 81174 16890
rect 81226 16838 81238 16890
rect 81290 16838 98808 16890
rect 1104 16816 98808 16838
rect 44726 16776 44732 16788
rect 8220 16748 12434 16776
rect 44687 16748 44732 16776
rect 6270 16668 6276 16720
rect 6328 16708 6334 16720
rect 8021 16711 8079 16717
rect 8021 16708 8033 16711
rect 6328 16680 8033 16708
rect 6328 16668 6334 16680
rect 8021 16677 8033 16680
rect 8067 16677 8079 16711
rect 8021 16671 8079 16677
rect 8220 16649 8248 16748
rect 8481 16711 8539 16717
rect 8481 16677 8493 16711
rect 8527 16708 8539 16711
rect 8570 16708 8576 16720
rect 8527 16680 8576 16708
rect 8527 16677 8539 16680
rect 8481 16671 8539 16677
rect 8570 16668 8576 16680
rect 8628 16668 8634 16720
rect 12406 16708 12434 16748
rect 44726 16736 44732 16748
rect 44784 16736 44790 16788
rect 47670 16776 47676 16788
rect 47631 16748 47676 16776
rect 47670 16736 47676 16748
rect 47728 16736 47734 16788
rect 48038 16776 48044 16788
rect 47872 16748 48044 16776
rect 24302 16708 24308 16720
rect 12406 16680 24308 16708
rect 24302 16668 24308 16680
rect 24360 16708 24366 16720
rect 24762 16708 24768 16720
rect 24360 16680 24768 16708
rect 24360 16668 24366 16680
rect 24762 16668 24768 16680
rect 24820 16668 24826 16720
rect 44450 16708 44456 16720
rect 31726 16680 44456 16708
rect 7837 16643 7895 16649
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8205 16643 8263 16649
rect 8205 16640 8217 16643
rect 7883 16612 8217 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8205 16609 8217 16612
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16640 8447 16643
rect 8938 16640 8944 16652
rect 8435 16612 8944 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 8938 16600 8944 16612
rect 8996 16600 9002 16652
rect 20254 16600 20260 16652
rect 20312 16640 20318 16652
rect 31726 16640 31754 16680
rect 44450 16668 44456 16680
rect 44508 16668 44514 16720
rect 44634 16708 44640 16720
rect 44595 16680 44640 16708
rect 44634 16668 44640 16680
rect 44692 16668 44698 16720
rect 20312 16612 31754 16640
rect 47872 16640 47900 16748
rect 48038 16736 48044 16748
rect 48096 16736 48102 16788
rect 48314 16736 48320 16788
rect 48372 16736 48378 16788
rect 58618 16776 58624 16788
rect 48700 16748 58624 16776
rect 48332 16649 48360 16736
rect 48498 16649 48504 16652
rect 48029 16643 48087 16649
rect 48029 16640 48041 16643
rect 47872 16612 48041 16640
rect 20312 16600 20318 16612
rect 48029 16609 48041 16612
rect 48075 16609 48087 16643
rect 48029 16603 48087 16609
rect 48317 16643 48375 16649
rect 48317 16609 48329 16643
rect 48363 16609 48375 16643
rect 48317 16603 48375 16609
rect 48455 16643 48504 16649
rect 48455 16609 48467 16643
rect 48501 16609 48504 16643
rect 48455 16603 48504 16609
rect 48498 16600 48504 16603
rect 48556 16600 48562 16652
rect 48700 16649 48728 16748
rect 58618 16736 58624 16748
rect 58676 16736 58682 16788
rect 68370 16736 68376 16788
rect 68428 16776 68434 16788
rect 97166 16776 97172 16788
rect 68428 16748 97172 16776
rect 68428 16736 68434 16748
rect 97166 16736 97172 16748
rect 97224 16736 97230 16788
rect 48685 16643 48743 16649
rect 48685 16609 48697 16643
rect 48731 16609 48743 16643
rect 48685 16603 48743 16609
rect 48961 16643 49019 16649
rect 48961 16609 48973 16643
rect 49007 16640 49019 16643
rect 49694 16640 49700 16652
rect 49007 16612 49700 16640
rect 49007 16609 49019 16612
rect 48961 16603 49019 16609
rect 49694 16600 49700 16612
rect 49752 16640 49758 16652
rect 50154 16640 50160 16652
rect 49752 16612 50160 16640
rect 49752 16600 49758 16612
rect 50154 16600 50160 16612
rect 50212 16600 50218 16652
rect 14550 16532 14556 16584
rect 14608 16572 14614 16584
rect 79410 16572 79416 16584
rect 14608 16544 38654 16572
rect 14608 16532 14614 16544
rect 38626 16504 38654 16544
rect 48286 16544 79416 16572
rect 48286 16504 48314 16544
rect 79410 16532 79416 16544
rect 79468 16532 79474 16584
rect 38626 16476 48314 16504
rect 46198 16396 46204 16448
rect 46256 16436 46262 16448
rect 67542 16436 67548 16448
rect 46256 16408 67548 16436
rect 46256 16396 46262 16408
rect 67542 16396 67548 16408
rect 67600 16396 67606 16448
rect 1104 16346 98808 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 65686 16346
rect 65738 16294 65750 16346
rect 65802 16294 65814 16346
rect 65866 16294 65878 16346
rect 65930 16294 96406 16346
rect 96458 16294 96470 16346
rect 96522 16294 96534 16346
rect 96586 16294 96598 16346
rect 96650 16294 98808 16346
rect 1104 16272 98808 16294
rect 25958 16192 25964 16244
rect 26016 16232 26022 16244
rect 42426 16232 42432 16244
rect 26016 16204 42432 16232
rect 26016 16192 26022 16204
rect 42426 16192 42432 16204
rect 42484 16192 42490 16244
rect 59262 16192 59268 16244
rect 59320 16232 59326 16244
rect 95970 16232 95976 16244
rect 59320 16204 95976 16232
rect 59320 16192 59326 16204
rect 95970 16192 95976 16204
rect 96028 16192 96034 16244
rect 37826 16124 37832 16176
rect 37884 16164 37890 16176
rect 85942 16164 85948 16176
rect 37884 16136 85948 16164
rect 37884 16124 37890 16136
rect 85942 16124 85948 16136
rect 86000 16124 86006 16176
rect 9858 16056 9864 16108
rect 9916 16096 9922 16108
rect 28994 16096 29000 16108
rect 9916 16068 29000 16096
rect 9916 16056 9922 16068
rect 28994 16056 29000 16068
rect 29052 16056 29058 16108
rect 40034 16056 40040 16108
rect 40092 16096 40098 16108
rect 89070 16096 89076 16108
rect 40092 16068 89076 16096
rect 40092 16056 40098 16068
rect 89070 16056 89076 16068
rect 89128 16056 89134 16108
rect 19242 15988 19248 16040
rect 19300 16028 19306 16040
rect 71406 16028 71412 16040
rect 19300 16000 71412 16028
rect 19300 15988 19306 16000
rect 71406 15988 71412 16000
rect 71464 15988 71470 16040
rect 2498 15920 2504 15972
rect 2556 15960 2562 15972
rect 13630 15960 13636 15972
rect 2556 15932 13636 15960
rect 2556 15920 2562 15932
rect 13630 15920 13636 15932
rect 13688 15920 13694 15972
rect 17770 15920 17776 15972
rect 17828 15960 17834 15972
rect 80330 15960 80336 15972
rect 17828 15932 80336 15960
rect 17828 15920 17834 15932
rect 80330 15920 80336 15932
rect 80388 15920 80394 15972
rect 2406 15852 2412 15904
rect 2464 15892 2470 15904
rect 69750 15892 69756 15904
rect 2464 15864 69756 15892
rect 2464 15852 2470 15864
rect 69750 15852 69756 15864
rect 69808 15852 69814 15904
rect 79410 15852 79416 15904
rect 79468 15892 79474 15904
rect 93854 15892 93860 15904
rect 79468 15864 93860 15892
rect 79468 15852 79474 15864
rect 93854 15852 93860 15864
rect 93912 15852 93918 15904
rect 1104 15802 98808 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 50326 15802
rect 50378 15750 50390 15802
rect 50442 15750 50454 15802
rect 50506 15750 50518 15802
rect 50570 15750 81046 15802
rect 81098 15750 81110 15802
rect 81162 15750 81174 15802
rect 81226 15750 81238 15802
rect 81290 15750 98808 15802
rect 1104 15728 98808 15750
rect 58066 15688 58072 15700
rect 58027 15660 58072 15688
rect 58066 15648 58072 15660
rect 58124 15648 58130 15700
rect 57974 15620 57980 15632
rect 57935 15592 57980 15620
rect 57974 15580 57980 15592
rect 58032 15580 58038 15632
rect 13630 15376 13636 15428
rect 13688 15416 13694 15428
rect 31662 15416 31668 15428
rect 13688 15388 31668 15416
rect 13688 15376 13694 15388
rect 31662 15376 31668 15388
rect 31720 15376 31726 15428
rect 21913 15351 21971 15357
rect 21913 15317 21925 15351
rect 21959 15348 21971 15351
rect 22189 15351 22247 15357
rect 22189 15348 22201 15351
rect 21959 15320 22201 15348
rect 21959 15317 21971 15320
rect 21913 15311 21971 15317
rect 22189 15317 22201 15320
rect 22235 15348 22247 15351
rect 92290 15348 92296 15360
rect 22235 15320 92296 15348
rect 22235 15317 22247 15320
rect 22189 15311 22247 15317
rect 92290 15308 92296 15320
rect 92348 15308 92354 15360
rect 1104 15258 98808 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 65686 15258
rect 65738 15206 65750 15258
rect 65802 15206 65814 15258
rect 65866 15206 65878 15258
rect 65930 15206 96406 15258
rect 96458 15206 96470 15258
rect 96522 15206 96534 15258
rect 96586 15206 96598 15258
rect 96650 15206 98808 15258
rect 1104 15184 98808 15206
rect 13998 15104 14004 15156
rect 14056 15144 14062 15156
rect 14550 15144 14556 15156
rect 14056 15116 14556 15144
rect 14056 15104 14062 15116
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 15562 15104 15568 15156
rect 15620 15144 15626 15156
rect 15620 15116 22094 15144
rect 15620 15104 15626 15116
rect 18690 15076 18696 15088
rect 13372 15048 18696 15076
rect 13372 14949 13400 15048
rect 18690 15036 18696 15048
rect 18748 15036 18754 15088
rect 22066 15076 22094 15116
rect 55766 15104 55772 15156
rect 55824 15144 55830 15156
rect 84378 15144 84384 15156
rect 55824 15116 84384 15144
rect 55824 15104 55830 15116
rect 84378 15104 84384 15116
rect 84436 15104 84442 15156
rect 59446 15076 59452 15088
rect 22066 15048 59452 15076
rect 59446 15036 59452 15048
rect 59504 15036 59510 15088
rect 61838 15036 61844 15088
rect 61896 15076 61902 15088
rect 97810 15076 97816 15088
rect 61896 15048 97816 15076
rect 61896 15036 61902 15048
rect 97810 15036 97816 15048
rect 97868 15036 97874 15088
rect 15930 15008 15936 15020
rect 13740 14980 15936 15008
rect 13357 14943 13415 14949
rect 13357 14909 13369 14943
rect 13403 14909 13415 14943
rect 13630 14940 13636 14952
rect 13591 14912 13636 14940
rect 13357 14903 13415 14909
rect 13630 14900 13636 14912
rect 13688 14900 13694 14952
rect 13740 14949 13768 14980
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 15008 16727 15011
rect 63402 15008 63408 15020
rect 16715 14980 63408 15008
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 63402 14968 63408 14980
rect 63460 14968 63466 15020
rect 71777 15011 71835 15017
rect 71777 14977 71789 15011
rect 71823 15008 71835 15011
rect 72053 15011 72111 15017
rect 72053 15008 72065 15011
rect 71823 14980 72065 15008
rect 71823 14977 71835 14980
rect 71777 14971 71835 14977
rect 72053 14977 72065 14980
rect 72099 15008 72111 15011
rect 72099 14980 80054 15008
rect 72099 14977 72111 14980
rect 72053 14971 72111 14977
rect 13725 14943 13783 14949
rect 13725 14909 13737 14943
rect 13771 14909 13783 14943
rect 13998 14940 14004 14952
rect 13959 14912 14004 14940
rect 13725 14903 13783 14909
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 14277 14943 14335 14949
rect 14277 14909 14289 14943
rect 14323 14940 14335 14943
rect 35250 14940 35256 14952
rect 14323 14912 35256 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 35250 14900 35256 14912
rect 35308 14900 35314 14952
rect 44818 14900 44824 14952
rect 44876 14940 44882 14952
rect 54757 14943 54815 14949
rect 54757 14940 54769 14943
rect 44876 14912 54769 14940
rect 44876 14900 44882 14912
rect 54757 14909 54769 14912
rect 54803 14909 54815 14943
rect 71593 14943 71651 14949
rect 71593 14940 71605 14943
rect 54757 14903 54815 14909
rect 70366 14912 71605 14940
rect 13814 14832 13820 14884
rect 13872 14872 13878 14884
rect 16669 14875 16727 14881
rect 16669 14872 16681 14875
rect 13872 14844 16681 14872
rect 13872 14832 13878 14844
rect 16669 14841 16681 14844
rect 16715 14841 16727 14875
rect 16669 14835 16727 14841
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 33962 14872 33968 14884
rect 17276 14844 33968 14872
rect 17276 14832 17282 14844
rect 33962 14832 33968 14844
rect 34020 14832 34026 14884
rect 54021 14875 54079 14881
rect 54021 14841 54033 14875
rect 54067 14872 54079 14875
rect 55214 14872 55220 14884
rect 54067 14844 55220 14872
rect 54067 14841 54079 14844
rect 54021 14835 54079 14841
rect 55214 14832 55220 14844
rect 55272 14832 55278 14884
rect 70366 14872 70394 14912
rect 71593 14909 71605 14912
rect 71639 14909 71651 14943
rect 80026 14940 80054 14980
rect 97902 14940 97908 14952
rect 80026 14912 97908 14940
rect 71593 14903 71651 14909
rect 97902 14900 97908 14912
rect 97960 14900 97966 14952
rect 96062 14872 96068 14884
rect 64846 14844 70394 14872
rect 71516 14844 96068 14872
rect 12989 14807 13047 14813
rect 12989 14773 13001 14807
rect 13035 14804 13047 14807
rect 64846 14804 64874 14844
rect 13035 14776 64874 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 66806 14764 66812 14816
rect 66864 14804 66870 14816
rect 71516 14804 71544 14844
rect 96062 14832 96068 14844
rect 96120 14832 96126 14884
rect 66864 14776 71544 14804
rect 71593 14807 71651 14813
rect 66864 14764 66870 14776
rect 71593 14773 71605 14807
rect 71639 14804 71651 14807
rect 87782 14804 87788 14816
rect 71639 14776 87788 14804
rect 71639 14773 71651 14776
rect 71593 14767 71651 14773
rect 87782 14764 87788 14776
rect 87840 14764 87846 14816
rect 1104 14714 98808 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 50326 14714
rect 50378 14662 50390 14714
rect 50442 14662 50454 14714
rect 50506 14662 50518 14714
rect 50570 14662 81046 14714
rect 81098 14662 81110 14714
rect 81162 14662 81174 14714
rect 81226 14662 81238 14714
rect 81290 14662 98808 14714
rect 1104 14640 98808 14662
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 81618 14600 81624 14612
rect 18564 14572 81624 14600
rect 18564 14560 18570 14572
rect 81618 14560 81624 14572
rect 81676 14560 81682 14612
rect 23014 14492 23020 14544
rect 23072 14532 23078 14544
rect 92106 14532 92112 14544
rect 23072 14504 92112 14532
rect 23072 14492 23078 14504
rect 92106 14492 92112 14504
rect 92164 14492 92170 14544
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 42978 14464 42984 14476
rect 13596 14436 42984 14464
rect 13596 14424 13602 14436
rect 42978 14424 42984 14436
rect 43036 14424 43042 14476
rect 44358 14464 44364 14476
rect 44319 14436 44364 14464
rect 44358 14424 44364 14436
rect 44416 14424 44422 14476
rect 44544 14467 44602 14473
rect 44544 14433 44556 14467
rect 44590 14433 44602 14467
rect 44726 14464 44732 14476
rect 44687 14436 44732 14464
rect 44544 14427 44602 14433
rect 44559 14340 44587 14427
rect 44726 14424 44732 14436
rect 44784 14424 44790 14476
rect 44818 14424 44824 14476
rect 44876 14473 44882 14476
rect 44876 14467 44925 14473
rect 44876 14433 44879 14467
rect 44913 14433 44925 14467
rect 44876 14427 44925 14433
rect 44876 14424 44882 14427
rect 45002 14424 45008 14476
rect 45060 14464 45066 14476
rect 74994 14464 75000 14476
rect 45060 14436 75000 14464
rect 45060 14424 45066 14436
rect 74994 14424 75000 14436
rect 75052 14424 75058 14476
rect 82906 14464 82912 14476
rect 82867 14436 82912 14464
rect 82906 14424 82912 14436
rect 82964 14424 82970 14476
rect 44637 14399 44695 14405
rect 44637 14365 44649 14399
rect 44683 14365 44695 14399
rect 45281 14399 45339 14405
rect 45281 14396 45293 14399
rect 44637 14359 44695 14365
rect 45020 14368 45293 14396
rect 22094 14288 22100 14340
rect 22152 14328 22158 14340
rect 44177 14331 44235 14337
rect 44177 14328 44189 14331
rect 22152 14300 44189 14328
rect 22152 14288 22158 14300
rect 44177 14297 44189 14300
rect 44223 14328 44235 14331
rect 44542 14328 44548 14340
rect 44223 14300 44548 14328
rect 44223 14297 44235 14300
rect 44177 14291 44235 14297
rect 44542 14288 44548 14300
rect 44600 14288 44606 14340
rect 44652 14328 44680 14359
rect 45020 14328 45048 14368
rect 45281 14365 45293 14368
rect 45327 14396 45339 14399
rect 77018 14396 77024 14408
rect 45327 14368 77024 14396
rect 45327 14365 45339 14368
rect 45281 14359 45339 14365
rect 77018 14356 77024 14368
rect 77076 14356 77082 14408
rect 44652 14300 45048 14328
rect 45370 14288 45376 14340
rect 45428 14328 45434 14340
rect 57238 14328 57244 14340
rect 45428 14300 57244 14328
rect 45428 14288 45434 14300
rect 57238 14288 57244 14300
rect 57296 14288 57302 14340
rect 61654 14288 61660 14340
rect 61712 14328 61718 14340
rect 67174 14328 67180 14340
rect 61712 14300 67180 14328
rect 61712 14288 61718 14300
rect 67174 14288 67180 14300
rect 67232 14288 67238 14340
rect 37734 14260 37740 14272
rect 37695 14232 37740 14260
rect 37734 14220 37740 14232
rect 37792 14220 37798 14272
rect 45005 14263 45063 14269
rect 45005 14229 45017 14263
rect 45051 14260 45063 14263
rect 46658 14260 46664 14272
rect 45051 14232 46664 14260
rect 45051 14229 45063 14232
rect 45005 14223 45063 14229
rect 46658 14220 46664 14232
rect 46716 14220 46722 14272
rect 49694 14220 49700 14272
rect 49752 14260 49758 14272
rect 54478 14260 54484 14272
rect 49752 14232 54484 14260
rect 49752 14220 49758 14232
rect 54478 14220 54484 14232
rect 54536 14220 54542 14272
rect 55214 14220 55220 14272
rect 55272 14260 55278 14272
rect 83093 14263 83151 14269
rect 83093 14260 83105 14263
rect 55272 14232 83105 14260
rect 55272 14220 55278 14232
rect 83093 14229 83105 14232
rect 83139 14229 83151 14263
rect 83093 14223 83151 14229
rect 1104 14170 98808 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 65686 14170
rect 65738 14118 65750 14170
rect 65802 14118 65814 14170
rect 65866 14118 65878 14170
rect 65930 14118 96406 14170
rect 96458 14118 96470 14170
rect 96522 14118 96534 14170
rect 96586 14118 96598 14170
rect 96650 14118 98808 14170
rect 1104 14096 98808 14118
rect 37734 14016 37740 14068
rect 37792 14056 37798 14068
rect 62482 14056 62488 14068
rect 37792 14028 62488 14056
rect 37792 14016 37798 14028
rect 62482 14016 62488 14028
rect 62540 14016 62546 14068
rect 8665 13991 8723 13997
rect 8665 13957 8677 13991
rect 8711 13988 8723 13991
rect 8849 13991 8907 13997
rect 8849 13988 8861 13991
rect 8711 13960 8861 13988
rect 8711 13957 8723 13960
rect 8665 13951 8723 13957
rect 8849 13957 8861 13960
rect 8895 13988 8907 13991
rect 9125 13991 9183 13997
rect 9125 13988 9137 13991
rect 8895 13960 9137 13988
rect 8895 13957 8907 13960
rect 8849 13951 8907 13957
rect 9125 13957 9137 13960
rect 9171 13988 9183 13991
rect 9309 13991 9367 13997
rect 9309 13988 9321 13991
rect 9171 13960 9321 13988
rect 9171 13957 9183 13960
rect 9125 13951 9183 13957
rect 9309 13957 9321 13960
rect 9355 13988 9367 13991
rect 49602 13988 49608 14000
rect 9355 13960 49608 13988
rect 9355 13957 9367 13960
rect 9309 13951 9367 13957
rect 49602 13948 49608 13960
rect 49660 13948 49666 14000
rect 46658 13880 46664 13932
rect 46716 13920 46722 13932
rect 49694 13920 49700 13932
rect 46716 13892 49700 13920
rect 46716 13880 46722 13892
rect 49694 13880 49700 13892
rect 49752 13880 49758 13932
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 16298 13852 16304 13864
rect 12216 13824 16304 13852
rect 12216 13812 12222 13824
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 20165 13855 20223 13861
rect 20165 13821 20177 13855
rect 20211 13852 20223 13855
rect 23198 13852 23204 13864
rect 20211 13824 23204 13852
rect 20211 13821 20223 13824
rect 20165 13815 20223 13821
rect 23198 13812 23204 13824
rect 23256 13812 23262 13864
rect 39758 13852 39764 13864
rect 39719 13824 39764 13852
rect 39758 13812 39764 13824
rect 39816 13812 39822 13864
rect 29362 13744 29368 13796
rect 29420 13784 29426 13796
rect 29730 13784 29736 13796
rect 29420 13756 29736 13784
rect 29420 13744 29426 13756
rect 29730 13744 29736 13756
rect 29788 13744 29794 13796
rect 92198 13744 92204 13796
rect 92256 13784 92262 13796
rect 94038 13784 94044 13796
rect 92256 13756 94044 13784
rect 92256 13744 92262 13756
rect 94038 13744 94044 13756
rect 94096 13744 94102 13796
rect 39945 13719 40003 13725
rect 39945 13685 39957 13719
rect 39991 13716 40003 13719
rect 44726 13716 44732 13728
rect 39991 13688 44732 13716
rect 39991 13685 40003 13688
rect 39945 13679 40003 13685
rect 44726 13676 44732 13688
rect 44784 13676 44790 13728
rect 1104 13626 98808 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 50326 13626
rect 50378 13574 50390 13626
rect 50442 13574 50454 13626
rect 50506 13574 50518 13626
rect 50570 13574 81046 13626
rect 81098 13574 81110 13626
rect 81162 13574 81174 13626
rect 81226 13574 81238 13626
rect 81290 13574 98808 13626
rect 1104 13552 98808 13574
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 36446 13512 36452 13524
rect 11020 13484 36452 13512
rect 11020 13472 11026 13484
rect 36446 13472 36452 13484
rect 36504 13512 36510 13524
rect 37182 13512 37188 13524
rect 36504 13484 37188 13512
rect 36504 13472 36510 13484
rect 37182 13472 37188 13484
rect 37240 13472 37246 13524
rect 11900 13416 12434 13444
rect 11422 13336 11428 13388
rect 11480 13376 11486 13388
rect 11900 13385 11928 13416
rect 11517 13379 11575 13385
rect 11517 13376 11529 13379
rect 11480 13348 11529 13376
rect 11480 13336 11486 13348
rect 11517 13345 11529 13348
rect 11563 13345 11575 13379
rect 11517 13339 11575 13345
rect 11885 13379 11943 13385
rect 11885 13345 11897 13379
rect 11931 13345 11943 13379
rect 12158 13376 12164 13388
rect 12119 13348 12164 13376
rect 11885 13339 11943 13345
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 12253 13379 12311 13385
rect 12253 13345 12265 13379
rect 12299 13345 12311 13379
rect 12406 13376 12434 13416
rect 12526 13404 12532 13456
rect 12584 13444 12590 13456
rect 19978 13444 19984 13456
rect 12584 13416 19984 13444
rect 12584 13404 12590 13416
rect 19978 13404 19984 13416
rect 20036 13404 20042 13456
rect 31018 13376 31024 13388
rect 12406 13348 31024 13376
rect 12253 13339 12311 13345
rect 9306 13268 9312 13320
rect 9364 13308 9370 13320
rect 11701 13311 11759 13317
rect 11701 13308 11713 13311
rect 9364 13280 11713 13308
rect 9364 13268 9370 13280
rect 11701 13277 11713 13280
rect 11747 13277 11759 13311
rect 12268 13308 12296 13339
rect 31018 13336 31024 13348
rect 31076 13336 31082 13388
rect 67358 13376 67364 13388
rect 67319 13348 67364 13376
rect 67358 13336 67364 13348
rect 67416 13336 67422 13388
rect 12526 13308 12532 13320
rect 12268 13280 12532 13308
rect 11701 13271 11759 13277
rect 11716 13172 11744 13271
rect 12526 13268 12532 13280
rect 12584 13268 12590 13320
rect 43254 13308 43260 13320
rect 12636 13280 43260 13308
rect 12636 13172 12664 13280
rect 43254 13268 43260 13280
rect 43312 13268 43318 13320
rect 61562 13268 61568 13320
rect 61620 13308 61626 13320
rect 69750 13308 69756 13320
rect 61620 13280 69756 13308
rect 61620 13268 61626 13280
rect 69750 13268 69756 13280
rect 69808 13268 69814 13320
rect 12713 13243 12771 13249
rect 12713 13209 12725 13243
rect 12759 13240 12771 13243
rect 39574 13240 39580 13252
rect 12759 13212 39580 13240
rect 12759 13209 12771 13212
rect 12713 13203 12771 13209
rect 39574 13200 39580 13212
rect 39632 13200 39638 13252
rect 41414 13200 41420 13252
rect 41472 13240 41478 13252
rect 61470 13240 61476 13252
rect 41472 13212 61476 13240
rect 41472 13200 41478 13212
rect 61470 13200 61476 13212
rect 61528 13200 61534 13252
rect 66622 13200 66628 13252
rect 66680 13240 66686 13252
rect 88242 13240 88248 13252
rect 66680 13212 88248 13240
rect 66680 13200 66686 13212
rect 88242 13200 88248 13212
rect 88300 13200 88306 13252
rect 16942 13172 16948 13184
rect 11716 13144 12664 13172
rect 16903 13144 16948 13172
rect 16942 13132 16948 13144
rect 17000 13132 17006 13184
rect 27709 13175 27767 13181
rect 27709 13141 27721 13175
rect 27755 13172 27767 13175
rect 28902 13172 28908 13184
rect 27755 13144 28908 13172
rect 27755 13141 27767 13144
rect 27709 13135 27767 13141
rect 28902 13132 28908 13144
rect 28960 13132 28966 13184
rect 52181 13175 52239 13181
rect 52181 13141 52193 13175
rect 52227 13172 52239 13175
rect 63770 13172 63776 13184
rect 52227 13144 63776 13172
rect 52227 13141 52239 13144
rect 52181 13135 52239 13141
rect 63770 13132 63776 13144
rect 63828 13132 63834 13184
rect 66346 13132 66352 13184
rect 66404 13172 66410 13184
rect 92198 13172 92204 13184
rect 66404 13144 92204 13172
rect 66404 13132 66410 13144
rect 92198 13132 92204 13144
rect 92256 13132 92262 13184
rect 1104 13082 98808 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 65686 13082
rect 65738 13030 65750 13082
rect 65802 13030 65814 13082
rect 65866 13030 65878 13082
rect 65930 13030 96406 13082
rect 96458 13030 96470 13082
rect 96522 13030 96534 13082
rect 96586 13030 96598 13082
rect 96650 13030 98808 13082
rect 1104 13008 98808 13030
rect 37182 12928 37188 12980
rect 37240 12968 37246 12980
rect 55950 12968 55956 12980
rect 37240 12940 55956 12968
rect 37240 12928 37246 12940
rect 55950 12928 55956 12940
rect 56008 12928 56014 12980
rect 60090 12928 60096 12980
rect 60148 12968 60154 12980
rect 60148 12940 69704 12968
rect 60148 12928 60154 12940
rect 6086 12860 6092 12912
rect 6144 12900 6150 12912
rect 6822 12900 6828 12912
rect 6144 12872 6828 12900
rect 6144 12860 6150 12872
rect 6822 12860 6828 12872
rect 6880 12900 6886 12912
rect 40589 12903 40647 12909
rect 40589 12900 40601 12903
rect 6880 12872 40601 12900
rect 6880 12860 6886 12872
rect 40589 12869 40601 12872
rect 40635 12900 40647 12903
rect 40911 12903 40969 12909
rect 40911 12900 40923 12903
rect 40635 12872 40923 12900
rect 40635 12869 40647 12872
rect 40589 12863 40647 12869
rect 40911 12869 40923 12872
rect 40957 12869 40969 12903
rect 41046 12900 41052 12912
rect 41007 12872 41052 12900
rect 40911 12863 40969 12869
rect 41046 12860 41052 12872
rect 41104 12860 41110 12912
rect 41156 12872 41552 12900
rect 41156 12844 41184 12872
rect 32490 12832 32496 12844
rect 18432 12804 32496 12832
rect 18432 12773 18460 12804
rect 32490 12792 32496 12804
rect 32548 12792 32554 12844
rect 41138 12832 41144 12844
rect 41051 12804 41144 12832
rect 41138 12792 41144 12804
rect 41196 12792 41202 12844
rect 41524 12832 41552 12872
rect 41598 12860 41604 12912
rect 41656 12900 41662 12912
rect 41656 12872 53144 12900
rect 41656 12860 41662 12872
rect 41524 12804 41736 12832
rect 18417 12767 18475 12773
rect 18417 12733 18429 12767
rect 18463 12733 18475 12767
rect 19058 12764 19064 12776
rect 19019 12736 19064 12764
rect 18417 12727 18475 12733
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 23106 12724 23112 12776
rect 23164 12764 23170 12776
rect 41598 12764 41604 12776
rect 23164 12736 41604 12764
rect 23164 12724 23170 12736
rect 41598 12724 41604 12736
rect 41656 12724 41662 12776
rect 41708 12773 41736 12804
rect 41693 12767 41751 12773
rect 41693 12733 41705 12767
rect 41739 12764 41751 12767
rect 53116 12764 53144 12872
rect 56134 12860 56140 12912
rect 56192 12900 56198 12912
rect 69201 12903 69259 12909
rect 69201 12900 69213 12903
rect 56192 12872 69213 12900
rect 56192 12860 56198 12872
rect 69201 12869 69213 12872
rect 69247 12869 69259 12903
rect 69676 12900 69704 12940
rect 69750 12928 69756 12980
rect 69808 12968 69814 12980
rect 69808 12940 97488 12968
rect 69808 12928 69814 12940
rect 69676 12872 97028 12900
rect 69201 12863 69259 12869
rect 55950 12792 55956 12844
rect 56008 12832 56014 12844
rect 96617 12835 96675 12841
rect 96617 12832 96629 12835
rect 56008 12804 96629 12832
rect 56008 12792 56014 12804
rect 96617 12801 96629 12804
rect 96663 12832 96675 12835
rect 96893 12835 96951 12841
rect 96893 12832 96905 12835
rect 96663 12804 96905 12832
rect 96663 12801 96675 12804
rect 96617 12795 96675 12801
rect 96893 12801 96905 12804
rect 96939 12801 96951 12835
rect 96893 12795 96951 12801
rect 56134 12764 56140 12776
rect 41739 12736 48314 12764
rect 53116 12736 56140 12764
rect 41739 12733 41751 12736
rect 41693 12727 41751 12733
rect 40770 12696 40776 12708
rect 40731 12668 40776 12696
rect 40770 12656 40776 12668
rect 40828 12656 40834 12708
rect 41509 12699 41567 12705
rect 41509 12665 41521 12699
rect 41555 12696 41567 12699
rect 48286 12696 48314 12736
rect 56134 12724 56140 12736
rect 56192 12724 56198 12776
rect 66257 12767 66315 12773
rect 66257 12733 66269 12767
rect 66303 12764 66315 12767
rect 66346 12764 66352 12776
rect 66303 12736 66352 12764
rect 66303 12733 66315 12736
rect 66257 12727 66315 12733
rect 66346 12724 66352 12736
rect 66404 12724 66410 12776
rect 66622 12764 66628 12776
rect 66583 12736 66628 12764
rect 66622 12724 66628 12736
rect 66680 12724 66686 12776
rect 66717 12767 66775 12773
rect 66717 12733 66729 12767
rect 66763 12764 66775 12767
rect 66806 12764 66812 12776
rect 66763 12736 66812 12764
rect 66763 12733 66775 12736
rect 66717 12727 66775 12733
rect 66806 12724 66812 12736
rect 66864 12724 66870 12776
rect 66990 12764 66996 12776
rect 66951 12736 66996 12764
rect 66990 12724 66996 12736
rect 67048 12724 67054 12776
rect 67082 12724 67088 12776
rect 67140 12764 67146 12776
rect 67177 12767 67235 12773
rect 67177 12764 67189 12767
rect 67140 12736 67189 12764
rect 67140 12724 67146 12736
rect 67177 12733 67189 12736
rect 67223 12733 67235 12767
rect 67542 12764 67548 12776
rect 67503 12736 67548 12764
rect 67177 12727 67235 12733
rect 67542 12724 67548 12736
rect 67600 12724 67606 12776
rect 69201 12767 69259 12773
rect 69201 12733 69213 12767
rect 69247 12764 69259 12767
rect 96706 12764 96712 12776
rect 69247 12736 89714 12764
rect 96667 12736 96712 12764
rect 69247 12733 69259 12736
rect 69201 12727 69259 12733
rect 82538 12696 82544 12708
rect 41555 12668 46244 12696
rect 48286 12668 82544 12696
rect 41555 12665 41567 12668
rect 41509 12659 41567 12665
rect 29730 12588 29736 12640
rect 29788 12628 29794 12640
rect 41046 12628 41052 12640
rect 29788 12600 41052 12628
rect 29788 12588 29794 12600
rect 41046 12588 41052 12600
rect 41104 12588 41110 12640
rect 46216 12628 46244 12668
rect 82538 12656 82544 12668
rect 82596 12656 82602 12708
rect 89686 12696 89714 12736
rect 96706 12724 96712 12736
rect 96764 12724 96770 12776
rect 97000 12764 97028 12872
rect 97460 12773 97488 12940
rect 97810 12900 97816 12912
rect 97771 12872 97816 12900
rect 97810 12860 97816 12872
rect 97868 12860 97874 12912
rect 97077 12767 97135 12773
rect 97077 12764 97089 12767
rect 97000 12736 97089 12764
rect 97077 12733 97089 12736
rect 97123 12733 97135 12767
rect 97077 12727 97135 12733
rect 97353 12767 97411 12773
rect 97353 12733 97365 12767
rect 97399 12733 97411 12767
rect 97353 12727 97411 12733
rect 97445 12767 97503 12773
rect 97445 12733 97457 12767
rect 97491 12733 97503 12767
rect 97445 12727 97503 12733
rect 97368 12696 97396 12727
rect 89686 12668 97396 12696
rect 84470 12628 84476 12640
rect 46216 12600 84476 12628
rect 84470 12588 84476 12600
rect 84528 12588 84534 12640
rect 1104 12538 98808 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 50326 12538
rect 50378 12486 50390 12538
rect 50442 12486 50454 12538
rect 50506 12486 50518 12538
rect 50570 12486 81046 12538
rect 81098 12486 81110 12538
rect 81162 12486 81174 12538
rect 81226 12486 81238 12538
rect 81290 12486 98808 12538
rect 1104 12464 98808 12486
rect 27706 12384 27712 12436
rect 27764 12424 27770 12436
rect 27982 12424 27988 12436
rect 27764 12396 27988 12424
rect 27764 12384 27770 12396
rect 27982 12384 27988 12396
rect 28040 12384 28046 12436
rect 63678 12424 63684 12436
rect 45526 12396 63684 12424
rect 38102 12288 38108 12300
rect 38063 12260 38108 12288
rect 38102 12248 38108 12260
rect 38160 12248 38166 12300
rect 38381 12291 38439 12297
rect 38381 12257 38393 12291
rect 38427 12288 38439 12291
rect 45526 12288 45554 12396
rect 63678 12384 63684 12396
rect 63736 12384 63742 12436
rect 67634 12384 67640 12436
rect 67692 12424 67698 12436
rect 67692 12396 96752 12424
rect 67692 12384 67698 12396
rect 67726 12316 67732 12368
rect 67784 12356 67790 12368
rect 67784 12328 89714 12356
rect 67784 12316 67790 12328
rect 38427 12260 45554 12288
rect 38427 12257 38439 12260
rect 38381 12251 38439 12257
rect 85666 12248 85672 12300
rect 85724 12288 85730 12300
rect 85761 12291 85819 12297
rect 85761 12288 85773 12291
rect 85724 12260 85773 12288
rect 85724 12248 85730 12260
rect 85761 12257 85773 12260
rect 85807 12257 85819 12291
rect 85761 12251 85819 12257
rect 85850 12248 85856 12300
rect 85908 12288 85914 12300
rect 85945 12291 86003 12297
rect 85945 12288 85957 12291
rect 85908 12260 85957 12288
rect 85908 12248 85914 12260
rect 85945 12257 85957 12260
rect 85991 12257 86003 12291
rect 85945 12251 86003 12257
rect 86129 12291 86187 12297
rect 86129 12257 86141 12291
rect 86175 12257 86187 12291
rect 86494 12288 86500 12300
rect 86455 12260 86500 12288
rect 86129 12251 86187 12257
rect 82170 12180 82176 12232
rect 82228 12220 82234 12232
rect 86144 12220 86172 12251
rect 86494 12248 86500 12260
rect 86552 12248 86558 12300
rect 86402 12220 86408 12232
rect 82228 12192 86172 12220
rect 86363 12192 86408 12220
rect 82228 12180 82234 12192
rect 86402 12180 86408 12192
rect 86460 12180 86466 12232
rect 3050 12112 3056 12164
rect 3108 12152 3114 12164
rect 86865 12155 86923 12161
rect 86865 12152 86877 12155
rect 3108 12124 26234 12152
rect 3108 12112 3114 12124
rect 26206 12084 26234 12124
rect 39592 12124 86877 12152
rect 39592 12084 39620 12124
rect 86865 12121 86877 12124
rect 86911 12121 86923 12155
rect 89686 12152 89714 12328
rect 95234 12248 95240 12300
rect 95292 12288 95298 12300
rect 96724 12297 96752 12396
rect 96341 12291 96399 12297
rect 96341 12288 96353 12291
rect 95292 12260 96353 12288
rect 95292 12248 95298 12260
rect 96341 12257 96353 12260
rect 96387 12257 96399 12291
rect 96341 12251 96399 12257
rect 96709 12291 96767 12297
rect 96709 12257 96721 12291
rect 96755 12257 96767 12291
rect 96709 12251 96767 12257
rect 97077 12291 97135 12297
rect 97077 12257 97089 12291
rect 97123 12257 97135 12291
rect 97077 12251 97135 12257
rect 96798 12220 96804 12232
rect 96759 12192 96804 12220
rect 96798 12180 96804 12192
rect 96856 12180 96862 12232
rect 96982 12220 96988 12232
rect 96943 12192 96988 12220
rect 96982 12180 96988 12192
rect 97040 12180 97046 12232
rect 97092 12152 97120 12251
rect 89686 12124 97120 12152
rect 86865 12115 86923 12121
rect 26206 12056 39620 12084
rect 39669 12087 39727 12093
rect 39669 12053 39681 12087
rect 39715 12084 39727 12087
rect 63586 12084 63592 12096
rect 39715 12056 63592 12084
rect 39715 12053 39727 12056
rect 39669 12047 39727 12053
rect 63586 12044 63592 12056
rect 63644 12044 63650 12096
rect 77110 12044 77116 12096
rect 77168 12084 77174 12096
rect 80698 12084 80704 12096
rect 77168 12056 80704 12084
rect 77168 12044 77174 12056
rect 80698 12044 80704 12056
rect 80756 12044 80762 12096
rect 97534 12084 97540 12096
rect 97495 12056 97540 12084
rect 97534 12044 97540 12056
rect 97592 12044 97598 12096
rect 1104 11994 98808 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 65686 11994
rect 65738 11942 65750 11994
rect 65802 11942 65814 11994
rect 65866 11942 65878 11994
rect 65930 11942 96406 11994
rect 96458 11942 96470 11994
rect 96522 11942 96534 11994
rect 96586 11942 96598 11994
rect 96650 11942 98808 11994
rect 1104 11920 98808 11942
rect 3418 11880 3424 11892
rect 3379 11852 3424 11880
rect 3418 11840 3424 11852
rect 3476 11840 3482 11892
rect 30190 11840 30196 11892
rect 30248 11880 30254 11892
rect 97534 11880 97540 11892
rect 30248 11852 97540 11880
rect 30248 11840 30254 11852
rect 97534 11840 97540 11852
rect 97592 11840 97598 11892
rect 19521 11815 19579 11821
rect 19521 11781 19533 11815
rect 19567 11812 19579 11815
rect 20622 11812 20628 11824
rect 19567 11784 20628 11812
rect 19567 11781 19579 11784
rect 19521 11775 19579 11781
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 48222 11772 48228 11824
rect 48280 11812 48286 11824
rect 80379 11815 80437 11821
rect 80379 11812 80391 11815
rect 48280 11784 80391 11812
rect 48280 11772 48286 11784
rect 80379 11781 80391 11784
rect 80425 11781 80437 11815
rect 80514 11812 80520 11824
rect 80475 11784 80520 11812
rect 80379 11775 80437 11781
rect 80514 11772 80520 11784
rect 80572 11772 80578 11824
rect 80698 11772 80704 11824
rect 80756 11812 80762 11824
rect 85298 11812 85304 11824
rect 80756 11784 85304 11812
rect 80756 11772 80762 11784
rect 85298 11772 85304 11784
rect 85356 11772 85362 11824
rect 3694 11744 3700 11756
rect 3655 11716 3700 11744
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 3835 11716 12434 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 3970 11685 3976 11688
rect 3513 11679 3571 11685
rect 3513 11645 3525 11679
rect 3559 11645 3571 11679
rect 3513 11639 3571 11645
rect 3917 11679 3976 11685
rect 3917 11645 3929 11679
rect 3963 11645 3976 11679
rect 3917 11639 3976 11645
rect 3237 11611 3295 11617
rect 3237 11577 3249 11611
rect 3283 11608 3295 11611
rect 3528 11608 3556 11639
rect 3970 11636 3976 11639
rect 4028 11636 4034 11688
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11676 4123 11679
rect 12066 11676 12072 11688
rect 4111 11648 12072 11676
rect 4111 11645 4123 11648
rect 4065 11639 4123 11645
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 12406 11676 12434 11716
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 35342 11744 35348 11756
rect 18012 11716 35348 11744
rect 18012 11704 18018 11716
rect 35342 11704 35348 11716
rect 35400 11704 35406 11756
rect 41230 11704 41236 11756
rect 41288 11744 41294 11756
rect 53834 11744 53840 11756
rect 41288 11716 53840 11744
rect 41288 11704 41294 11716
rect 53834 11704 53840 11716
rect 53892 11704 53898 11756
rect 79965 11747 80023 11753
rect 79965 11744 79977 11747
rect 77220 11716 79977 11744
rect 77110 11676 77116 11688
rect 12406 11648 77116 11676
rect 77110 11636 77116 11648
rect 77168 11636 77174 11688
rect 17954 11608 17960 11620
rect 3283 11580 17960 11608
rect 3283 11577 3295 11580
rect 3237 11571 3295 11577
rect 17954 11568 17960 11580
rect 18012 11568 18018 11620
rect 27706 11568 27712 11620
rect 27764 11608 27770 11620
rect 33778 11608 33784 11620
rect 27764 11580 33784 11608
rect 27764 11568 27770 11580
rect 33778 11568 33784 11580
rect 33836 11568 33842 11620
rect 37550 11568 37556 11620
rect 37608 11608 37614 11620
rect 44174 11608 44180 11620
rect 37608 11580 44180 11608
rect 37608 11568 37614 11580
rect 44174 11568 44180 11580
rect 44232 11568 44238 11620
rect 51074 11568 51080 11620
rect 51132 11608 51138 11620
rect 51994 11608 52000 11620
rect 51132 11580 52000 11608
rect 51132 11568 51138 11580
rect 51994 11568 52000 11580
rect 52052 11608 52058 11620
rect 77220 11608 77248 11716
rect 79965 11713 79977 11716
rect 80011 11744 80023 11747
rect 80057 11747 80115 11753
rect 80057 11744 80069 11747
rect 80011 11716 80069 11744
rect 80011 11713 80023 11716
rect 79965 11707 80023 11713
rect 80057 11713 80069 11716
rect 80103 11713 80115 11747
rect 80057 11707 80115 11713
rect 80609 11747 80667 11753
rect 80609 11713 80621 11747
rect 80655 11744 80667 11747
rect 80882 11744 80888 11756
rect 80655 11716 80888 11744
rect 80655 11713 80667 11716
rect 80609 11707 80667 11713
rect 80882 11704 80888 11716
rect 80940 11704 80946 11756
rect 52052 11580 77248 11608
rect 77312 11648 84194 11676
rect 52052 11568 52058 11580
rect 31662 11500 31668 11552
rect 31720 11540 31726 11552
rect 77312 11540 77340 11648
rect 79965 11611 80023 11617
rect 79965 11577 79977 11611
rect 80011 11608 80023 11611
rect 80241 11611 80299 11617
rect 80241 11608 80253 11611
rect 80011 11580 80253 11608
rect 80011 11577 80023 11580
rect 79965 11571 80023 11577
rect 80241 11577 80253 11580
rect 80287 11577 80299 11611
rect 80241 11571 80299 11577
rect 80882 11540 80888 11552
rect 31720 11512 77340 11540
rect 80843 11512 80888 11540
rect 31720 11500 31726 11512
rect 80882 11500 80888 11512
rect 80940 11500 80946 11552
rect 84166 11540 84194 11648
rect 96982 11540 96988 11552
rect 84166 11512 96988 11540
rect 96982 11500 96988 11512
rect 97040 11500 97046 11552
rect 1104 11450 98808 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 50326 11450
rect 50378 11398 50390 11450
rect 50442 11398 50454 11450
rect 50506 11398 50518 11450
rect 50570 11398 81046 11450
rect 81098 11398 81110 11450
rect 81162 11398 81174 11450
rect 81226 11398 81238 11450
rect 81290 11398 98808 11450
rect 1104 11376 98808 11398
rect 26973 11339 27031 11345
rect 26973 11305 26985 11339
rect 27019 11336 27031 11339
rect 89346 11336 89352 11348
rect 27019 11308 89352 11336
rect 27019 11305 27031 11308
rect 26973 11299 27031 11305
rect 89346 11296 89352 11308
rect 89404 11296 89410 11348
rect 8754 11228 8760 11280
rect 8812 11268 8818 11280
rect 27982 11268 27988 11280
rect 8812 11240 27384 11268
rect 8812 11228 8818 11240
rect 27154 11200 27160 11212
rect 26206 11172 26924 11200
rect 27115 11172 27160 11200
rect 5718 11132 5724 11144
rect 5679 11104 5724 11132
rect 5718 11092 5724 11104
rect 5776 11092 5782 11144
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11132 6055 11135
rect 26206 11132 26234 11172
rect 6043 11104 26234 11132
rect 26896 11132 26924 11172
rect 27154 11160 27160 11172
rect 27212 11160 27218 11212
rect 27356 11209 27384 11240
rect 27908 11240 27988 11268
rect 27341 11203 27399 11209
rect 27341 11169 27353 11203
rect 27387 11169 27399 11203
rect 27706 11200 27712 11212
rect 27667 11172 27712 11200
rect 27341 11163 27399 11169
rect 27706 11160 27712 11172
rect 27764 11160 27770 11212
rect 27908 11209 27936 11240
rect 27982 11228 27988 11240
rect 28040 11228 28046 11280
rect 44450 11228 44456 11280
rect 44508 11268 44514 11280
rect 47210 11268 47216 11280
rect 44508 11240 47216 11268
rect 44508 11228 44514 11240
rect 47210 11228 47216 11240
rect 47268 11268 47274 11280
rect 48222 11268 48228 11280
rect 47268 11240 48228 11268
rect 47268 11228 47274 11240
rect 48222 11228 48228 11240
rect 48280 11228 48286 11280
rect 50798 11228 50804 11280
rect 50856 11268 50862 11280
rect 80790 11268 80796 11280
rect 50856 11240 53604 11268
rect 50856 11228 50862 11240
rect 27893 11203 27951 11209
rect 27893 11169 27905 11203
rect 27939 11169 27951 11203
rect 37366 11200 37372 11212
rect 27893 11163 27951 11169
rect 35866 11172 37372 11200
rect 35866 11132 35894 11172
rect 37366 11160 37372 11172
rect 37424 11160 37430 11212
rect 42794 11160 42800 11212
rect 42852 11200 42858 11212
rect 42889 11203 42947 11209
rect 42889 11200 42901 11203
rect 42852 11172 42901 11200
rect 42852 11160 42858 11172
rect 42889 11169 42901 11172
rect 42935 11200 42947 11203
rect 44082 11200 44088 11212
rect 42935 11172 44088 11200
rect 42935 11169 42947 11172
rect 42889 11163 42947 11169
rect 44082 11160 44088 11172
rect 44140 11160 44146 11212
rect 44174 11160 44180 11212
rect 44232 11200 44238 11212
rect 53576 11209 53604 11240
rect 53668 11240 80796 11268
rect 53377 11203 53435 11209
rect 53377 11200 53389 11203
rect 44232 11172 53389 11200
rect 44232 11160 44238 11172
rect 53377 11169 53389 11172
rect 53423 11169 53435 11203
rect 53377 11163 53435 11169
rect 53561 11203 53619 11209
rect 53561 11169 53573 11203
rect 53607 11169 53619 11203
rect 53561 11163 53619 11169
rect 26896 11104 35894 11132
rect 43165 11135 43223 11141
rect 6043 11101 6055 11104
rect 5997 11095 6055 11101
rect 43165 11101 43177 11135
rect 43211 11132 43223 11135
rect 47486 11132 47492 11144
rect 43211 11104 47492 11132
rect 43211 11101 43223 11104
rect 43165 11095 43223 11101
rect 47486 11092 47492 11104
rect 47544 11092 47550 11144
rect 7285 11067 7343 11073
rect 7285 11033 7297 11067
rect 7331 11064 7343 11067
rect 38010 11064 38016 11076
rect 7331 11036 38016 11064
rect 7331 11033 7343 11036
rect 7285 11027 7343 11033
rect 38010 11024 38016 11036
rect 38068 11024 38074 11076
rect 44192 11036 44404 11064
rect 19150 10956 19156 11008
rect 19208 10996 19214 11008
rect 44192 10996 44220 11036
rect 19208 10968 44220 10996
rect 44376 10996 44404 11036
rect 44450 11024 44456 11076
rect 44508 11064 44514 11076
rect 53190 11064 53196 11076
rect 44508 11036 44553 11064
rect 53151 11036 53196 11064
rect 44508 11024 44514 11036
rect 53190 11024 53196 11036
rect 53248 11064 53254 11076
rect 53668 11064 53696 11240
rect 53834 11200 53840 11212
rect 53795 11172 53840 11200
rect 53834 11160 53840 11172
rect 53892 11160 53898 11212
rect 53944 11209 53972 11240
rect 80790 11228 80796 11240
rect 80848 11228 80854 11280
rect 53930 11203 53988 11209
rect 53930 11169 53942 11203
rect 53976 11169 53988 11203
rect 53930 11163 53988 11169
rect 54113 11203 54171 11209
rect 54113 11169 54125 11203
rect 54159 11200 54171 11203
rect 54294 11200 54300 11212
rect 54159 11172 54300 11200
rect 54159 11169 54171 11172
rect 54113 11163 54171 11169
rect 54294 11160 54300 11172
rect 54352 11160 54358 11212
rect 53745 11135 53803 11141
rect 53745 11101 53757 11135
rect 53791 11101 53803 11135
rect 53852 11132 53880 11160
rect 55030 11132 55036 11144
rect 53852 11104 55036 11132
rect 53745 11095 53803 11101
rect 53248 11036 53696 11064
rect 53760 11064 53788 11095
rect 55030 11092 55036 11104
rect 55088 11092 55094 11144
rect 55214 11064 55220 11076
rect 53760 11036 55220 11064
rect 53248 11024 53254 11036
rect 55214 11024 55220 11036
rect 55272 11024 55278 11076
rect 51074 10996 51080 11008
rect 44376 10968 51080 10996
rect 19208 10956 19214 10968
rect 51074 10956 51080 10968
rect 51132 10956 51138 11008
rect 1104 10906 98808 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 65686 10906
rect 65738 10854 65750 10906
rect 65802 10854 65814 10906
rect 65866 10854 65878 10906
rect 65930 10854 96406 10906
rect 96458 10854 96470 10906
rect 96522 10854 96534 10906
rect 96586 10854 96598 10906
rect 96650 10854 98808 10906
rect 1104 10832 98808 10854
rect 5718 10792 5724 10804
rect 1688 10764 5724 10792
rect 1688 10665 1716 10764
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 55214 10792 55220 10804
rect 17000 10764 55220 10792
rect 17000 10752 17006 10764
rect 55214 10752 55220 10764
rect 55272 10752 55278 10804
rect 14458 10724 14464 10736
rect 4448 10696 14464 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10625 1731 10659
rect 3878 10656 3884 10668
rect 3839 10628 3884 10656
rect 1673 10619 1731 10625
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 1946 10588 1952 10600
rect 1907 10560 1952 10588
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 4448 10597 4476 10696
rect 14458 10684 14464 10696
rect 14516 10684 14522 10736
rect 36909 10727 36967 10733
rect 36909 10693 36921 10727
rect 36955 10724 36967 10727
rect 78858 10724 78864 10736
rect 36955 10696 78864 10724
rect 36955 10693 36967 10696
rect 36909 10687 36967 10693
rect 78858 10684 78864 10696
rect 78916 10684 78922 10736
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 6178 10656 6184 10668
rect 4525 10619 4583 10625
rect 4816 10628 6184 10656
rect 4433 10591 4491 10597
rect 4433 10557 4445 10591
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 4540 10520 4568 10619
rect 4816 10597 4844 10628
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 12894 10656 12900 10668
rect 8628 10628 12434 10656
rect 12855 10628 12900 10656
rect 8628 10616 8634 10628
rect 4801 10591 4859 10597
rect 4801 10557 4813 10591
rect 4847 10557 4859 10591
rect 4801 10551 4859 10557
rect 4985 10591 5043 10597
rect 4985 10557 4997 10591
rect 5031 10588 5043 10591
rect 6638 10588 6644 10600
rect 5031 10560 6644 10588
rect 5031 10557 5043 10560
rect 4985 10551 5043 10557
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 12069 10591 12127 10597
rect 12069 10557 12081 10591
rect 12115 10557 12127 10591
rect 12406 10588 12434 10628
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 39853 10659 39911 10665
rect 22066 10628 39804 10656
rect 22066 10588 22094 10628
rect 24026 10588 24032 10600
rect 12406 10560 22094 10588
rect 23987 10560 24032 10588
rect 12069 10551 12127 10557
rect 11330 10520 11336 10532
rect 4540 10492 11336 10520
rect 11330 10480 11336 10492
rect 11388 10520 11394 10532
rect 12084 10520 12112 10551
rect 24026 10548 24032 10560
rect 24084 10548 24090 10600
rect 24302 10548 24308 10600
rect 24360 10588 24366 10600
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 24360 10560 24685 10588
rect 24360 10548 24366 10560
rect 24673 10557 24685 10560
rect 24719 10557 24731 10591
rect 36354 10588 36360 10600
rect 36315 10560 36360 10588
rect 24673 10551 24731 10557
rect 36354 10548 36360 10560
rect 36412 10548 36418 10600
rect 36630 10588 36636 10600
rect 36591 10560 36636 10588
rect 36630 10548 36636 10560
rect 36688 10548 36694 10600
rect 36722 10548 36728 10600
rect 36780 10597 36786 10600
rect 36780 10588 36788 10597
rect 39776 10588 39804 10628
rect 39853 10625 39865 10659
rect 39899 10656 39911 10659
rect 40129 10659 40187 10665
rect 40129 10656 40141 10659
rect 39899 10628 40141 10656
rect 39899 10625 39911 10628
rect 39853 10619 39911 10625
rect 40129 10625 40141 10628
rect 40175 10656 40187 10659
rect 93210 10656 93216 10668
rect 40175 10628 93216 10656
rect 40175 10625 40187 10628
rect 40129 10619 40187 10625
rect 93210 10616 93216 10628
rect 93268 10616 93274 10668
rect 36780 10560 36825 10588
rect 39776 10560 45554 10588
rect 36780 10551 36788 10560
rect 36780 10548 36786 10551
rect 11388 10492 12112 10520
rect 36541 10523 36599 10529
rect 11388 10480 11394 10492
rect 36541 10489 36553 10523
rect 36587 10520 36599 10523
rect 40678 10520 40684 10532
rect 36587 10492 40684 10520
rect 36587 10489 36599 10492
rect 36541 10483 36599 10489
rect 40678 10480 40684 10492
rect 40736 10480 40742 10532
rect 45526 10520 45554 10560
rect 54294 10548 54300 10600
rect 54352 10588 54358 10600
rect 54665 10591 54723 10597
rect 54665 10588 54677 10591
rect 54352 10560 54677 10588
rect 54352 10548 54358 10560
rect 54665 10557 54677 10560
rect 54711 10557 54723 10591
rect 54665 10551 54723 10557
rect 54849 10591 54907 10597
rect 54849 10557 54861 10591
rect 54895 10557 54907 10591
rect 55030 10588 55036 10600
rect 54991 10560 55036 10588
rect 54849 10551 54907 10557
rect 54481 10523 54539 10529
rect 54481 10520 54493 10523
rect 45526 10492 54493 10520
rect 54481 10489 54493 10492
rect 54527 10520 54539 10523
rect 54864 10520 54892 10551
rect 55030 10548 55036 10560
rect 55088 10548 55094 10600
rect 55306 10548 55312 10600
rect 55364 10588 55370 10600
rect 55401 10591 55459 10597
rect 55401 10588 55413 10591
rect 55364 10560 55413 10588
rect 55364 10548 55370 10560
rect 55401 10557 55413 10560
rect 55447 10557 55459 10591
rect 55582 10588 55588 10600
rect 55543 10560 55588 10588
rect 55401 10551 55459 10557
rect 55582 10548 55588 10560
rect 55640 10548 55646 10600
rect 75178 10520 75184 10532
rect 54527 10492 75184 10520
rect 54527 10489 54539 10492
rect 54481 10483 54539 10489
rect 75178 10480 75184 10492
rect 75236 10480 75242 10532
rect 3237 10455 3295 10461
rect 3237 10421 3249 10455
rect 3283 10452 3295 10455
rect 13170 10452 13176 10464
rect 3283 10424 13176 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 30098 10412 30104 10464
rect 30156 10452 30162 10464
rect 38194 10452 38200 10464
rect 30156 10424 38200 10452
rect 30156 10412 30162 10424
rect 38194 10412 38200 10424
rect 38252 10412 38258 10464
rect 55861 10455 55919 10461
rect 55861 10421 55873 10455
rect 55907 10452 55919 10455
rect 93578 10452 93584 10464
rect 55907 10424 93584 10452
rect 55907 10421 55919 10424
rect 55861 10415 55919 10421
rect 93578 10412 93584 10424
rect 93636 10412 93642 10464
rect 1104 10362 98808 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 50326 10362
rect 50378 10310 50390 10362
rect 50442 10310 50454 10362
rect 50506 10310 50518 10362
rect 50570 10310 81046 10362
rect 81098 10310 81110 10362
rect 81162 10310 81174 10362
rect 81226 10310 81238 10362
rect 81290 10310 98808 10362
rect 1104 10288 98808 10310
rect 17129 10251 17187 10257
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 17175 10220 19656 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 4798 10140 4804 10192
rect 4856 10180 4862 10192
rect 19628 10180 19656 10220
rect 20622 10208 20628 10260
rect 20680 10248 20686 10260
rect 40218 10248 40224 10260
rect 20680 10220 40224 10248
rect 20680 10208 20686 10220
rect 40218 10208 40224 10220
rect 40276 10208 40282 10260
rect 61746 10248 61752 10260
rect 61707 10220 61752 10248
rect 61746 10208 61752 10220
rect 61804 10208 61810 10260
rect 62206 10248 62212 10260
rect 62167 10220 62212 10248
rect 62206 10208 62212 10220
rect 62264 10208 62270 10260
rect 62684 10220 63540 10248
rect 4856 10152 17356 10180
rect 19628 10152 26234 10180
rect 4856 10140 4862 10152
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10112 17187 10115
rect 17221 10115 17279 10121
rect 17221 10112 17233 10115
rect 17175 10084 17233 10112
rect 17175 10081 17187 10084
rect 17129 10075 17187 10081
rect 17221 10081 17233 10084
rect 17267 10081 17279 10115
rect 17328 10112 17356 10152
rect 23569 10115 23627 10121
rect 23569 10112 23581 10115
rect 17328 10084 23581 10112
rect 17221 10075 17279 10081
rect 23569 10081 23581 10084
rect 23615 10081 23627 10115
rect 26206 10112 26234 10152
rect 35526 10140 35532 10192
rect 35584 10180 35590 10192
rect 39942 10180 39948 10192
rect 35584 10152 39948 10180
rect 35584 10140 35590 10152
rect 39942 10140 39948 10152
rect 40000 10140 40006 10192
rect 61764 10180 61792 10208
rect 62684 10180 62712 10220
rect 61764 10152 62712 10180
rect 63319 10115 63377 10121
rect 26206 10084 63080 10112
rect 23569 10075 23627 10081
rect 17560 10047 17618 10053
rect 17560 10044 17572 10047
rect 17236 10016 17572 10044
rect 17236 9988 17264 10016
rect 17560 10013 17572 10016
rect 17606 10013 17618 10047
rect 17560 10007 17618 10013
rect 17678 10004 17684 10056
rect 17736 10044 17742 10056
rect 62942 10044 62948 10056
rect 17736 10016 62948 10044
rect 17736 10004 17742 10016
rect 62942 10004 62948 10016
rect 63000 10004 63006 10056
rect 63052 10044 63080 10084
rect 63319 10081 63331 10115
rect 63365 10112 63377 10115
rect 63512 10112 63540 10220
rect 63678 10140 63684 10192
rect 63736 10180 63742 10192
rect 63736 10152 67634 10180
rect 63736 10140 63742 10152
rect 63365 10084 63540 10112
rect 63582 10115 63640 10121
rect 63365 10081 63377 10084
rect 63319 10075 63377 10081
rect 63582 10081 63594 10115
rect 63628 10081 63640 10115
rect 67606 10112 67634 10152
rect 80882 10112 80888 10124
rect 67606 10084 80888 10112
rect 63582 10075 63640 10081
rect 63402 10044 63408 10056
rect 63052 10016 63408 10044
rect 63402 10004 63408 10016
rect 63460 10004 63466 10056
rect 63604 9988 63632 10075
rect 80882 10072 80888 10084
rect 80940 10072 80946 10124
rect 91465 10115 91523 10121
rect 91465 10081 91477 10115
rect 91511 10112 91523 10115
rect 91741 10115 91799 10121
rect 91741 10112 91753 10115
rect 91511 10084 91753 10112
rect 91511 10081 91523 10084
rect 91465 10075 91523 10081
rect 91741 10081 91753 10084
rect 91787 10112 91799 10115
rect 93394 10112 93400 10124
rect 91787 10084 93400 10112
rect 91787 10081 91799 10084
rect 91741 10075 91799 10081
rect 93394 10072 93400 10084
rect 93452 10072 93458 10124
rect 63862 10004 63868 10056
rect 63920 10044 63926 10056
rect 92750 10044 92756 10056
rect 63920 10016 92756 10044
rect 63920 10004 63926 10016
rect 92750 10004 92756 10016
rect 92808 10004 92814 10056
rect 17218 9936 17224 9988
rect 17276 9936 17282 9988
rect 17386 9979 17444 9985
rect 17386 9945 17398 9979
rect 17432 9976 17444 9979
rect 17432 9948 62712 9976
rect 17432 9945 17444 9948
rect 17386 9939 17444 9945
rect 17497 9911 17555 9917
rect 17497 9877 17509 9911
rect 17543 9908 17555 9911
rect 17678 9908 17684 9920
rect 17543 9880 17684 9908
rect 17543 9877 17555 9880
rect 17497 9871 17555 9877
rect 17678 9868 17684 9880
rect 17736 9868 17742 9920
rect 17862 9908 17868 9920
rect 17823 9880 17868 9908
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 23753 9911 23811 9917
rect 23753 9877 23765 9911
rect 23799 9908 23811 9911
rect 24026 9908 24032 9920
rect 23799 9880 24032 9908
rect 23799 9877 23811 9880
rect 23753 9871 23811 9877
rect 24026 9868 24032 9880
rect 24084 9908 24090 9920
rect 24394 9908 24400 9920
rect 24084 9880 24400 9908
rect 24084 9868 24090 9880
rect 24394 9868 24400 9880
rect 24452 9868 24458 9920
rect 62684 9908 62712 9948
rect 63586 9936 63592 9988
rect 63644 9936 63650 9988
rect 94130 9976 94136 9988
rect 70366 9948 94136 9976
rect 70366 9908 70394 9948
rect 94130 9936 94136 9948
rect 94188 9936 94194 9988
rect 62684 9880 70394 9908
rect 1104 9818 98808 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 65686 9818
rect 65738 9766 65750 9818
rect 65802 9766 65814 9818
rect 65866 9766 65878 9818
rect 65930 9766 96406 9818
rect 96458 9766 96470 9818
rect 96522 9766 96534 9818
rect 96586 9766 96598 9818
rect 96650 9766 98808 9818
rect 1104 9744 98808 9766
rect 1946 9664 1952 9716
rect 2004 9704 2010 9716
rect 91002 9704 91008 9716
rect 2004 9676 91008 9704
rect 2004 9664 2010 9676
rect 91002 9664 91008 9676
rect 91060 9664 91066 9716
rect 48958 9636 48964 9648
rect 45112 9608 48964 9636
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 27062 9568 27068 9580
rect 13228 9540 27068 9568
rect 13228 9528 13234 9540
rect 27062 9528 27068 9540
rect 27120 9528 27126 9580
rect 23198 9460 23204 9512
rect 23256 9500 23262 9512
rect 44358 9500 44364 9512
rect 23256 9472 44364 9500
rect 23256 9460 23262 9472
rect 44358 9460 44364 9472
rect 44416 9460 44422 9512
rect 45112 9509 45140 9608
rect 48958 9596 48964 9608
rect 49016 9596 49022 9648
rect 92566 9596 92572 9648
rect 92624 9636 92630 9648
rect 94225 9639 94283 9645
rect 94225 9636 94237 9639
rect 92624 9608 94237 9636
rect 92624 9596 92630 9608
rect 94225 9605 94237 9608
rect 94271 9605 94283 9639
rect 94225 9599 94283 9605
rect 45480 9540 49280 9568
rect 45097 9503 45155 9509
rect 45097 9469 45109 9503
rect 45143 9469 45155 9503
rect 45278 9500 45284 9512
rect 45239 9472 45284 9500
rect 45097 9463 45155 9469
rect 45278 9460 45284 9472
rect 45336 9460 45342 9512
rect 45480 9509 45508 9540
rect 45465 9503 45523 9509
rect 45465 9469 45477 9503
rect 45511 9469 45523 9503
rect 45465 9463 45523 9469
rect 45646 9460 45652 9512
rect 45704 9500 45710 9512
rect 46477 9503 46535 9509
rect 46477 9500 46489 9503
rect 45704 9472 46489 9500
rect 45704 9460 45710 9472
rect 46477 9469 46489 9472
rect 46523 9469 46535 9503
rect 49252 9500 49280 9540
rect 53098 9528 53104 9580
rect 53156 9568 53162 9580
rect 58066 9568 58072 9580
rect 53156 9540 58072 9568
rect 53156 9528 53162 9540
rect 58066 9528 58072 9540
rect 58124 9528 58130 9580
rect 60182 9528 60188 9580
rect 60240 9568 60246 9580
rect 86402 9568 86408 9580
rect 60240 9540 86408 9568
rect 60240 9528 60246 9540
rect 86402 9528 86408 9540
rect 86460 9528 86466 9580
rect 55582 9500 55588 9512
rect 49252 9472 55588 9500
rect 46477 9463 46535 9469
rect 55582 9460 55588 9472
rect 55640 9460 55646 9512
rect 61105 9503 61163 9509
rect 61105 9469 61117 9503
rect 61151 9500 61163 9503
rect 63402 9500 63408 9512
rect 61151 9472 63408 9500
rect 61151 9469 61163 9472
rect 61105 9463 61163 9469
rect 63402 9460 63408 9472
rect 63460 9460 63466 9512
rect 68278 9460 68284 9512
rect 68336 9500 68342 9512
rect 92842 9500 92848 9512
rect 68336 9472 92848 9500
rect 68336 9460 68342 9472
rect 92842 9460 92848 9472
rect 92900 9460 92906 9512
rect 20530 9392 20536 9444
rect 20588 9432 20594 9444
rect 44450 9432 44456 9444
rect 20588 9404 44456 9432
rect 20588 9392 20594 9404
rect 44450 9392 44456 9404
rect 44508 9392 44514 9444
rect 44637 9435 44695 9441
rect 44637 9401 44649 9435
rect 44683 9432 44695 9435
rect 70762 9432 70768 9444
rect 44683 9404 70768 9432
rect 44683 9401 44695 9404
rect 44637 9395 44695 9401
rect 70762 9392 70768 9404
rect 70820 9392 70826 9444
rect 73798 9392 73804 9444
rect 73856 9432 73862 9444
rect 82814 9432 82820 9444
rect 73856 9404 82820 9432
rect 73856 9392 73862 9404
rect 82814 9392 82820 9404
rect 82872 9392 82878 9444
rect 94038 9432 94044 9444
rect 93951 9404 94044 9432
rect 94038 9392 94044 9404
rect 94096 9432 94102 9444
rect 94406 9432 94412 9444
rect 94096 9404 94412 9432
rect 94096 9392 94102 9404
rect 94406 9392 94412 9404
rect 94464 9392 94470 9444
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 40862 9364 40868 9376
rect 16724 9336 40868 9364
rect 16724 9324 16730 9336
rect 40862 9324 40868 9336
rect 40920 9324 40926 9376
rect 47578 9324 47584 9376
rect 47636 9364 47642 9376
rect 79502 9364 79508 9376
rect 47636 9336 79508 9364
rect 47636 9324 47642 9336
rect 79502 9324 79508 9336
rect 79560 9324 79566 9376
rect 83458 9324 83464 9376
rect 83516 9364 83522 9376
rect 91278 9364 91284 9376
rect 83516 9336 91284 9364
rect 83516 9324 83522 9336
rect 91278 9324 91284 9336
rect 91336 9324 91342 9376
rect 1104 9274 98808 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 50326 9274
rect 50378 9222 50390 9274
rect 50442 9222 50454 9274
rect 50506 9222 50518 9274
rect 50570 9222 81046 9274
rect 81098 9222 81110 9274
rect 81162 9222 81174 9274
rect 81226 9222 81238 9274
rect 81290 9222 98808 9274
rect 1104 9200 98808 9222
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 39666 9160 39672 9172
rect 3292 9132 39672 9160
rect 3292 9120 3298 9132
rect 39666 9120 39672 9132
rect 39724 9120 39730 9172
rect 49050 9120 49056 9172
rect 49108 9160 49114 9172
rect 91462 9160 91468 9172
rect 49108 9132 91468 9160
rect 49108 9120 49114 9132
rect 91462 9120 91468 9132
rect 91520 9120 91526 9172
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 53190 9092 53196 9104
rect 9824 9064 53196 9092
rect 9824 9052 9830 9064
rect 53190 9052 53196 9064
rect 53248 9052 53254 9104
rect 56042 9052 56048 9104
rect 56100 9092 56106 9104
rect 97442 9092 97448 9104
rect 56100 9064 97448 9092
rect 56100 9052 56106 9064
rect 97442 9052 97448 9064
rect 97500 9052 97506 9104
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 40770 9024 40776 9036
rect 4028 8996 40776 9024
rect 4028 8984 4034 8996
rect 40770 8984 40776 8996
rect 40828 8984 40834 9036
rect 49602 8984 49608 9036
rect 49660 9024 49666 9036
rect 96890 9024 96896 9036
rect 49660 8996 96896 9024
rect 49660 8984 49666 8996
rect 96890 8984 96896 8996
rect 96948 8984 96954 9036
rect 25406 8916 25412 8968
rect 25464 8956 25470 8968
rect 96062 8956 96068 8968
rect 25464 8928 96068 8956
rect 25464 8916 25470 8928
rect 96062 8916 96068 8928
rect 96120 8916 96126 8968
rect 1104 8730 98808 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 65686 8730
rect 65738 8678 65750 8730
rect 65802 8678 65814 8730
rect 65866 8678 65878 8730
rect 65930 8678 96406 8730
rect 96458 8678 96470 8730
rect 96522 8678 96534 8730
rect 96586 8678 96598 8730
rect 96650 8678 98808 8730
rect 1104 8656 98808 8678
rect 4798 8616 4804 8628
rect 4759 8588 4804 8616
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 12342 8616 12348 8628
rect 11756 8588 12348 8616
rect 11756 8576 11762 8588
rect 12342 8576 12348 8588
rect 12400 8616 12406 8628
rect 12400 8588 26234 8616
rect 12400 8576 12406 8588
rect 13909 8551 13967 8557
rect 13909 8517 13921 8551
rect 13955 8548 13967 8551
rect 16761 8551 16819 8557
rect 16761 8548 16773 8551
rect 13955 8520 16773 8548
rect 13955 8517 13967 8520
rect 13909 8511 13967 8517
rect 16761 8517 16773 8520
rect 16807 8517 16819 8551
rect 26206 8548 26234 8588
rect 60182 8548 60188 8560
rect 26206 8520 60188 8548
rect 16761 8511 16819 8517
rect 60182 8508 60188 8520
rect 60240 8508 60246 8560
rect 32858 8480 32864 8492
rect 5092 8452 32864 8480
rect 5092 8421 5120 8452
rect 32858 8440 32864 8452
rect 32916 8440 32922 8492
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8381 5135 8415
rect 75086 8412 75092 8424
rect 5077 8375 5135 8381
rect 12406 8384 75092 8412
rect 4062 8304 4068 8356
rect 4120 8344 4126 8356
rect 4433 8347 4491 8353
rect 4433 8344 4445 8347
rect 4120 8316 4445 8344
rect 4120 8304 4126 8316
rect 4433 8313 4445 8316
rect 4479 8344 4491 8347
rect 4908 8344 4936 8375
rect 12406 8344 12434 8384
rect 75086 8372 75092 8384
rect 75144 8372 75150 8424
rect 4479 8316 12434 8344
rect 16761 8347 16819 8353
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 16761 8313 16773 8347
rect 16807 8344 16819 8347
rect 50706 8344 50712 8356
rect 16807 8316 50712 8344
rect 16807 8313 16819 8316
rect 16761 8307 16819 8313
rect 50706 8304 50712 8316
rect 50764 8304 50770 8356
rect 63770 8304 63776 8356
rect 63828 8344 63834 8356
rect 67082 8344 67088 8356
rect 63828 8316 67088 8344
rect 63828 8304 63834 8316
rect 67082 8304 67088 8316
rect 67140 8304 67146 8356
rect 20622 8236 20628 8288
rect 20680 8276 20686 8288
rect 22922 8276 22928 8288
rect 20680 8248 22928 8276
rect 20680 8236 20686 8248
rect 22922 8236 22928 8248
rect 22980 8236 22986 8288
rect 23842 8236 23848 8288
rect 23900 8276 23906 8288
rect 25498 8276 25504 8288
rect 23900 8248 25504 8276
rect 23900 8236 23906 8248
rect 25498 8236 25504 8248
rect 25556 8236 25562 8288
rect 1104 8186 98808 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 50326 8186
rect 50378 8134 50390 8186
rect 50442 8134 50454 8186
rect 50506 8134 50518 8186
rect 50570 8134 81046 8186
rect 81098 8134 81110 8186
rect 81162 8134 81174 8186
rect 81226 8134 81238 8186
rect 81290 8134 98808 8186
rect 1104 8112 98808 8134
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 22830 8072 22836 8084
rect 18932 8044 22836 8072
rect 18932 8032 18938 8044
rect 22830 8032 22836 8044
rect 22888 8032 22894 8084
rect 28902 8032 28908 8084
rect 28960 8072 28966 8084
rect 74810 8072 74816 8084
rect 28960 8044 74816 8072
rect 28960 8032 28966 8044
rect 74810 8032 74816 8044
rect 74868 8032 74874 8084
rect 96798 8072 96804 8084
rect 94516 8044 96804 8072
rect 21450 7964 21456 8016
rect 21508 8004 21514 8016
rect 22094 8004 22100 8016
rect 21508 7976 22100 8004
rect 21508 7964 21514 7976
rect 22094 7964 22100 7976
rect 22152 7964 22158 8016
rect 64414 8004 64420 8016
rect 64327 7976 64420 8004
rect 64414 7964 64420 7976
rect 64472 8004 64478 8016
rect 79134 8004 79140 8016
rect 64472 7976 79140 8004
rect 64472 7964 64478 7976
rect 79134 7964 79140 7976
rect 79192 7964 79198 8016
rect 94516 8004 94544 8044
rect 96798 8032 96804 8044
rect 96856 8032 96862 8084
rect 94241 7976 94544 8004
rect 93854 7936 93860 7948
rect 93815 7908 93860 7936
rect 93854 7896 93860 7908
rect 93912 7896 93918 7948
rect 94241 7945 94269 7976
rect 94133 7939 94191 7945
rect 94133 7936 94145 7939
rect 93964 7908 94145 7936
rect 50982 7828 50988 7880
rect 51040 7868 51046 7880
rect 61378 7868 61384 7880
rect 51040 7840 61384 7868
rect 51040 7828 51046 7840
rect 61378 7828 61384 7840
rect 61436 7828 61442 7880
rect 62758 7868 62764 7880
rect 62719 7840 62764 7868
rect 62758 7828 62764 7840
rect 62816 7828 62822 7880
rect 63037 7871 63095 7877
rect 63037 7837 63049 7871
rect 63083 7868 63095 7871
rect 79226 7868 79232 7880
rect 63083 7840 79232 7868
rect 63083 7837 63095 7840
rect 63037 7831 63095 7837
rect 79226 7828 79232 7840
rect 79284 7828 79290 7880
rect 79686 7828 79692 7880
rect 79744 7868 79750 7880
rect 93964 7868 93992 7908
rect 94133 7905 94145 7908
rect 94179 7905 94191 7939
rect 94133 7899 94191 7905
rect 94226 7939 94284 7945
rect 94226 7905 94238 7939
rect 94272 7905 94284 7939
rect 94406 7936 94412 7948
rect 94367 7908 94412 7936
rect 94226 7899 94284 7905
rect 94406 7896 94412 7908
rect 94464 7896 94470 7948
rect 79744 7840 93992 7868
rect 94041 7871 94099 7877
rect 79744 7828 79750 7840
rect 94041 7837 94053 7871
rect 94087 7837 94099 7871
rect 94041 7831 94099 7837
rect 2958 7760 2964 7812
rect 3016 7800 3022 7812
rect 3016 7772 12434 7800
rect 3016 7760 3022 7772
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 9122 7732 9128 7744
rect 8812 7704 9128 7732
rect 8812 7692 8818 7704
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 12406 7732 12434 7772
rect 24486 7760 24492 7812
rect 24544 7800 24550 7812
rect 31110 7800 31116 7812
rect 24544 7772 31116 7800
rect 24544 7760 24550 7772
rect 31110 7760 31116 7772
rect 31168 7760 31174 7812
rect 45094 7760 45100 7812
rect 45152 7800 45158 7812
rect 59354 7800 59360 7812
rect 45152 7772 59360 7800
rect 45152 7760 45158 7772
rect 59354 7760 59360 7772
rect 59412 7760 59418 7812
rect 64064 7772 70394 7800
rect 29914 7732 29920 7744
rect 12406 7704 29920 7732
rect 29914 7692 29920 7704
rect 29972 7692 29978 7744
rect 39758 7692 39764 7744
rect 39816 7732 39822 7744
rect 64064 7732 64092 7772
rect 39816 7704 64092 7732
rect 70366 7732 70394 7772
rect 78490 7760 78496 7812
rect 78548 7800 78554 7812
rect 93673 7803 93731 7809
rect 93673 7800 93685 7803
rect 78548 7772 93685 7800
rect 78548 7760 78554 7772
rect 93673 7769 93685 7772
rect 93719 7769 93731 7803
rect 94056 7800 94084 7831
rect 93673 7763 93731 7769
rect 93964 7772 94084 7800
rect 93489 7735 93547 7741
rect 93489 7732 93501 7735
rect 70366 7704 93501 7732
rect 39816 7692 39822 7704
rect 93489 7701 93501 7704
rect 93535 7732 93547 7735
rect 93964 7732 93992 7772
rect 93535 7704 93992 7732
rect 93535 7701 93547 7704
rect 93489 7695 93547 7701
rect 94406 7692 94412 7744
rect 94464 7732 94470 7744
rect 94516 7741 94544 7976
rect 94501 7735 94559 7741
rect 94501 7732 94513 7735
rect 94464 7704 94513 7732
rect 94464 7692 94470 7704
rect 94501 7701 94513 7704
rect 94547 7701 94559 7735
rect 94501 7695 94559 7701
rect 1104 7642 98808 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 65686 7642
rect 65738 7590 65750 7642
rect 65802 7590 65814 7642
rect 65866 7590 65878 7642
rect 65930 7590 96406 7642
rect 96458 7590 96470 7642
rect 96522 7590 96534 7642
rect 96586 7590 96598 7642
rect 96650 7590 98808 7642
rect 1104 7568 98808 7590
rect 16206 7488 16212 7540
rect 16264 7528 16270 7540
rect 64414 7528 64420 7540
rect 16264 7500 64420 7528
rect 16264 7488 16270 7500
rect 64414 7488 64420 7500
rect 64472 7488 64478 7540
rect 41046 7420 41052 7472
rect 41104 7460 41110 7472
rect 43717 7463 43775 7469
rect 43717 7460 43729 7463
rect 41104 7432 43729 7460
rect 41104 7420 41110 7432
rect 43717 7429 43729 7432
rect 43763 7429 43775 7463
rect 43717 7423 43775 7429
rect 17862 7352 17868 7404
rect 17920 7392 17926 7404
rect 17920 7364 45554 7392
rect 17920 7352 17926 7364
rect 13081 7327 13139 7333
rect 13081 7293 13093 7327
rect 13127 7324 13139 7327
rect 45005 7327 45063 7333
rect 45005 7324 45017 7327
rect 13127 7296 22094 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 22066 7256 22094 7296
rect 43456 7296 45017 7324
rect 43346 7256 43352 7268
rect 22066 7228 43352 7256
rect 43346 7216 43352 7228
rect 43404 7216 43410 7268
rect 13354 7148 13360 7200
rect 13412 7188 13418 7200
rect 16390 7188 16396 7200
rect 13412 7160 16396 7188
rect 13412 7148 13418 7160
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 29638 7148 29644 7200
rect 29696 7188 29702 7200
rect 43456 7197 43484 7296
rect 45005 7293 45017 7296
rect 45051 7293 45063 7327
rect 45005 7287 45063 7293
rect 45281 7327 45339 7333
rect 45281 7293 45293 7327
rect 45327 7293 45339 7327
rect 45281 7287 45339 7293
rect 43441 7191 43499 7197
rect 43441 7188 43453 7191
rect 29696 7160 43453 7188
rect 29696 7148 29702 7160
rect 43441 7157 43453 7160
rect 43487 7157 43499 7191
rect 43441 7151 43499 7157
rect 44082 7148 44088 7200
rect 44140 7188 44146 7200
rect 45296 7188 45324 7287
rect 45526 7256 45554 7364
rect 57348 7364 60734 7392
rect 57348 7333 57376 7364
rect 57333 7327 57391 7333
rect 57333 7293 57345 7327
rect 57379 7293 57391 7327
rect 57333 7287 57391 7293
rect 57425 7327 57483 7333
rect 57425 7293 57437 7327
rect 57471 7293 57483 7327
rect 60706 7324 60734 7364
rect 84746 7324 84752 7336
rect 60706 7296 84752 7324
rect 57425 7287 57483 7293
rect 57440 7256 57468 7287
rect 84746 7284 84752 7296
rect 84804 7284 84810 7336
rect 85574 7284 85580 7336
rect 85632 7324 85638 7336
rect 90913 7327 90971 7333
rect 90913 7324 90925 7327
rect 85632 7296 90925 7324
rect 85632 7284 85638 7296
rect 90913 7293 90925 7296
rect 90959 7293 90971 7327
rect 90913 7287 90971 7293
rect 45526 7228 57468 7256
rect 44140 7160 45324 7188
rect 57793 7191 57851 7197
rect 44140 7148 44146 7160
rect 57793 7157 57805 7191
rect 57839 7188 57851 7191
rect 87966 7188 87972 7200
rect 57839 7160 87972 7188
rect 57839 7157 57851 7160
rect 57793 7151 57851 7157
rect 87966 7148 87972 7160
rect 88024 7148 88030 7200
rect 1104 7098 98808 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 50326 7098
rect 50378 7046 50390 7098
rect 50442 7046 50454 7098
rect 50506 7046 50518 7098
rect 50570 7046 81046 7098
rect 81098 7046 81110 7098
rect 81162 7046 81174 7098
rect 81226 7046 81238 7098
rect 81290 7046 98808 7098
rect 1104 7024 98808 7046
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 94406 6984 94412 6996
rect 2648 6956 94412 6984
rect 2648 6944 2654 6956
rect 94406 6944 94412 6956
rect 94464 6944 94470 6996
rect 13906 6876 13912 6928
rect 13964 6916 13970 6928
rect 16114 6916 16120 6928
rect 13964 6888 16120 6916
rect 13964 6876 13970 6888
rect 16114 6876 16120 6888
rect 16172 6876 16178 6928
rect 59648 6888 60044 6916
rect 50525 6851 50583 6857
rect 45526 6820 50384 6848
rect 45186 6740 45192 6792
rect 45244 6780 45250 6792
rect 45526 6780 45554 6820
rect 50249 6783 50307 6789
rect 50249 6780 50261 6783
rect 45244 6752 45554 6780
rect 49068 6752 50261 6780
rect 45244 6740 45250 6752
rect 38746 6672 38752 6724
rect 38804 6712 38810 6724
rect 48961 6715 49019 6721
rect 48961 6712 48973 6715
rect 38804 6684 48973 6712
rect 38804 6672 38810 6684
rect 48961 6681 48973 6684
rect 49007 6681 49019 6715
rect 48961 6675 49019 6681
rect 48682 6644 48688 6656
rect 48643 6616 48688 6644
rect 48682 6604 48688 6616
rect 48740 6644 48746 6656
rect 49068 6644 49096 6752
rect 50249 6749 50261 6752
rect 50295 6749 50307 6783
rect 50356 6780 50384 6820
rect 50525 6817 50537 6851
rect 50571 6848 50583 6851
rect 59648 6848 59676 6888
rect 50571 6820 59676 6848
rect 50571 6817 50583 6820
rect 50525 6811 50583 6817
rect 59722 6808 59728 6860
rect 59780 6848 59786 6860
rect 59909 6851 59967 6857
rect 59909 6848 59921 6851
rect 59780 6820 59921 6848
rect 59780 6808 59786 6820
rect 59909 6817 59921 6820
rect 59955 6817 59967 6851
rect 60016 6848 60044 6888
rect 62758 6848 62764 6860
rect 60016 6820 62764 6848
rect 59909 6811 59967 6817
rect 62758 6808 62764 6820
rect 62816 6808 62822 6860
rect 97537 6851 97595 6857
rect 97537 6817 97549 6851
rect 97583 6848 97595 6851
rect 98270 6848 98276 6860
rect 97583 6820 98276 6848
rect 97583 6817 97595 6820
rect 97537 6811 97595 6817
rect 98270 6808 98276 6820
rect 98328 6808 98334 6860
rect 60277 6783 60335 6789
rect 60277 6780 60289 6783
rect 50356 6752 60289 6780
rect 50249 6743 50307 6749
rect 60277 6749 60289 6752
rect 60323 6749 60335 6783
rect 60277 6743 60335 6749
rect 53558 6672 53564 6724
rect 53616 6712 53622 6724
rect 60047 6715 60105 6721
rect 60047 6712 60059 6715
rect 53616 6684 60059 6712
rect 53616 6672 53622 6684
rect 60047 6681 60059 6684
rect 60093 6681 60105 6715
rect 60182 6712 60188 6724
rect 60143 6684 60188 6712
rect 60047 6675 60105 6681
rect 60182 6672 60188 6684
rect 60240 6672 60246 6724
rect 84654 6712 84660 6724
rect 60706 6684 84660 6712
rect 56962 6644 56968 6656
rect 48740 6616 49096 6644
rect 56923 6616 56968 6644
rect 48740 6604 48746 6616
rect 56962 6604 56968 6616
rect 57020 6604 57026 6656
rect 59722 6644 59728 6656
rect 59683 6616 59728 6644
rect 59722 6604 59728 6616
rect 59780 6604 59786 6656
rect 60553 6647 60611 6653
rect 60553 6613 60565 6647
rect 60599 6644 60611 6647
rect 60706 6644 60734 6684
rect 84654 6672 84660 6684
rect 84712 6672 84718 6724
rect 60599 6616 60734 6644
rect 60599 6613 60611 6616
rect 60553 6607 60611 6613
rect 78030 6604 78036 6656
rect 78088 6644 78094 6656
rect 81621 6647 81679 6653
rect 81621 6644 81633 6647
rect 78088 6616 81633 6644
rect 78088 6604 78094 6616
rect 81621 6613 81633 6616
rect 81667 6613 81679 6647
rect 81621 6607 81679 6613
rect 96893 6647 96951 6653
rect 96893 6613 96905 6647
rect 96939 6644 96951 6647
rect 97534 6644 97540 6656
rect 96939 6616 97540 6644
rect 96939 6613 96951 6616
rect 96893 6607 96951 6613
rect 97534 6604 97540 6616
rect 97592 6604 97598 6656
rect 1104 6554 98808 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 65686 6554
rect 65738 6502 65750 6554
rect 65802 6502 65814 6554
rect 65866 6502 65878 6554
rect 65930 6502 96406 6554
rect 96458 6502 96470 6554
rect 96522 6502 96534 6554
rect 96586 6502 96598 6554
rect 96650 6502 98808 6554
rect 1104 6480 98808 6502
rect 14182 6400 14188 6452
rect 14240 6440 14246 6452
rect 48682 6440 48688 6452
rect 14240 6412 48688 6440
rect 14240 6400 14246 6412
rect 48682 6400 48688 6412
rect 48740 6400 48746 6452
rect 53834 6400 53840 6452
rect 53892 6440 53898 6452
rect 78030 6440 78036 6452
rect 53892 6412 78036 6440
rect 53892 6400 53898 6412
rect 78030 6400 78036 6412
rect 78088 6400 78094 6452
rect 92106 6440 92112 6452
rect 92067 6412 92112 6440
rect 92106 6400 92112 6412
rect 92164 6400 92170 6452
rect 13998 6264 14004 6316
rect 14056 6304 14062 6316
rect 38746 6304 38752 6316
rect 14056 6276 38752 6304
rect 14056 6264 14062 6276
rect 38746 6264 38752 6276
rect 38804 6264 38810 6316
rect 92124 6304 92152 6400
rect 93673 6307 93731 6313
rect 93673 6304 93685 6307
rect 92124 6276 93685 6304
rect 93673 6273 93685 6276
rect 93719 6273 93731 6307
rect 93673 6267 93731 6273
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6236 14703 6239
rect 52454 6236 52460 6248
rect 14691 6208 52460 6236
rect 14691 6205 14703 6208
rect 14645 6199 14703 6205
rect 52454 6196 52460 6208
rect 52512 6196 52518 6248
rect 61930 6196 61936 6248
rect 61988 6236 61994 6248
rect 71038 6236 71044 6248
rect 61988 6208 71044 6236
rect 61988 6196 61994 6208
rect 71038 6196 71044 6208
rect 71096 6196 71102 6248
rect 90450 6196 90456 6248
rect 90508 6236 90514 6248
rect 93949 6239 94007 6245
rect 93949 6236 93961 6239
rect 90508 6208 93961 6236
rect 90508 6196 90514 6208
rect 93949 6205 93961 6208
rect 93995 6205 94007 6239
rect 93949 6199 94007 6205
rect 96985 6239 97043 6245
rect 96985 6205 96997 6239
rect 97031 6205 97043 6239
rect 97626 6236 97632 6248
rect 97587 6208 97632 6236
rect 96985 6199 97043 6205
rect 8386 6128 8392 6180
rect 8444 6168 8450 6180
rect 53558 6168 53564 6180
rect 8444 6140 53564 6168
rect 8444 6128 8450 6140
rect 53558 6128 53564 6140
rect 53616 6128 53622 6180
rect 59630 6128 59636 6180
rect 59688 6168 59694 6180
rect 73522 6168 73528 6180
rect 59688 6140 73528 6168
rect 59688 6128 59694 6140
rect 73522 6128 73528 6140
rect 73580 6128 73586 6180
rect 92293 6171 92351 6177
rect 92293 6168 92305 6171
rect 84166 6140 92305 6168
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 21726 6100 21732 6112
rect 20772 6072 21732 6100
rect 20772 6060 20778 6072
rect 21726 6060 21732 6072
rect 21784 6100 21790 6112
rect 59722 6100 59728 6112
rect 21784 6072 59728 6100
rect 21784 6060 21790 6072
rect 59722 6060 59728 6072
rect 59780 6060 59786 6112
rect 72694 6060 72700 6112
rect 72752 6100 72758 6112
rect 84166 6100 84194 6140
rect 92293 6137 92305 6140
rect 92339 6137 92351 6171
rect 97000 6168 97028 6199
rect 97626 6196 97632 6208
rect 97684 6196 97690 6248
rect 98822 6168 98828 6180
rect 97000 6140 98828 6168
rect 92293 6131 92351 6137
rect 98822 6128 98828 6140
rect 98880 6128 98886 6180
rect 72752 6072 84194 6100
rect 72752 6060 72758 6072
rect 1104 6010 98808 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 50326 6010
rect 50378 5958 50390 6010
rect 50442 5958 50454 6010
rect 50506 5958 50518 6010
rect 50570 5958 81046 6010
rect 81098 5958 81110 6010
rect 81162 5958 81174 6010
rect 81226 5958 81238 6010
rect 81290 5958 98808 6010
rect 1104 5936 98808 5958
rect 50154 5856 50160 5908
rect 50212 5896 50218 5908
rect 50341 5899 50399 5905
rect 50341 5896 50353 5899
rect 50212 5868 50353 5896
rect 50212 5856 50218 5868
rect 50341 5865 50353 5868
rect 50387 5865 50399 5899
rect 50341 5859 50399 5865
rect 82446 5856 82452 5908
rect 82504 5896 82510 5908
rect 84930 5896 84936 5908
rect 82504 5868 84936 5896
rect 82504 5856 82510 5868
rect 84930 5856 84936 5868
rect 84988 5856 84994 5908
rect 85206 5896 85212 5908
rect 85167 5868 85212 5896
rect 85206 5856 85212 5868
rect 85264 5856 85270 5908
rect 50062 5788 50068 5840
rect 50120 5828 50126 5840
rect 50249 5831 50307 5837
rect 50249 5828 50261 5831
rect 50120 5800 50261 5828
rect 50120 5788 50126 5800
rect 50249 5797 50261 5800
rect 50295 5797 50307 5831
rect 50249 5791 50307 5797
rect 88978 5788 88984 5840
rect 89036 5828 89042 5840
rect 91189 5831 91247 5837
rect 91189 5828 91201 5831
rect 89036 5800 91201 5828
rect 89036 5788 89042 5800
rect 91189 5797 91201 5800
rect 91235 5797 91247 5831
rect 91189 5791 91247 5797
rect 2682 5760 2688 5772
rect 2643 5732 2688 5760
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 69658 5720 69664 5772
rect 69716 5760 69722 5772
rect 84102 5760 84108 5772
rect 69716 5732 83964 5760
rect 84063 5732 84108 5760
rect 69716 5720 69722 5732
rect 80238 5652 80244 5704
rect 80296 5692 80302 5704
rect 83829 5695 83887 5701
rect 83829 5692 83841 5695
rect 80296 5664 83841 5692
rect 80296 5652 80302 5664
rect 83829 5661 83841 5664
rect 83875 5661 83887 5695
rect 83936 5692 83964 5732
rect 84102 5720 84108 5732
rect 84160 5720 84166 5772
rect 91646 5760 91652 5772
rect 91607 5732 91652 5760
rect 91646 5720 91652 5732
rect 91704 5720 91710 5772
rect 91833 5763 91891 5769
rect 91833 5729 91845 5763
rect 91879 5760 91891 5763
rect 91922 5760 91928 5772
rect 91879 5732 91928 5760
rect 91879 5729 91891 5732
rect 91833 5723 91891 5729
rect 91922 5720 91928 5732
rect 91980 5720 91986 5772
rect 92017 5763 92075 5769
rect 92017 5729 92029 5763
rect 92063 5729 92075 5763
rect 92017 5723 92075 5729
rect 96249 5763 96307 5769
rect 96249 5729 96261 5763
rect 96295 5729 96307 5763
rect 96249 5723 96307 5729
rect 96893 5763 96951 5769
rect 96893 5729 96905 5763
rect 96939 5760 96951 5763
rect 96982 5760 96988 5772
rect 96939 5732 96988 5760
rect 96939 5729 96951 5732
rect 96893 5723 96951 5729
rect 92032 5692 92060 5723
rect 83936 5664 92060 5692
rect 96264 5692 96292 5723
rect 96982 5720 96988 5732
rect 97040 5720 97046 5772
rect 97537 5763 97595 5769
rect 97537 5729 97549 5763
rect 97583 5760 97595 5763
rect 99006 5760 99012 5772
rect 97583 5732 99012 5760
rect 97583 5729 97595 5732
rect 97537 5723 97595 5729
rect 99006 5720 99012 5732
rect 99064 5720 99070 5772
rect 99466 5692 99472 5704
rect 96264 5664 99472 5692
rect 83829 5655 83887 5661
rect 13722 5516 13728 5568
rect 13780 5556 13786 5568
rect 14274 5556 14280 5568
rect 13780 5528 14280 5556
rect 13780 5516 13786 5528
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 83844 5556 83872 5655
rect 99466 5652 99472 5664
rect 99524 5652 99530 5704
rect 90450 5556 90456 5568
rect 83844 5528 90456 5556
rect 90450 5516 90456 5528
rect 90508 5516 90514 5568
rect 1104 5466 98808 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 65686 5466
rect 65738 5414 65750 5466
rect 65802 5414 65814 5466
rect 65866 5414 65878 5466
rect 65930 5414 96406 5466
rect 96458 5414 96470 5466
rect 96522 5414 96534 5466
rect 96586 5414 96598 5466
rect 96650 5414 98808 5466
rect 1104 5392 98808 5414
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 68462 5352 68468 5364
rect 6696 5324 68468 5352
rect 6696 5312 6702 5324
rect 68462 5312 68468 5324
rect 68520 5312 68526 5364
rect 82262 5312 82268 5364
rect 82320 5352 82326 5364
rect 85022 5352 85028 5364
rect 82320 5324 85028 5352
rect 82320 5312 82326 5324
rect 85022 5312 85028 5324
rect 85080 5312 85086 5364
rect 16298 5244 16304 5296
rect 16356 5284 16362 5296
rect 46290 5284 46296 5296
rect 16356 5256 46296 5284
rect 16356 5244 16362 5256
rect 46290 5244 46296 5256
rect 46348 5244 46354 5296
rect 67358 5244 67364 5296
rect 67416 5284 67422 5296
rect 80606 5284 80612 5296
rect 67416 5256 80612 5284
rect 67416 5244 67422 5256
rect 80606 5244 80612 5256
rect 80664 5244 80670 5296
rect 3510 5176 3516 5228
rect 3568 5216 3574 5228
rect 3568 5188 4108 5216
rect 3568 5176 3574 5188
rect 1854 5108 1860 5160
rect 1912 5148 1918 5160
rect 4080 5157 4108 5188
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 16942 5216 16948 5228
rect 7524 5188 16948 5216
rect 7524 5176 7530 5188
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 17126 5176 17132 5228
rect 17184 5216 17190 5228
rect 35434 5216 35440 5228
rect 17184 5188 35440 5216
rect 17184 5176 17190 5188
rect 35434 5176 35440 5188
rect 35492 5176 35498 5228
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 1912 5120 2513 5148
rect 1912 5108 1918 5120
rect 2501 5117 2513 5120
rect 2547 5117 2559 5151
rect 4065 5151 4123 5157
rect 2501 5111 2559 5117
rect 2746 5120 4016 5148
rect 1673 5083 1731 5089
rect 1673 5049 1685 5083
rect 1719 5080 1731 5083
rect 1949 5083 2007 5089
rect 1949 5080 1961 5083
rect 1719 5052 1961 5080
rect 1719 5049 1731 5052
rect 1673 5043 1731 5049
rect 1949 5049 1961 5052
rect 1995 5080 2007 5083
rect 2746 5080 2774 5120
rect 3326 5080 3332 5092
rect 1995 5052 2774 5080
rect 3287 5052 3332 5080
rect 1995 5049 2007 5052
rect 1949 5043 2007 5049
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3513 5083 3571 5089
rect 3513 5049 3525 5083
rect 3559 5080 3571 5083
rect 3602 5080 3608 5092
rect 3559 5052 3608 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 474 4972 480 5024
rect 532 5012 538 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 532 4984 1869 5012
rect 532 4972 538 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 1857 4975 1915 4981
rect 3237 5015 3295 5021
rect 3237 4981 3249 5015
rect 3283 5012 3295 5015
rect 3528 5012 3556 5043
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 3988 5080 4016 5120
rect 4065 5117 4077 5151
rect 4111 5117 4123 5151
rect 4065 5111 4123 5117
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 4798 5148 4804 5160
rect 4755 5120 4804 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 7006 5148 7012 5160
rect 6967 5120 7012 5148
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 10594 5148 10600 5160
rect 10555 5120 10600 5148
rect 10594 5108 10600 5120
rect 10652 5108 10658 5160
rect 11882 5108 11888 5160
rect 11940 5148 11946 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11940 5120 12081 5148
rect 11940 5108 11946 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 13078 5148 13084 5160
rect 13039 5120 13084 5148
rect 12069 5111 12127 5117
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 14274 5148 14280 5160
rect 14235 5120 14280 5148
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 15470 5148 15476 5160
rect 15431 5120 15476 5148
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 16850 5108 16856 5160
rect 16908 5148 16914 5160
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 16908 5120 17325 5148
rect 16908 5108 16914 5120
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 18598 5148 18604 5160
rect 18559 5120 18604 5148
rect 17313 5111 17371 5117
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 24394 5148 24400 5160
rect 24355 5120 24400 5148
rect 24394 5108 24400 5120
rect 24452 5108 24458 5160
rect 80514 5148 80520 5160
rect 80475 5120 80520 5148
rect 80514 5108 80520 5120
rect 80572 5108 80578 5160
rect 96246 5108 96252 5160
rect 96304 5148 96310 5160
rect 96433 5151 96491 5157
rect 96433 5148 96445 5151
rect 96304 5120 96445 5148
rect 96304 5108 96310 5120
rect 96433 5117 96445 5120
rect 96479 5117 96491 5151
rect 96433 5111 96491 5117
rect 97169 5151 97227 5157
rect 97169 5117 97181 5151
rect 97215 5117 97227 5151
rect 97810 5148 97816 5160
rect 97771 5120 97816 5148
rect 97169 5111 97227 5117
rect 43438 5080 43444 5092
rect 3988 5052 43444 5080
rect 43438 5040 43444 5052
rect 43496 5040 43502 5092
rect 56962 5040 56968 5092
rect 57020 5080 57026 5092
rect 73706 5080 73712 5092
rect 57020 5052 73712 5080
rect 57020 5040 57026 5052
rect 73706 5040 73712 5052
rect 73764 5040 73770 5092
rect 97184 5080 97212 5111
rect 97810 5108 97816 5120
rect 97868 5108 97874 5160
rect 98454 5080 98460 5092
rect 97184 5052 98460 5080
rect 98454 5040 98460 5052
rect 98512 5040 98518 5092
rect 3283 4984 3556 5012
rect 3283 4981 3295 4984
rect 3237 4975 3295 4981
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 17218 5012 17224 5024
rect 5224 4984 17224 5012
rect 5224 4972 5230 4984
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 24578 5012 24584 5024
rect 24539 4984 24584 5012
rect 24578 4972 24584 4984
rect 24636 4972 24642 5024
rect 52454 4972 52460 5024
rect 52512 5012 52518 5024
rect 86954 5012 86960 5024
rect 52512 4984 86960 5012
rect 52512 4972 52518 4984
rect 86954 4972 86960 4984
rect 87012 4972 87018 5024
rect 1104 4922 98808 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 50326 4922
rect 50378 4870 50390 4922
rect 50442 4870 50454 4922
rect 50506 4870 50518 4922
rect 50570 4870 81046 4922
rect 81098 4870 81110 4922
rect 81162 4870 81174 4922
rect 81226 4870 81238 4922
rect 81290 4870 98808 4922
rect 1104 4848 98808 4870
rect 15194 4808 15200 4820
rect 4448 4780 12434 4808
rect 15155 4780 15200 4808
rect 1673 4743 1731 4749
rect 1673 4709 1685 4743
rect 1719 4740 1731 4743
rect 1762 4740 1768 4752
rect 1719 4712 1768 4740
rect 1719 4709 1731 4712
rect 1673 4703 1731 4709
rect 1762 4700 1768 4712
rect 1820 4700 1826 4752
rect 4448 4749 4476 4780
rect 4157 4743 4215 4749
rect 4157 4709 4169 4743
rect 4203 4740 4215 4743
rect 4433 4743 4491 4749
rect 4433 4740 4445 4743
rect 4203 4712 4445 4740
rect 4203 4709 4215 4712
rect 4157 4703 4215 4709
rect 4433 4709 4445 4712
rect 4479 4709 4491 4743
rect 4433 4703 4491 4709
rect 4893 4743 4951 4749
rect 4893 4709 4905 4743
rect 4939 4740 4951 4743
rect 5166 4740 5172 4752
rect 4939 4712 5172 4740
rect 4939 4709 4951 4712
rect 4893 4703 4951 4709
rect 5166 4700 5172 4712
rect 5224 4700 5230 4752
rect 5629 4743 5687 4749
rect 5629 4709 5641 4743
rect 5675 4740 5687 4743
rect 5902 4740 5908 4752
rect 5675 4712 5908 4740
rect 5675 4709 5687 4712
rect 5629 4703 5687 4709
rect 5902 4700 5908 4712
rect 5960 4700 5966 4752
rect 6365 4743 6423 4749
rect 6365 4709 6377 4743
rect 6411 4740 6423 4743
rect 6638 4740 6644 4752
rect 6411 4712 6644 4740
rect 6411 4709 6423 4712
rect 6365 4703 6423 4709
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 7466 4740 7472 4752
rect 7427 4712 7472 4740
rect 7466 4700 7472 4712
rect 7524 4700 7530 4752
rect 11146 4740 11152 4752
rect 11107 4712 11152 4740
rect 11146 4700 11152 4712
rect 11204 4700 11210 4752
rect 11330 4740 11336 4752
rect 11291 4712 11336 4740
rect 11330 4700 11336 4712
rect 11388 4700 11394 4752
rect 11790 4700 11796 4752
rect 11848 4740 11854 4752
rect 11885 4743 11943 4749
rect 11885 4740 11897 4743
rect 11848 4712 11897 4740
rect 11848 4700 11854 4712
rect 11885 4709 11897 4712
rect 11931 4709 11943 4743
rect 12406 4740 12434 4780
rect 15194 4768 15200 4780
rect 15252 4768 15258 4820
rect 17218 4768 17224 4820
rect 17276 4808 17282 4820
rect 32398 4808 32404 4820
rect 17276 4780 32404 4808
rect 17276 4768 17282 4780
rect 32398 4768 32404 4780
rect 32456 4768 32462 4820
rect 43346 4768 43352 4820
rect 43404 4808 43410 4820
rect 43404 4780 60734 4808
rect 43404 4768 43410 4780
rect 41138 4740 41144 4752
rect 12406 4712 41144 4740
rect 11885 4703 11943 4709
rect 41138 4700 41144 4712
rect 41196 4700 41202 4752
rect 60706 4740 60734 4780
rect 79318 4768 79324 4820
rect 79376 4808 79382 4820
rect 81526 4808 81532 4820
rect 79376 4780 81532 4808
rect 79376 4768 79382 4780
rect 81526 4768 81532 4780
rect 81584 4768 81590 4820
rect 82078 4768 82084 4820
rect 82136 4808 82142 4820
rect 84562 4808 84568 4820
rect 82136 4780 84568 4808
rect 82136 4768 82142 4780
rect 84562 4768 84568 4780
rect 84620 4768 84626 4820
rect 80146 4740 80152 4752
rect 60706 4712 80152 4740
rect 80146 4700 80152 4712
rect 80204 4700 80210 4752
rect 842 4632 848 4684
rect 900 4672 906 4684
rect 1397 4675 1455 4681
rect 1397 4672 1409 4675
rect 900 4644 1409 4672
rect 900 4632 906 4644
rect 1397 4641 1409 4644
rect 1443 4641 1455 4675
rect 2314 4672 2320 4684
rect 2275 4644 2320 4672
rect 1397 4635 1455 4641
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 8113 4675 8171 4681
rect 8113 4672 8125 4675
rect 7616 4644 8125 4672
rect 7616 4632 7622 4644
rect 8113 4641 8125 4644
rect 8159 4641 8171 4675
rect 10042 4672 10048 4684
rect 10003 4644 10048 4672
rect 8113 4635 8171 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 12526 4672 12532 4684
rect 12487 4644 12532 4672
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 13173 4675 13231 4681
rect 13173 4641 13185 4675
rect 13219 4641 13231 4675
rect 13173 4635 13231 4641
rect 14921 4675 14979 4681
rect 14921 4641 14933 4675
rect 14967 4672 14979 4675
rect 15105 4675 15163 4681
rect 15105 4672 15117 4675
rect 14967 4644 15117 4672
rect 14967 4641 14979 4644
rect 14921 4635 14979 4641
rect 15105 4641 15117 4644
rect 15151 4641 15163 4675
rect 15746 4672 15752 4684
rect 15707 4644 15752 4672
rect 15105 4635 15163 4641
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 2639 4576 2774 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 2746 4536 2774 4576
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5592 4576 5733 4604
rect 5592 4564 5598 4576
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6236 4576 6469 4604
rect 6236 4564 6242 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 13188 4604 13216 4635
rect 12492 4576 13216 4604
rect 15120 4604 15148 4635
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 16114 4632 16120 4684
rect 16172 4672 16178 4684
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 16172 4644 16405 4672
rect 16172 4632 16178 4644
rect 16393 4641 16405 4644
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 17126 4632 17132 4684
rect 17184 4672 17190 4684
rect 17221 4675 17279 4681
rect 17221 4672 17233 4675
rect 17184 4644 17233 4672
rect 17184 4632 17190 4644
rect 17221 4641 17233 4644
rect 17267 4641 17279 4675
rect 17221 4635 17279 4641
rect 17310 4632 17316 4684
rect 17368 4672 17374 4684
rect 17865 4675 17923 4681
rect 17865 4672 17877 4675
rect 17368 4644 17877 4672
rect 17368 4632 17374 4644
rect 17865 4641 17877 4644
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 17954 4632 17960 4684
rect 18012 4672 18018 4684
rect 18509 4675 18567 4681
rect 18509 4672 18521 4675
rect 18012 4644 18521 4672
rect 18012 4632 18018 4644
rect 18509 4641 18521 4644
rect 18555 4641 18567 4675
rect 18509 4635 18567 4641
rect 19426 4632 19432 4684
rect 19484 4672 19490 4684
rect 19981 4675 20039 4681
rect 19981 4672 19993 4675
rect 19484 4644 19993 4672
rect 19484 4632 19490 4644
rect 19981 4641 19993 4644
rect 20027 4641 20039 4675
rect 19981 4635 20039 4641
rect 20346 4632 20352 4684
rect 20404 4672 20410 4684
rect 20625 4675 20683 4681
rect 20625 4672 20637 4675
rect 20404 4644 20637 4672
rect 20404 4632 20410 4644
rect 20625 4641 20637 4644
rect 20671 4641 20683 4675
rect 20625 4635 20683 4641
rect 21082 4632 21088 4684
rect 21140 4672 21146 4684
rect 21269 4675 21327 4681
rect 21269 4672 21281 4675
rect 21140 4644 21281 4672
rect 21140 4632 21146 4644
rect 21269 4641 21281 4644
rect 21315 4641 21327 4675
rect 21269 4635 21327 4641
rect 25038 4632 25044 4684
rect 25096 4672 25102 4684
rect 25225 4675 25283 4681
rect 25225 4672 25237 4675
rect 25096 4644 25237 4672
rect 25096 4632 25102 4644
rect 25225 4641 25237 4644
rect 25271 4641 25283 4675
rect 25225 4635 25283 4641
rect 25682 4632 25688 4684
rect 25740 4672 25746 4684
rect 25869 4675 25927 4681
rect 25869 4672 25881 4675
rect 25740 4644 25881 4672
rect 25740 4632 25746 4644
rect 25869 4641 25881 4644
rect 25915 4641 25927 4675
rect 25869 4635 25927 4641
rect 26418 4632 26424 4684
rect 26476 4672 26482 4684
rect 26513 4675 26571 4681
rect 26513 4672 26525 4675
rect 26476 4644 26525 4672
rect 26476 4632 26482 4644
rect 26513 4641 26525 4644
rect 26559 4641 26571 4675
rect 26513 4635 26571 4641
rect 26878 4632 26884 4684
rect 26936 4672 26942 4684
rect 27157 4675 27215 4681
rect 27157 4672 27169 4675
rect 26936 4644 27169 4672
rect 26936 4632 26942 4644
rect 27157 4641 27169 4644
rect 27203 4641 27215 4675
rect 37274 4672 37280 4684
rect 37235 4644 37280 4672
rect 27157 4635 27215 4641
rect 37274 4632 37280 4644
rect 37332 4632 37338 4684
rect 39114 4672 39120 4684
rect 39075 4644 39120 4672
rect 39114 4632 39120 4644
rect 39172 4632 39178 4684
rect 39666 4632 39672 4684
rect 39724 4672 39730 4684
rect 39761 4675 39819 4681
rect 39761 4672 39773 4675
rect 39724 4644 39773 4672
rect 39724 4632 39730 4644
rect 39761 4641 39773 4644
rect 39807 4641 39819 4675
rect 39761 4635 39819 4641
rect 41693 4675 41751 4681
rect 41693 4641 41705 4675
rect 41739 4672 41751 4675
rect 44082 4672 44088 4684
rect 41739 4644 44088 4672
rect 41739 4641 41751 4644
rect 41693 4635 41751 4641
rect 44082 4632 44088 4644
rect 44140 4632 44146 4684
rect 44542 4672 44548 4684
rect 44503 4644 44548 4672
rect 44542 4632 44548 4644
rect 44600 4632 44606 4684
rect 45830 4632 45836 4684
rect 45888 4672 45894 4684
rect 46201 4675 46259 4681
rect 46201 4672 46213 4675
rect 45888 4644 46213 4672
rect 45888 4632 45894 4644
rect 46201 4641 46213 4644
rect 46247 4641 46259 4675
rect 47026 4672 47032 4684
rect 46987 4644 47032 4672
rect 46201 4635 46259 4641
rect 47026 4632 47032 4644
rect 47084 4632 47090 4684
rect 47578 4632 47584 4684
rect 47636 4672 47642 4684
rect 47673 4675 47731 4681
rect 47673 4672 47685 4675
rect 47636 4644 47685 4672
rect 47636 4632 47642 4644
rect 47673 4641 47685 4644
rect 47719 4641 47731 4675
rect 47673 4635 47731 4641
rect 48222 4632 48228 4684
rect 48280 4672 48286 4684
rect 48317 4675 48375 4681
rect 48317 4672 48329 4675
rect 48280 4644 48329 4672
rect 48280 4632 48286 4644
rect 48317 4641 48329 4644
rect 48363 4641 48375 4675
rect 52546 4672 52552 4684
rect 52507 4644 52552 4672
rect 48317 4635 48375 4641
rect 52546 4632 52552 4644
rect 52604 4632 52610 4684
rect 53098 4632 53104 4684
rect 53156 4672 53162 4684
rect 53193 4675 53251 4681
rect 53193 4672 53205 4675
rect 53156 4644 53205 4672
rect 53156 4632 53162 4644
rect 53193 4641 53205 4644
rect 53239 4641 53251 4675
rect 62850 4672 62856 4684
rect 62811 4644 62856 4672
rect 53193 4635 53251 4641
rect 62850 4632 62856 4644
rect 62908 4632 62914 4684
rect 73798 4672 73804 4684
rect 73759 4644 73804 4672
rect 73798 4632 73804 4644
rect 73856 4632 73862 4684
rect 78766 4672 78772 4684
rect 78727 4644 78772 4672
rect 78766 4632 78772 4644
rect 78824 4632 78830 4684
rect 79318 4632 79324 4684
rect 79376 4672 79382 4684
rect 79413 4675 79471 4681
rect 79413 4672 79425 4675
rect 79376 4644 79425 4672
rect 79376 4632 79382 4644
rect 79413 4641 79425 4644
rect 79459 4641 79471 4675
rect 80054 4672 80060 4684
rect 80015 4644 80060 4672
rect 79413 4635 79471 4641
rect 80054 4632 80060 4644
rect 80112 4632 80118 4684
rect 80790 4672 80796 4684
rect 80751 4644 80796 4672
rect 80790 4632 80796 4644
rect 80848 4632 80854 4684
rect 81434 4672 81440 4684
rect 81395 4644 81440 4672
rect 81434 4632 81440 4644
rect 81492 4632 81498 4684
rect 82906 4672 82912 4684
rect 82867 4644 82912 4672
rect 82906 4632 82912 4644
rect 82964 4632 82970 4684
rect 89714 4632 89720 4684
rect 89772 4672 89778 4684
rect 90177 4675 90235 4681
rect 90177 4672 90189 4675
rect 89772 4644 90189 4672
rect 89772 4632 89778 4644
rect 90177 4641 90189 4644
rect 90223 4641 90235 4675
rect 93394 4672 93400 4684
rect 93355 4644 93400 4672
rect 90177 4635 90235 4641
rect 93394 4632 93400 4644
rect 93452 4632 93458 4684
rect 93946 4632 93952 4684
rect 94004 4672 94010 4684
rect 94041 4675 94099 4681
rect 94041 4672 94053 4675
rect 94004 4644 94053 4672
rect 94004 4632 94010 4644
rect 94041 4641 94053 4644
rect 94087 4641 94099 4675
rect 94041 4635 94099 4641
rect 94590 4632 94596 4684
rect 94648 4672 94654 4684
rect 94685 4675 94743 4681
rect 94685 4672 94697 4675
rect 94648 4644 94697 4672
rect 94648 4632 94654 4644
rect 94685 4641 94697 4644
rect 94731 4641 94743 4675
rect 94685 4635 94743 4641
rect 95234 4632 95240 4684
rect 95292 4672 95298 4684
rect 95329 4675 95387 4681
rect 95329 4672 95341 4675
rect 95292 4644 95341 4672
rect 95292 4632 95298 4644
rect 95329 4641 95341 4644
rect 95375 4641 95387 4675
rect 95329 4635 95387 4641
rect 95786 4632 95792 4684
rect 95844 4672 95850 4684
rect 95973 4675 96031 4681
rect 95973 4672 95985 4675
rect 95844 4644 95985 4672
rect 95844 4632 95850 4644
rect 95973 4641 95985 4644
rect 96019 4641 96031 4675
rect 95973 4635 96031 4641
rect 96617 4675 96675 4681
rect 96617 4641 96629 4675
rect 96663 4672 96675 4675
rect 96706 4672 96712 4684
rect 96663 4644 96712 4672
rect 96663 4641 96675 4644
rect 96617 4635 96675 4641
rect 96706 4632 96712 4644
rect 96764 4632 96770 4684
rect 97258 4672 97264 4684
rect 97219 4644 97264 4672
rect 97258 4632 97264 4644
rect 97316 4632 97322 4684
rect 16298 4604 16304 4616
rect 15120 4576 16304 4604
rect 12492 4564 12498 4576
rect 16298 4564 16304 4576
rect 16356 4564 16362 4616
rect 16942 4564 16948 4616
rect 17000 4604 17006 4616
rect 20714 4604 20720 4616
rect 17000 4576 20720 4604
rect 17000 4564 17006 4576
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 41969 4607 42027 4613
rect 41969 4573 41981 4607
rect 42015 4604 42027 4607
rect 58526 4604 58532 4616
rect 42015 4576 58532 4604
rect 42015 4573 42027 4576
rect 41969 4567 42027 4573
rect 58526 4564 58532 4576
rect 58584 4564 58590 4616
rect 18506 4536 18512 4548
rect 2746 4508 18512 4536
rect 18506 4496 18512 4508
rect 18564 4496 18570 4548
rect 43257 4539 43315 4545
rect 43257 4505 43269 4539
rect 43303 4536 43315 4539
rect 55858 4536 55864 4548
rect 43303 4508 55864 4536
rect 43303 4505 43315 4508
rect 43257 4499 43315 4505
rect 55858 4496 55864 4508
rect 55916 4496 55922 4548
rect 60706 4508 74534 4536
rect 4341 4471 4399 4477
rect 4341 4437 4353 4471
rect 4387 4468 4399 4471
rect 4614 4468 4620 4480
rect 4387 4440 4620 4468
rect 4387 4437 4399 4440
rect 4341 4431 4399 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 5074 4468 5080 4480
rect 5035 4440 5080 4468
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 7561 4471 7619 4477
rect 7561 4468 7573 4471
rect 7524 4440 7573 4468
rect 7524 4428 7530 4440
rect 7561 4437 7573 4440
rect 7607 4437 7619 4471
rect 7561 4431 7619 4437
rect 11606 4428 11612 4480
rect 11664 4468 11670 4480
rect 11977 4471 12035 4477
rect 11977 4468 11989 4471
rect 11664 4440 11989 4468
rect 11664 4428 11670 4440
rect 11977 4437 11989 4440
rect 12023 4437 12035 4471
rect 11977 4431 12035 4437
rect 17126 4428 17132 4480
rect 17184 4468 17190 4480
rect 17313 4471 17371 4477
rect 17313 4468 17325 4471
rect 17184 4440 17325 4468
rect 17184 4428 17190 4440
rect 17313 4437 17325 4440
rect 17359 4437 17371 4471
rect 17313 4431 17371 4437
rect 48498 4428 48504 4480
rect 48556 4468 48562 4480
rect 60706 4468 60734 4508
rect 65150 4468 65156 4480
rect 48556 4440 60734 4468
rect 65111 4440 65156 4468
rect 48556 4428 48562 4440
rect 65150 4428 65156 4440
rect 65208 4428 65214 4480
rect 74506 4468 74534 4508
rect 89717 4471 89775 4477
rect 89717 4468 89729 4471
rect 74506 4440 89729 4468
rect 89717 4437 89729 4440
rect 89763 4437 89775 4471
rect 89717 4431 89775 4437
rect 1104 4378 98808 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 65686 4378
rect 65738 4326 65750 4378
rect 65802 4326 65814 4378
rect 65866 4326 65878 4378
rect 65930 4326 96406 4378
rect 96458 4326 96470 4378
rect 96522 4326 96534 4378
rect 96586 4326 96598 4378
rect 96650 4326 98808 4378
rect 1104 4304 98808 4326
rect 3602 4224 3608 4276
rect 3660 4264 3666 4276
rect 29730 4264 29736 4276
rect 3660 4236 29736 4264
rect 3660 4224 3666 4236
rect 29730 4224 29736 4236
rect 29788 4224 29794 4276
rect 48130 4224 48136 4276
rect 48188 4264 48194 4276
rect 65150 4264 65156 4276
rect 48188 4236 65156 4264
rect 48188 4224 48194 4236
rect 65150 4224 65156 4236
rect 65208 4224 65214 4276
rect 69934 4224 69940 4276
rect 69992 4224 69998 4276
rect 69952 4196 69980 4224
rect 70670 4196 70676 4208
rect 69952 4168 70676 4196
rect 70670 4156 70676 4168
rect 70728 4156 70734 4208
rect 82354 4156 82360 4208
rect 82412 4196 82418 4208
rect 84746 4196 84752 4208
rect 82412 4168 84752 4196
rect 82412 4156 82418 4168
rect 84746 4156 84752 4168
rect 84804 4156 84810 4208
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 2590 4128 2596 4140
rect 1719 4100 2452 4128
rect 2551 4100 2596 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 658 4020 664 4072
rect 716 4060 722 4072
rect 1397 4063 1455 4069
rect 1397 4060 1409 4063
rect 716 4032 1409 4060
rect 716 4020 722 4032
rect 1397 4029 1409 4032
rect 1443 4029 1455 4063
rect 1397 4023 1455 4029
rect 1486 4020 1492 4072
rect 1544 4060 1550 4072
rect 2317 4063 2375 4069
rect 2317 4060 2329 4063
rect 1544 4032 2329 4060
rect 1544 4020 1550 4032
rect 2317 4029 2329 4032
rect 2363 4029 2375 4063
rect 2424 4060 2452 4100
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 3418 4128 3424 4140
rect 2700 4100 3424 4128
rect 2700 4060 2728 4100
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 11974 4128 11980 4140
rect 11935 4100 11980 4128
rect 11974 4088 11980 4100
rect 12032 4128 12038 4140
rect 12032 4100 12296 4128
rect 12032 4088 12038 4100
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 2424 4032 2728 4060
rect 3252 4032 4261 4060
rect 2317 4023 2375 4029
rect 2498 3952 2504 4004
rect 2556 3992 2562 4004
rect 3252 3992 3280 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 5166 4060 5172 4072
rect 5127 4032 5172 4060
rect 4249 4023 4307 4029
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 6362 4020 6368 4072
rect 6420 4060 6426 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6420 4032 6837 4060
rect 6420 4020 6426 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 7650 4060 7656 4072
rect 7611 4032 7656 4060
rect 6825 4023 6883 4029
rect 7650 4020 7656 4032
rect 7708 4020 7714 4072
rect 8386 4060 8392 4072
rect 8347 4032 8392 4060
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8846 4020 8852 4072
rect 8904 4060 8910 4072
rect 9033 4063 9091 4069
rect 9033 4060 9045 4063
rect 8904 4032 9045 4060
rect 8904 4020 8910 4032
rect 9033 4029 9045 4032
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9456 4032 9689 4060
rect 9456 4020 9462 4032
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 10502 4060 10508 4072
rect 10463 4032 10508 4060
rect 9677 4023 9735 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 12268 4069 12296 4100
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 13541 4131 13599 4137
rect 13541 4128 13553 4131
rect 13044 4100 13553 4128
rect 13044 4088 13050 4100
rect 13541 4097 13553 4100
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 69934 4088 69940 4140
rect 69992 4128 69998 4140
rect 81618 4128 81624 4140
rect 69992 4100 80652 4128
rect 81579 4100 81624 4128
rect 69992 4088 69998 4100
rect 12253 4063 12311 4069
rect 12253 4029 12265 4063
rect 12299 4029 12311 4063
rect 12253 4023 12311 4029
rect 12710 4020 12716 4072
rect 12768 4060 12774 4072
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12768 4032 12909 4060
rect 12768 4020 12774 4032
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 13449 4063 13507 4069
rect 13449 4029 13461 4063
rect 13495 4060 13507 4063
rect 13722 4060 13728 4072
rect 13495 4032 13728 4060
rect 13495 4029 13507 4032
rect 13449 4023 13507 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 14366 4060 14372 4072
rect 14327 4032 14372 4060
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4029 15071 4063
rect 16022 4060 16028 4072
rect 15983 4032 16028 4060
rect 15013 4023 15071 4029
rect 2556 3964 3280 3992
rect 3329 3995 3387 4001
rect 2556 3952 2562 3964
rect 3329 3961 3341 3995
rect 3375 3992 3387 3995
rect 3970 3992 3976 4004
rect 3375 3964 3976 3992
rect 3375 3961 3387 3964
rect 3329 3955 3387 3961
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 4065 3995 4123 4001
rect 4065 3961 4077 3995
rect 4111 3992 4123 3995
rect 6086 3992 6092 4004
rect 4111 3964 6092 3992
rect 4111 3961 4123 3964
rect 4065 3955 4123 3961
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 6730 3952 6736 4004
rect 6788 3992 6794 4004
rect 7837 3995 7895 4001
rect 7837 3992 7849 3995
rect 6788 3964 7849 3992
rect 6788 3952 6794 3964
rect 7837 3961 7849 3964
rect 7883 3961 7895 3995
rect 7837 3955 7895 3961
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 12069 3995 12127 4001
rect 12069 3992 12081 3995
rect 11112 3964 12081 3992
rect 11112 3952 11118 3964
rect 12069 3961 12081 3964
rect 12115 3961 12127 3995
rect 12069 3955 12127 3961
rect 13630 3952 13636 4004
rect 13688 3992 13694 4004
rect 15028 3992 15056 4023
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 17402 4060 17408 4072
rect 17363 4032 17408 4060
rect 17402 4020 17408 4032
rect 17460 4020 17466 4072
rect 18046 4020 18052 4072
rect 18104 4060 18110 4072
rect 18141 4063 18199 4069
rect 18141 4060 18153 4063
rect 18104 4032 18153 4060
rect 18104 4020 18110 4032
rect 18141 4029 18153 4032
rect 18187 4029 18199 4063
rect 18874 4060 18880 4072
rect 18835 4032 18880 4060
rect 18141 4023 18199 4029
rect 18874 4020 18880 4032
rect 18932 4020 18938 4072
rect 19613 4063 19671 4069
rect 19613 4029 19625 4063
rect 19659 4060 19671 4063
rect 19886 4060 19892 4072
rect 19659 4032 19892 4060
rect 19659 4029 19671 4032
rect 19613 4023 19671 4029
rect 19886 4020 19892 4032
rect 19944 4020 19950 4072
rect 20070 4020 20076 4072
rect 20128 4060 20134 4072
rect 20993 4063 21051 4069
rect 20993 4060 21005 4063
rect 20128 4032 21005 4060
rect 20128 4020 20134 4032
rect 20993 4029 21005 4032
rect 21039 4029 21051 4063
rect 20993 4023 21051 4029
rect 22002 4020 22008 4072
rect 22060 4060 22066 4072
rect 22557 4063 22615 4069
rect 22557 4060 22569 4063
rect 22060 4032 22569 4060
rect 22060 4020 22066 4032
rect 22557 4029 22569 4032
rect 22603 4029 22615 4063
rect 22557 4023 22615 4029
rect 22830 4020 22836 4072
rect 22888 4060 22894 4072
rect 23201 4063 23259 4069
rect 23201 4060 23213 4063
rect 22888 4032 23213 4060
rect 22888 4020 22894 4032
rect 23201 4029 23213 4032
rect 23247 4029 23259 4063
rect 23201 4023 23259 4029
rect 23290 4020 23296 4072
rect 23348 4060 23354 4072
rect 23845 4063 23903 4069
rect 23845 4060 23857 4063
rect 23348 4032 23857 4060
rect 23348 4020 23354 4032
rect 23845 4029 23857 4032
rect 23891 4029 23903 4063
rect 23845 4023 23903 4029
rect 23934 4020 23940 4072
rect 23992 4060 23998 4072
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 23992 4032 24501 4060
rect 23992 4020 23998 4032
rect 24489 4029 24501 4032
rect 24535 4029 24547 4063
rect 24489 4023 24547 4029
rect 24578 4020 24584 4072
rect 24636 4060 24642 4072
rect 25133 4063 25191 4069
rect 25133 4060 25145 4063
rect 24636 4032 25145 4060
rect 24636 4020 24642 4032
rect 25133 4029 25145 4032
rect 25179 4029 25191 4063
rect 25866 4060 25872 4072
rect 25827 4032 25872 4060
rect 25133 4023 25191 4029
rect 25866 4020 25872 4032
rect 25924 4020 25930 4072
rect 26510 4060 26516 4072
rect 26471 4032 26516 4060
rect 26510 4020 26516 4032
rect 26568 4020 26574 4072
rect 27522 4020 27528 4072
rect 27580 4060 27586 4072
rect 27801 4063 27859 4069
rect 27801 4060 27813 4063
rect 27580 4032 27813 4060
rect 27580 4020 27586 4032
rect 27801 4029 27813 4032
rect 27847 4029 27859 4063
rect 28718 4060 28724 4072
rect 28679 4032 28724 4060
rect 27801 4023 27859 4029
rect 28718 4020 28724 4032
rect 28776 4020 28782 4072
rect 29362 4060 29368 4072
rect 29323 4032 29368 4060
rect 29362 4020 29368 4032
rect 29420 4020 29426 4072
rect 30558 4060 30564 4072
rect 30519 4032 30564 4060
rect 30558 4020 30564 4032
rect 30616 4020 30622 4072
rect 31202 4060 31208 4072
rect 31163 4032 31208 4060
rect 31202 4020 31208 4032
rect 31260 4020 31266 4072
rect 31754 4020 31760 4072
rect 31812 4060 31818 4072
rect 31849 4063 31907 4069
rect 31849 4060 31861 4063
rect 31812 4032 31861 4060
rect 31812 4020 31818 4032
rect 31849 4029 31861 4032
rect 31895 4029 31907 4063
rect 33594 4060 33600 4072
rect 33555 4032 33600 4060
rect 31849 4023 31907 4029
rect 33594 4020 33600 4032
rect 33652 4020 33658 4072
rect 34238 4060 34244 4072
rect 34199 4032 34244 4060
rect 34238 4020 34244 4032
rect 34296 4020 34302 4072
rect 34790 4020 34796 4072
rect 34848 4060 34854 4072
rect 34885 4063 34943 4069
rect 34885 4060 34897 4063
rect 34848 4032 34897 4060
rect 34848 4020 34854 4032
rect 34885 4029 34897 4032
rect 34931 4029 34943 4063
rect 34885 4023 34943 4029
rect 35434 4020 35440 4072
rect 35492 4060 35498 4072
rect 35529 4063 35587 4069
rect 35529 4060 35541 4063
rect 35492 4032 35541 4060
rect 35492 4020 35498 4032
rect 35529 4029 35541 4032
rect 35575 4029 35587 4063
rect 35529 4023 35587 4029
rect 36078 4020 36084 4072
rect 36136 4060 36142 4072
rect 36173 4063 36231 4069
rect 36173 4060 36185 4063
rect 36136 4032 36185 4060
rect 36136 4020 36142 4032
rect 36173 4029 36185 4032
rect 36219 4029 36231 4063
rect 36173 4023 36231 4029
rect 36630 4020 36636 4072
rect 36688 4060 36694 4072
rect 36817 4063 36875 4069
rect 36817 4060 36829 4063
rect 36688 4032 36829 4060
rect 36688 4020 36694 4032
rect 36817 4029 36829 4032
rect 36863 4029 36875 4063
rect 36817 4023 36875 4029
rect 37826 4020 37832 4072
rect 37884 4060 37890 4072
rect 38289 4063 38347 4069
rect 38289 4060 38301 4063
rect 37884 4032 38301 4060
rect 37884 4020 37890 4032
rect 38289 4029 38301 4032
rect 38335 4029 38347 4063
rect 38289 4023 38347 4029
rect 38470 4020 38476 4072
rect 38528 4060 38534 4072
rect 38933 4063 38991 4069
rect 38933 4060 38945 4063
rect 38528 4032 38945 4060
rect 38528 4020 38534 4032
rect 38933 4029 38945 4032
rect 38979 4029 38991 4063
rect 39942 4060 39948 4072
rect 39903 4032 39948 4060
rect 38933 4023 38991 4029
rect 39942 4020 39948 4032
rect 40000 4020 40006 4072
rect 40310 4020 40316 4072
rect 40368 4060 40374 4072
rect 40589 4063 40647 4069
rect 40589 4060 40601 4063
rect 40368 4032 40601 4060
rect 40368 4020 40374 4032
rect 40589 4029 40601 4032
rect 40635 4029 40647 4063
rect 40589 4023 40647 4029
rect 40954 4020 40960 4072
rect 41012 4060 41018 4072
rect 41233 4063 41291 4069
rect 41233 4060 41245 4063
rect 41012 4032 41245 4060
rect 41012 4020 41018 4032
rect 41233 4029 41245 4032
rect 41279 4029 41291 4063
rect 41233 4023 41291 4029
rect 41506 4020 41512 4072
rect 41564 4060 41570 4072
rect 41877 4063 41935 4069
rect 41877 4060 41889 4063
rect 41564 4032 41889 4060
rect 41564 4020 41570 4032
rect 41877 4029 41889 4032
rect 41923 4029 41935 4063
rect 41877 4023 41935 4029
rect 42702 4020 42708 4072
rect 42760 4060 42766 4072
rect 43533 4063 43591 4069
rect 43533 4060 43545 4063
rect 42760 4032 43545 4060
rect 42760 4020 42766 4032
rect 43533 4029 43545 4032
rect 43579 4029 43591 4063
rect 43533 4023 43591 4029
rect 44177 4063 44235 4069
rect 44177 4029 44189 4063
rect 44223 4029 44235 4063
rect 44177 4023 44235 4029
rect 44821 4063 44879 4069
rect 44821 4029 44833 4063
rect 44867 4029 44879 4063
rect 46014 4060 46020 4072
rect 45975 4032 46020 4060
rect 44821 4023 44879 4029
rect 13688 3964 15056 3992
rect 20349 3995 20407 4001
rect 13688 3952 13694 3964
rect 20349 3961 20361 3995
rect 20395 3992 20407 3995
rect 20622 3992 20628 4004
rect 20395 3964 20628 3992
rect 20395 3961 20407 3964
rect 20349 3955 20407 3961
rect 20622 3952 20628 3964
rect 20680 3952 20686 4004
rect 43346 3952 43352 4004
rect 43404 3992 43410 4004
rect 44192 3992 44220 4023
rect 43404 3964 44220 3992
rect 43404 3952 43410 3964
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 1820 3896 3433 3924
rect 1820 3884 1826 3896
rect 3421 3893 3433 3896
rect 3467 3893 3479 3927
rect 5350 3924 5356 3936
rect 5311 3896 5356 3924
rect 3421 3887 3479 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 7009 3927 7067 3933
rect 7009 3893 7021 3927
rect 7055 3924 7067 3927
rect 7190 3924 7196 3936
rect 7055 3896 7196 3924
rect 7055 3893 7067 3896
rect 7009 3887 7067 3893
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 8481 3927 8539 3933
rect 8481 3924 8493 3927
rect 8076 3896 8493 3924
rect 8076 3884 8082 3896
rect 8481 3893 8493 3896
rect 8527 3893 8539 3927
rect 8481 3887 8539 3893
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 10597 3927 10655 3933
rect 10597 3924 10609 3927
rect 10560 3896 10609 3924
rect 10560 3884 10566 3896
rect 10597 3893 10609 3896
rect 10643 3893 10655 3927
rect 10597 3887 10655 3893
rect 12342 3884 12348 3936
rect 12400 3924 12406 3936
rect 12989 3927 13047 3933
rect 12989 3924 13001 3927
rect 12400 3896 13001 3924
rect 12400 3884 12406 3896
rect 12989 3893 13001 3896
rect 13035 3893 13047 3927
rect 12989 3887 13047 3893
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 14461 3927 14519 3933
rect 14461 3924 14473 3927
rect 13504 3896 14473 3924
rect 13504 3884 13510 3896
rect 14461 3893 14473 3896
rect 14507 3893 14519 3927
rect 14461 3887 14519 3893
rect 15930 3884 15936 3936
rect 15988 3924 15994 3936
rect 16117 3927 16175 3933
rect 16117 3924 16129 3927
rect 15988 3896 16129 3924
rect 15988 3884 15994 3896
rect 16117 3893 16129 3896
rect 16163 3893 16175 3927
rect 16117 3887 16175 3893
rect 16390 3884 16396 3936
rect 16448 3924 16454 3936
rect 17497 3927 17555 3933
rect 17497 3924 17509 3927
rect 16448 3896 17509 3924
rect 16448 3884 16454 3896
rect 17497 3893 17509 3896
rect 17543 3893 17555 3927
rect 17497 3887 17555 3893
rect 17770 3884 17776 3936
rect 17828 3924 17834 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 17828 3896 18245 3924
rect 17828 3884 17834 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18233 3887 18291 3893
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 18969 3927 19027 3933
rect 18969 3924 18981 3927
rect 18380 3896 18981 3924
rect 18380 3884 18386 3896
rect 18969 3893 18981 3896
rect 19015 3893 19027 3927
rect 18969 3887 19027 3893
rect 19058 3884 19064 3936
rect 19116 3924 19122 3936
rect 19705 3927 19763 3933
rect 19705 3924 19717 3927
rect 19116 3896 19717 3924
rect 19116 3884 19122 3896
rect 19705 3893 19717 3896
rect 19751 3893 19763 3927
rect 19705 3887 19763 3893
rect 19978 3884 19984 3936
rect 20036 3924 20042 3936
rect 20441 3927 20499 3933
rect 20441 3924 20453 3927
rect 20036 3896 20453 3924
rect 20036 3884 20042 3896
rect 20441 3893 20453 3896
rect 20487 3893 20499 3927
rect 20441 3887 20499 3893
rect 43990 3884 43996 3936
rect 44048 3924 44054 3936
rect 44836 3924 44864 4023
rect 46014 4020 46020 4032
rect 46072 4020 46078 4072
rect 46661 4063 46719 4069
rect 46661 4029 46673 4063
rect 46707 4029 46719 4063
rect 46661 4023 46719 4029
rect 47305 4063 47363 4069
rect 47305 4029 47317 4063
rect 47351 4029 47363 4063
rect 47305 4023 47363 4029
rect 45186 3952 45192 4004
rect 45244 3992 45250 4004
rect 46676 3992 46704 4023
rect 45244 3964 46704 3992
rect 45244 3952 45250 3964
rect 44048 3896 44864 3924
rect 44048 3884 44054 3896
rect 46382 3884 46388 3936
rect 46440 3924 46446 3936
rect 47320 3924 47348 4023
rect 48406 4020 48412 4072
rect 48464 4060 48470 4072
rect 48777 4063 48835 4069
rect 48777 4060 48789 4063
rect 48464 4032 48789 4060
rect 48464 4020 48470 4032
rect 48777 4029 48789 4032
rect 48823 4029 48835 4063
rect 48777 4023 48835 4029
rect 48866 4020 48872 4072
rect 48924 4060 48930 4072
rect 49421 4063 49479 4069
rect 49421 4060 49433 4063
rect 48924 4032 49433 4060
rect 48924 4020 48930 4032
rect 49421 4029 49433 4032
rect 49467 4029 49479 4063
rect 49421 4023 49479 4029
rect 49602 4020 49608 4072
rect 49660 4060 49666 4072
rect 50065 4063 50123 4069
rect 50065 4060 50077 4063
rect 49660 4032 50077 4060
rect 49660 4020 49666 4032
rect 50065 4029 50077 4032
rect 50111 4029 50123 4063
rect 50065 4023 50123 4029
rect 50154 4020 50160 4072
rect 50212 4060 50218 4072
rect 50709 4063 50767 4069
rect 50709 4060 50721 4063
rect 50212 4032 50721 4060
rect 50212 4020 50218 4032
rect 50709 4029 50721 4032
rect 50755 4029 50767 4063
rect 50709 4023 50767 4029
rect 50798 4020 50804 4072
rect 50856 4060 50862 4072
rect 51353 4063 51411 4069
rect 51353 4060 51365 4063
rect 50856 4032 51365 4060
rect 50856 4020 50862 4032
rect 51353 4029 51365 4032
rect 51399 4029 51411 4063
rect 51353 4023 51411 4029
rect 51442 4020 51448 4072
rect 51500 4060 51506 4072
rect 51997 4063 52055 4069
rect 51997 4060 52009 4063
rect 51500 4032 52009 4060
rect 51500 4020 51506 4032
rect 51997 4029 52009 4032
rect 52043 4029 52055 4063
rect 51997 4023 52055 4029
rect 52641 4063 52699 4069
rect 52641 4029 52653 4063
rect 52687 4029 52699 4063
rect 52641 4023 52699 4029
rect 51902 3952 51908 4004
rect 51960 3992 51966 4004
rect 52656 3992 52684 4023
rect 53742 4020 53748 4072
rect 53800 4060 53806 4072
rect 54021 4063 54079 4069
rect 54021 4060 54033 4063
rect 53800 4032 54033 4060
rect 53800 4020 53806 4032
rect 54021 4029 54033 4032
rect 54067 4029 54079 4063
rect 54021 4023 54079 4029
rect 54294 4020 54300 4072
rect 54352 4060 54358 4072
rect 54665 4063 54723 4069
rect 54665 4060 54677 4063
rect 54352 4032 54677 4060
rect 54352 4020 54358 4032
rect 54665 4029 54677 4032
rect 54711 4029 54723 4063
rect 54665 4023 54723 4029
rect 54938 4020 54944 4072
rect 54996 4060 55002 4072
rect 55309 4063 55367 4069
rect 55309 4060 55321 4063
rect 54996 4032 55321 4060
rect 54996 4020 55002 4032
rect 55309 4029 55321 4032
rect 55355 4029 55367 4063
rect 55309 4023 55367 4029
rect 55582 4020 55588 4072
rect 55640 4060 55646 4072
rect 55953 4063 56011 4069
rect 55953 4060 55965 4063
rect 55640 4032 55965 4060
rect 55640 4020 55646 4032
rect 55953 4029 55965 4032
rect 55999 4029 56011 4063
rect 55953 4023 56011 4029
rect 56134 4020 56140 4072
rect 56192 4060 56198 4072
rect 56597 4063 56655 4069
rect 56597 4060 56609 4063
rect 56192 4032 56609 4060
rect 56192 4020 56198 4032
rect 56597 4029 56609 4032
rect 56643 4029 56655 4063
rect 56597 4023 56655 4029
rect 56778 4020 56784 4072
rect 56836 4060 56842 4072
rect 57241 4063 57299 4069
rect 57241 4060 57253 4063
rect 56836 4032 57253 4060
rect 56836 4020 56842 4032
rect 57241 4029 57253 4032
rect 57287 4029 57299 4063
rect 57241 4023 57299 4029
rect 57422 4020 57428 4072
rect 57480 4060 57486 4072
rect 57885 4063 57943 4069
rect 57885 4060 57897 4063
rect 57480 4032 57897 4060
rect 57480 4020 57486 4032
rect 57885 4029 57897 4032
rect 57931 4029 57943 4063
rect 57885 4023 57943 4029
rect 58618 4020 58624 4072
rect 58676 4060 58682 4072
rect 59265 4063 59323 4069
rect 59265 4060 59277 4063
rect 58676 4032 59277 4060
rect 58676 4020 58682 4032
rect 59265 4029 59277 4032
rect 59311 4029 59323 4063
rect 59909 4063 59967 4069
rect 59909 4060 59921 4063
rect 59265 4023 59323 4029
rect 59372 4032 59921 4060
rect 51960 3964 52684 3992
rect 51960 3952 51966 3964
rect 59170 3952 59176 4004
rect 59228 3992 59234 4004
rect 59372 3992 59400 4032
rect 59909 4029 59921 4032
rect 59955 4029 59967 4063
rect 59909 4023 59967 4029
rect 60553 4063 60611 4069
rect 60553 4029 60565 4063
rect 60599 4029 60611 4063
rect 61197 4063 61255 4069
rect 61197 4060 61209 4063
rect 60553 4023 60611 4029
rect 60706 4032 61209 4060
rect 59228 3964 59400 3992
rect 59228 3952 59234 3964
rect 59814 3952 59820 4004
rect 59872 3992 59878 4004
rect 60568 3992 60596 4023
rect 59872 3964 60596 3992
rect 59872 3952 59878 3964
rect 46440 3896 47348 3924
rect 46440 3884 46446 3896
rect 60458 3884 60464 3936
rect 60516 3924 60522 3936
rect 60706 3924 60734 4032
rect 61197 4029 61209 4032
rect 61243 4029 61255 4063
rect 61841 4063 61899 4069
rect 61841 4060 61853 4063
rect 61197 4023 61255 4029
rect 61304 4032 61853 4060
rect 61010 3952 61016 4004
rect 61068 3992 61074 4004
rect 61304 3992 61332 4032
rect 61841 4029 61853 4032
rect 61887 4029 61899 4063
rect 61841 4023 61899 4029
rect 62485 4063 62543 4069
rect 62485 4029 62497 4063
rect 62531 4029 62543 4063
rect 62485 4023 62543 4029
rect 63129 4063 63187 4069
rect 63129 4029 63141 4063
rect 63175 4029 63187 4063
rect 63129 4023 63187 4029
rect 61068 3964 61332 3992
rect 61068 3952 61074 3964
rect 61746 3952 61752 4004
rect 61804 3992 61810 4004
rect 62500 3992 62528 4023
rect 61804 3964 62528 3992
rect 61804 3952 61810 3964
rect 60516 3896 60734 3924
rect 60516 3884 60522 3896
rect 62298 3884 62304 3936
rect 62356 3924 62362 3936
rect 63144 3924 63172 4023
rect 64138 4020 64144 4072
rect 64196 4060 64202 4072
rect 64509 4063 64567 4069
rect 64509 4060 64521 4063
rect 64196 4032 64521 4060
rect 64196 4020 64202 4032
rect 64509 4029 64521 4032
rect 64555 4029 64567 4063
rect 64509 4023 64567 4029
rect 64782 4020 64788 4072
rect 64840 4060 64846 4072
rect 65153 4063 65211 4069
rect 65153 4060 65165 4063
rect 64840 4032 65165 4060
rect 64840 4020 64846 4032
rect 65153 4029 65165 4032
rect 65199 4029 65211 4063
rect 65153 4023 65211 4029
rect 65889 4063 65947 4069
rect 65889 4029 65901 4063
rect 65935 4060 65947 4063
rect 65978 4060 65984 4072
rect 65935 4032 65984 4060
rect 65935 4029 65947 4032
rect 65889 4023 65947 4029
rect 65978 4020 65984 4032
rect 66036 4020 66042 4072
rect 66530 4060 66536 4072
rect 66491 4032 66536 4060
rect 66530 4020 66536 4032
rect 66588 4020 66594 4072
rect 67174 4060 67180 4072
rect 67135 4032 67180 4060
rect 67174 4020 67180 4032
rect 67232 4020 67238 4072
rect 67726 4020 67732 4072
rect 67784 4060 67790 4072
rect 67821 4063 67879 4069
rect 67821 4060 67833 4063
rect 67784 4032 67833 4060
rect 67784 4020 67790 4032
rect 67821 4029 67833 4032
rect 67867 4029 67879 4063
rect 68462 4060 68468 4072
rect 68423 4032 68468 4060
rect 67821 4023 67879 4029
rect 68462 4020 68468 4032
rect 68520 4020 68526 4072
rect 68922 4020 68928 4072
rect 68980 4060 68986 4072
rect 69753 4063 69811 4069
rect 69753 4060 69765 4063
rect 68980 4032 69765 4060
rect 68980 4020 68986 4032
rect 69753 4029 69765 4032
rect 69799 4029 69811 4063
rect 69753 4023 69811 4029
rect 70397 4063 70455 4069
rect 70397 4029 70409 4063
rect 70443 4029 70455 4063
rect 70397 4023 70455 4029
rect 69566 3952 69572 4004
rect 69624 3992 69630 4004
rect 70412 3992 70440 4023
rect 70762 4020 70768 4072
rect 70820 4060 70826 4072
rect 71041 4063 71099 4069
rect 71041 4060 71053 4063
rect 70820 4032 71053 4060
rect 70820 4020 70826 4032
rect 71041 4029 71053 4032
rect 71087 4029 71099 4063
rect 71041 4023 71099 4029
rect 71406 4020 71412 4072
rect 71464 4060 71470 4072
rect 71685 4063 71743 4069
rect 71685 4060 71697 4063
rect 71464 4032 71697 4060
rect 71464 4020 71470 4032
rect 71685 4029 71697 4032
rect 71731 4029 71743 4063
rect 71685 4023 71743 4029
rect 72050 4020 72056 4072
rect 72108 4060 72114 4072
rect 72329 4063 72387 4069
rect 72329 4060 72341 4063
rect 72108 4032 72341 4060
rect 72108 4020 72114 4032
rect 72329 4029 72341 4032
rect 72375 4029 72387 4063
rect 72329 4023 72387 4029
rect 72602 4020 72608 4072
rect 72660 4060 72666 4072
rect 72973 4063 73031 4069
rect 72973 4060 72985 4063
rect 72660 4032 72985 4060
rect 72660 4020 72666 4032
rect 72973 4029 72985 4032
rect 73019 4029 73031 4063
rect 72973 4023 73031 4029
rect 73246 4020 73252 4072
rect 73304 4060 73310 4072
rect 73617 4063 73675 4069
rect 73617 4060 73629 4063
rect 73304 4032 73629 4060
rect 73304 4020 73310 4032
rect 73617 4029 73629 4032
rect 73663 4029 73675 4063
rect 73617 4023 73675 4029
rect 74442 4020 74448 4072
rect 74500 4060 74506 4072
rect 74997 4063 75055 4069
rect 74997 4060 75009 4063
rect 74500 4032 75009 4060
rect 74500 4020 74506 4032
rect 74997 4029 75009 4032
rect 75043 4029 75055 4063
rect 74997 4023 75055 4029
rect 75086 4020 75092 4072
rect 75144 4060 75150 4072
rect 75641 4063 75699 4069
rect 75641 4060 75653 4063
rect 75144 4032 75653 4060
rect 75144 4020 75150 4032
rect 75641 4029 75653 4032
rect 75687 4029 75699 4063
rect 75641 4023 75699 4029
rect 75730 4020 75736 4072
rect 75788 4060 75794 4072
rect 76285 4063 76343 4069
rect 76285 4060 76297 4063
rect 75788 4032 76297 4060
rect 75788 4020 75794 4032
rect 76285 4029 76297 4032
rect 76331 4029 76343 4063
rect 76285 4023 76343 4029
rect 76374 4020 76380 4072
rect 76432 4060 76438 4072
rect 76929 4063 76987 4069
rect 76929 4060 76941 4063
rect 76432 4032 76941 4060
rect 76432 4020 76438 4032
rect 76929 4029 76941 4032
rect 76975 4029 76987 4063
rect 76929 4023 76987 4029
rect 77018 4020 77024 4072
rect 77076 4060 77082 4072
rect 77573 4063 77631 4069
rect 77573 4060 77585 4063
rect 77076 4032 77585 4060
rect 77076 4020 77082 4032
rect 77573 4029 77585 4032
rect 77619 4029 77631 4063
rect 77573 4023 77631 4029
rect 77662 4020 77668 4072
rect 77720 4060 77726 4072
rect 78217 4063 78275 4069
rect 78217 4060 78229 4063
rect 77720 4032 78229 4060
rect 77720 4020 77726 4032
rect 78217 4029 78229 4032
rect 78263 4029 78275 4063
rect 78217 4023 78275 4029
rect 78861 4063 78919 4069
rect 78861 4029 78873 4063
rect 78907 4029 78919 4063
rect 80238 4060 80244 4072
rect 80199 4032 80244 4060
rect 78861 4023 78919 4029
rect 69624 3964 70440 3992
rect 69624 3952 69630 3964
rect 78122 3952 78128 4004
rect 78180 3992 78186 4004
rect 78876 3992 78904 4023
rect 80238 4020 80244 4032
rect 80296 4020 80302 4072
rect 80330 4020 80336 4072
rect 80388 4060 80394 4072
rect 80517 4063 80575 4069
rect 80517 4060 80529 4063
rect 80388 4032 80529 4060
rect 80388 4020 80394 4032
rect 80517 4029 80529 4032
rect 80563 4029 80575 4063
rect 80624 4060 80652 4100
rect 81618 4088 81624 4100
rect 81676 4088 81682 4140
rect 83550 4128 83556 4140
rect 81728 4100 83556 4128
rect 81728 4060 81756 4100
rect 83550 4088 83556 4100
rect 83608 4088 83614 4140
rect 96801 4131 96859 4137
rect 96801 4097 96813 4131
rect 96847 4128 96859 4131
rect 96890 4128 96896 4140
rect 96847 4100 96896 4128
rect 96847 4097 96859 4100
rect 96801 4091 96859 4097
rect 96890 4088 96896 4100
rect 96948 4088 96954 4140
rect 97445 4131 97503 4137
rect 97445 4128 97457 4131
rect 97184 4100 97457 4128
rect 80624 4032 81756 4060
rect 80517 4023 80575 4029
rect 81986 4020 81992 4072
rect 82044 4060 82050 4072
rect 82357 4063 82415 4069
rect 82357 4060 82369 4063
rect 82044 4032 82369 4060
rect 82044 4020 82050 4032
rect 82357 4029 82369 4032
rect 82403 4029 82415 4063
rect 82357 4023 82415 4029
rect 83001 4063 83059 4069
rect 83001 4029 83013 4063
rect 83047 4029 83059 4063
rect 83642 4060 83648 4072
rect 83603 4032 83648 4060
rect 83001 4023 83059 4029
rect 78180 3964 78904 3992
rect 78180 3952 78186 3964
rect 81802 3952 81808 4004
rect 81860 3992 81866 4004
rect 83016 3992 83044 4023
rect 83642 4020 83648 4032
rect 83700 4020 83706 4072
rect 84194 4020 84200 4072
rect 84252 4060 84258 4072
rect 84289 4063 84347 4069
rect 84289 4060 84301 4063
rect 84252 4032 84301 4060
rect 84252 4020 84258 4032
rect 84289 4029 84301 4032
rect 84335 4029 84347 4063
rect 84289 4023 84347 4029
rect 84838 4020 84844 4072
rect 84896 4060 84902 4072
rect 85485 4063 85543 4069
rect 85485 4060 85497 4063
rect 84896 4032 85497 4060
rect 84896 4020 84902 4032
rect 85485 4029 85497 4032
rect 85531 4029 85543 4063
rect 85485 4023 85543 4029
rect 86129 4063 86187 4069
rect 86129 4029 86141 4063
rect 86175 4029 86187 4063
rect 86129 4023 86187 4029
rect 81860 3964 83044 3992
rect 81860 3952 81866 3964
rect 85390 3952 85396 4004
rect 85448 3992 85454 4004
rect 86144 3992 86172 4023
rect 86678 4020 86684 4072
rect 86736 4060 86742 4072
rect 86773 4063 86831 4069
rect 86773 4060 86785 4063
rect 86736 4032 86785 4060
rect 86736 4020 86742 4032
rect 86773 4029 86785 4032
rect 86819 4029 86831 4063
rect 86773 4023 86831 4029
rect 87230 4020 87236 4072
rect 87288 4060 87294 4072
rect 87417 4063 87475 4069
rect 87417 4060 87429 4063
rect 87288 4032 87429 4060
rect 87288 4020 87294 4032
rect 87417 4029 87429 4032
rect 87463 4029 87475 4063
rect 88518 4060 88524 4072
rect 88479 4032 88524 4060
rect 87417 4023 87475 4029
rect 88518 4020 88524 4032
rect 88576 4020 88582 4072
rect 89070 4020 89076 4072
rect 89128 4060 89134 4072
rect 89165 4063 89223 4069
rect 89165 4060 89177 4063
rect 89128 4032 89177 4060
rect 89128 4020 89134 4032
rect 89165 4029 89177 4032
rect 89211 4029 89223 4063
rect 89165 4023 89223 4029
rect 90266 4020 90272 4072
rect 90324 4060 90330 4072
rect 90729 4063 90787 4069
rect 90729 4060 90741 4063
rect 90324 4032 90741 4060
rect 90324 4020 90330 4032
rect 90729 4029 90741 4032
rect 90775 4029 90787 4063
rect 90729 4023 90787 4029
rect 90910 4020 90916 4072
rect 90968 4060 90974 4072
rect 91373 4063 91431 4069
rect 91373 4060 91385 4063
rect 90968 4032 91385 4060
rect 90968 4020 90974 4032
rect 91373 4029 91385 4032
rect 91419 4029 91431 4063
rect 91373 4023 91431 4029
rect 91554 4020 91560 4072
rect 91612 4060 91618 4072
rect 92017 4063 92075 4069
rect 92017 4060 92029 4063
rect 91612 4032 92029 4060
rect 91612 4020 91618 4032
rect 92017 4029 92029 4032
rect 92063 4029 92075 4063
rect 92017 4023 92075 4029
rect 92106 4020 92112 4072
rect 92164 4060 92170 4072
rect 92661 4063 92719 4069
rect 92661 4060 92673 4063
rect 92164 4032 92673 4060
rect 92164 4020 92170 4032
rect 92661 4029 92673 4032
rect 92707 4029 92719 4063
rect 92661 4023 92719 4029
rect 92750 4020 92756 4072
rect 92808 4060 92814 4072
rect 93305 4063 93363 4069
rect 93305 4060 93317 4063
rect 92808 4032 93317 4060
rect 92808 4020 92814 4032
rect 93305 4029 93317 4032
rect 93351 4029 93363 4063
rect 94130 4060 94136 4072
rect 94091 4032 94136 4060
rect 93305 4023 93363 4029
rect 94130 4020 94136 4032
rect 94188 4020 94194 4072
rect 94774 4060 94780 4072
rect 94735 4032 94780 4060
rect 94774 4020 94780 4032
rect 94832 4020 94838 4072
rect 95970 4060 95976 4072
rect 95931 4032 95976 4060
rect 95970 4020 95976 4032
rect 96028 4020 96034 4072
rect 96908 4060 96936 4088
rect 97184 4069 97212 4100
rect 97445 4097 97457 4100
rect 97491 4097 97503 4131
rect 97445 4091 97503 4097
rect 97169 4063 97227 4069
rect 97169 4060 97181 4063
rect 96908 4032 97181 4060
rect 97169 4029 97181 4032
rect 97215 4029 97227 4063
rect 97169 4023 97227 4029
rect 97353 4063 97411 4069
rect 97353 4029 97365 4063
rect 97399 4060 97411 4063
rect 99282 4060 99288 4072
rect 97399 4032 99288 4060
rect 97399 4029 97411 4032
rect 97353 4023 97411 4029
rect 99282 4020 99288 4032
rect 99340 4020 99346 4072
rect 85448 3964 86172 3992
rect 85448 3952 85454 3964
rect 97442 3952 97448 4004
rect 97500 3992 97506 4004
rect 97629 3995 97687 4001
rect 97629 3992 97641 3995
rect 97500 3964 97641 3992
rect 97500 3952 97506 3964
rect 97629 3961 97641 3964
rect 97675 3992 97687 3995
rect 97905 3995 97963 4001
rect 97905 3992 97917 3995
rect 97675 3964 97917 3992
rect 97675 3961 97687 3964
rect 97629 3955 97687 3961
rect 97905 3961 97917 3964
rect 97951 3961 97963 3995
rect 97905 3955 97963 3961
rect 62356 3896 63172 3924
rect 62356 3884 62362 3896
rect 78214 3884 78220 3936
rect 78272 3924 78278 3936
rect 90174 3924 90180 3936
rect 78272 3896 90180 3924
rect 78272 3884 78278 3896
rect 90174 3884 90180 3896
rect 90232 3884 90238 3936
rect 97994 3924 98000 3936
rect 97955 3896 98000 3924
rect 97994 3884 98000 3896
rect 98052 3884 98058 3936
rect 1104 3834 98808 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 50326 3834
rect 50378 3782 50390 3834
rect 50442 3782 50454 3834
rect 50506 3782 50518 3834
rect 50570 3782 81046 3834
rect 81098 3782 81110 3834
rect 81162 3782 81174 3834
rect 81226 3782 81238 3834
rect 81290 3782 98808 3834
rect 1104 3760 98808 3782
rect 106 3680 112 3732
rect 164 3720 170 3732
rect 1118 3720 1124 3732
rect 164 3692 1124 3720
rect 164 3680 170 3692
rect 1118 3680 1124 3692
rect 1176 3680 1182 3732
rect 2958 3720 2964 3732
rect 2919 3692 2964 3720
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 12069 3723 12127 3729
rect 12069 3689 12081 3723
rect 12115 3720 12127 3723
rect 13354 3720 13360 3732
rect 12115 3692 13360 3720
rect 12115 3689 12127 3692
rect 12069 3683 12127 3689
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 14918 3680 14924 3732
rect 14976 3720 14982 3732
rect 15746 3720 15752 3732
rect 14976 3692 15752 3720
rect 14976 3680 14982 3692
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 68646 3680 68652 3732
rect 68704 3720 68710 3732
rect 85022 3720 85028 3732
rect 68704 3692 84194 3720
rect 84983 3692 85028 3720
rect 68704 3680 68710 3692
rect 2041 3655 2099 3661
rect 2041 3621 2053 3655
rect 2087 3652 2099 3655
rect 4062 3652 4068 3664
rect 2087 3624 4068 3652
rect 2087 3621 2099 3624
rect 2041 3615 2099 3621
rect 4062 3612 4068 3624
rect 4120 3612 4126 3664
rect 5353 3655 5411 3661
rect 5353 3621 5365 3655
rect 5399 3652 5411 3655
rect 6270 3652 6276 3664
rect 5399 3624 6276 3652
rect 5399 3621 5411 3624
rect 5353 3615 5411 3621
rect 6270 3612 6276 3624
rect 6328 3612 6334 3664
rect 6454 3652 6460 3664
rect 6415 3624 6460 3652
rect 6454 3612 6460 3624
rect 6512 3612 6518 3664
rect 7374 3612 7380 3664
rect 7432 3652 7438 3664
rect 7469 3655 7527 3661
rect 7469 3652 7481 3655
rect 7432 3624 7481 3652
rect 7432 3612 7438 3624
rect 7469 3621 7481 3624
rect 7515 3621 7527 3655
rect 7469 3615 7527 3621
rect 8389 3655 8447 3661
rect 8389 3621 8401 3655
rect 8435 3652 8447 3655
rect 8570 3652 8576 3664
rect 8435 3624 8576 3652
rect 8435 3621 8447 3624
rect 8389 3615 8447 3621
rect 8570 3612 8576 3624
rect 8628 3612 8634 3664
rect 9766 3652 9772 3664
rect 9727 3624 9772 3652
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 10689 3655 10747 3661
rect 10689 3621 10701 3655
rect 10735 3652 10747 3655
rect 10778 3652 10784 3664
rect 10735 3624 10784 3652
rect 10735 3621 10747 3624
rect 10689 3615 10747 3621
rect 10778 3612 10784 3624
rect 10836 3612 10842 3664
rect 13262 3652 13268 3664
rect 13223 3624 13268 3652
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 15378 3652 15384 3664
rect 15339 3624 15384 3652
rect 15378 3612 15384 3624
rect 15436 3612 15442 3664
rect 16482 3652 16488 3664
rect 16443 3624 16488 3652
rect 16482 3612 16488 3624
rect 16540 3612 16546 3664
rect 18230 3612 18236 3664
rect 18288 3652 18294 3664
rect 18601 3655 18659 3661
rect 18601 3652 18613 3655
rect 18288 3624 18613 3652
rect 18288 3612 18294 3624
rect 18601 3621 18613 3624
rect 18647 3621 18659 3655
rect 18601 3615 18659 3621
rect 20162 3612 20168 3664
rect 20220 3652 20226 3664
rect 20257 3655 20315 3661
rect 20257 3652 20269 3655
rect 20220 3624 20269 3652
rect 20220 3612 20226 3624
rect 20257 3621 20269 3624
rect 20303 3621 20315 3655
rect 20990 3652 20996 3664
rect 20951 3624 20996 3652
rect 20257 3615 20315 3621
rect 20990 3612 20996 3624
rect 21048 3612 21054 3664
rect 21729 3655 21787 3661
rect 21729 3621 21741 3655
rect 21775 3652 21787 3655
rect 21910 3652 21916 3664
rect 21775 3624 21916 3652
rect 21775 3621 21787 3624
rect 21729 3615 21787 3621
rect 21910 3612 21916 3624
rect 21968 3612 21974 3664
rect 26605 3655 26663 3661
rect 26605 3621 26617 3655
rect 26651 3652 26663 3655
rect 26881 3655 26939 3661
rect 26881 3652 26893 3655
rect 26651 3624 26893 3652
rect 26651 3621 26663 3624
rect 26605 3615 26663 3621
rect 26881 3621 26893 3624
rect 26927 3652 26939 3655
rect 26970 3652 26976 3664
rect 26927 3624 26976 3652
rect 26927 3621 26939 3624
rect 26881 3615 26939 3621
rect 26970 3612 26976 3624
rect 27028 3612 27034 3664
rect 31570 3612 31576 3664
rect 31628 3652 31634 3664
rect 31665 3655 31723 3661
rect 31665 3652 31677 3655
rect 31628 3624 31677 3652
rect 31628 3612 31634 3624
rect 31665 3621 31677 3624
rect 31711 3621 31723 3655
rect 39758 3652 39764 3664
rect 31665 3615 31723 3621
rect 31864 3624 39764 3652
rect 1118 3544 1124 3596
rect 1176 3584 1182 3596
rect 1489 3587 1547 3593
rect 1489 3584 1501 3587
rect 1176 3556 1501 3584
rect 1176 3544 1182 3556
rect 1489 3553 1501 3556
rect 1535 3553 1547 3587
rect 1489 3547 1547 3553
rect 2222 3544 2228 3596
rect 2280 3584 2286 3596
rect 2685 3587 2743 3593
rect 2685 3584 2697 3587
rect 2280 3556 2697 3584
rect 2280 3544 2286 3556
rect 2685 3553 2697 3556
rect 2731 3553 2743 3587
rect 2685 3547 2743 3553
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 4801 3587 4859 3593
rect 4801 3584 4813 3587
rect 4764 3556 4813 3584
rect 4764 3544 4770 3556
rect 4801 3553 4813 3556
rect 4847 3553 4859 3587
rect 4801 3547 4859 3553
rect 5442 3544 5448 3596
rect 5500 3584 5506 3596
rect 5997 3587 6055 3593
rect 5997 3584 6009 3587
rect 5500 3556 6009 3584
rect 5500 3544 5506 3556
rect 5997 3553 6009 3556
rect 6043 3553 6055 3587
rect 7190 3584 7196 3596
rect 7151 3556 7196 3584
rect 5997 3547 6055 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 7742 3544 7748 3596
rect 7800 3584 7806 3596
rect 8113 3587 8171 3593
rect 8113 3584 8125 3587
rect 7800 3556 8125 3584
rect 7800 3544 7806 3556
rect 8113 3553 8125 3556
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 9493 3587 9551 3593
rect 9493 3584 9505 3587
rect 9180 3556 9505 3584
rect 9180 3544 9186 3556
rect 9493 3553 9505 3556
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 10284 3556 10425 3584
rect 10284 3544 10290 3556
rect 10413 3553 10425 3556
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 11793 3587 11851 3593
rect 11793 3553 11805 3587
rect 11839 3584 11851 3587
rect 12066 3584 12072 3596
rect 11839 3556 12072 3584
rect 11839 3553 11851 3556
rect 11793 3547 11851 3553
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 12618 3544 12624 3596
rect 12676 3584 12682 3596
rect 12713 3587 12771 3593
rect 12713 3584 12725 3587
rect 12676 3556 12725 3584
rect 12676 3544 12682 3556
rect 12713 3553 12725 3556
rect 12759 3553 12771 3587
rect 12713 3547 12771 3553
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 14829 3587 14887 3593
rect 14829 3584 14841 3587
rect 14516 3556 14841 3584
rect 14516 3544 14522 3556
rect 14829 3553 14841 3556
rect 14875 3553 14887 3587
rect 14829 3547 14887 3553
rect 15010 3544 15016 3596
rect 15068 3584 15074 3596
rect 16025 3587 16083 3593
rect 16025 3584 16037 3587
rect 15068 3556 16037 3584
rect 15068 3544 15074 3556
rect 16025 3553 16037 3556
rect 16071 3553 16083 3587
rect 16025 3547 16083 3553
rect 16298 3544 16304 3596
rect 16356 3584 16362 3596
rect 17221 3587 17279 3593
rect 17221 3584 17233 3587
rect 16356 3556 17233 3584
rect 16356 3544 16362 3556
rect 17221 3553 17233 3556
rect 17267 3553 17279 3587
rect 17221 3547 17279 3553
rect 18138 3544 18144 3596
rect 18196 3584 18202 3596
rect 18325 3587 18383 3593
rect 18325 3584 18337 3587
rect 18196 3556 18337 3584
rect 18196 3544 18202 3556
rect 18325 3553 18337 3556
rect 18371 3553 18383 3587
rect 19978 3584 19984 3596
rect 19939 3556 19984 3584
rect 18325 3547 18383 3553
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 22186 3544 22192 3596
rect 22244 3584 22250 3596
rect 23017 3587 23075 3593
rect 23017 3584 23029 3587
rect 22244 3556 23029 3584
rect 22244 3544 22250 3556
rect 23017 3553 23029 3556
rect 23063 3553 23075 3587
rect 23017 3547 23075 3553
rect 23474 3544 23480 3596
rect 23532 3584 23538 3596
rect 23661 3587 23719 3593
rect 23661 3584 23673 3587
rect 23532 3556 23673 3584
rect 23532 3544 23538 3556
rect 23661 3553 23673 3556
rect 23707 3553 23719 3587
rect 23661 3547 23719 3553
rect 24670 3544 24676 3596
rect 24728 3584 24734 3596
rect 25225 3587 25283 3593
rect 25225 3584 25237 3587
rect 24728 3556 25237 3584
rect 24728 3544 24734 3556
rect 25225 3553 25237 3556
rect 25271 3553 25283 3587
rect 25225 3547 25283 3553
rect 25869 3587 25927 3593
rect 25869 3553 25881 3587
rect 25915 3553 25927 3587
rect 25869 3547 25927 3553
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3516 17831 3519
rect 21358 3516 21364 3528
rect 17819 3488 21364 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 20806 3408 20812 3460
rect 20864 3448 20870 3460
rect 21913 3451 21971 3457
rect 21913 3448 21925 3451
rect 20864 3420 21925 3448
rect 20864 3408 20870 3420
rect 21913 3417 21925 3420
rect 21959 3417 21971 3451
rect 21913 3411 21971 3417
rect 25222 3408 25228 3460
rect 25280 3448 25286 3460
rect 25884 3448 25912 3547
rect 27062 3544 27068 3596
rect 27120 3584 27126 3596
rect 27433 3587 27491 3593
rect 27433 3584 27445 3587
rect 27120 3556 27445 3584
rect 27120 3544 27126 3556
rect 27433 3553 27445 3556
rect 27479 3553 27491 3587
rect 28074 3584 28080 3596
rect 28035 3556 28080 3584
rect 27433 3547 27491 3553
rect 28074 3544 28080 3556
rect 28132 3544 28138 3596
rect 28902 3584 28908 3596
rect 28863 3556 28908 3584
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 29914 3544 29920 3596
rect 29972 3584 29978 3596
rect 30469 3587 30527 3593
rect 30469 3584 30481 3587
rect 29972 3556 30481 3584
rect 29972 3544 29978 3556
rect 30469 3553 30481 3556
rect 30515 3553 30527 3587
rect 30469 3547 30527 3553
rect 31297 3587 31355 3593
rect 31297 3553 31309 3587
rect 31343 3584 31355 3587
rect 31864 3584 31892 3624
rect 39758 3612 39764 3624
rect 39816 3612 39822 3664
rect 46750 3652 46756 3664
rect 46711 3624 46756 3652
rect 46750 3612 46756 3624
rect 46808 3612 46814 3664
rect 62390 3612 62396 3664
rect 62448 3652 62454 3664
rect 81437 3655 81495 3661
rect 62448 3624 74534 3652
rect 62448 3612 62454 3624
rect 31343 3556 31892 3584
rect 31343 3553 31355 3556
rect 31297 3547 31355 3553
rect 31938 3544 31944 3596
rect 31996 3584 32002 3596
rect 32401 3587 32459 3593
rect 32401 3584 32413 3587
rect 31996 3556 32413 3584
rect 31996 3544 32002 3556
rect 32401 3553 32413 3556
rect 32447 3553 32459 3587
rect 32401 3547 32459 3553
rect 32490 3544 32496 3596
rect 32548 3584 32554 3596
rect 33045 3587 33103 3593
rect 33045 3584 33057 3587
rect 32548 3556 33057 3584
rect 32548 3544 32554 3556
rect 33045 3553 33057 3556
rect 33091 3553 33103 3587
rect 33045 3547 33103 3553
rect 33689 3587 33747 3593
rect 33689 3553 33701 3587
rect 33735 3553 33747 3587
rect 34422 3584 34428 3596
rect 34383 3556 34428 3584
rect 33689 3547 33747 3553
rect 32950 3476 32956 3528
rect 33008 3516 33014 3528
rect 33704 3516 33732 3547
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 35618 3544 35624 3596
rect 35676 3584 35682 3596
rect 35713 3587 35771 3593
rect 35713 3584 35725 3587
rect 35676 3556 35725 3584
rect 35676 3544 35682 3556
rect 35713 3553 35725 3556
rect 35759 3553 35771 3587
rect 36814 3584 36820 3596
rect 36775 3556 36820 3584
rect 35713 3547 35771 3553
rect 36814 3544 36820 3556
rect 36872 3544 36878 3596
rect 37458 3584 37464 3596
rect 37419 3556 37464 3584
rect 37458 3544 37464 3556
rect 37516 3544 37522 3596
rect 38102 3584 38108 3596
rect 38063 3556 38108 3584
rect 38102 3544 38108 3556
rect 38160 3544 38166 3596
rect 39298 3584 39304 3596
rect 39259 3556 39304 3584
rect 39298 3544 39304 3556
rect 39356 3544 39362 3596
rect 40494 3544 40500 3596
rect 40552 3584 40558 3596
rect 40957 3587 41015 3593
rect 40957 3584 40969 3587
rect 40552 3556 40969 3584
rect 40552 3544 40558 3556
rect 40957 3553 40969 3556
rect 41003 3553 41015 3587
rect 41690 3584 41696 3596
rect 41651 3556 41696 3584
rect 40957 3547 41015 3553
rect 41690 3544 41696 3556
rect 41748 3544 41754 3596
rect 42334 3584 42340 3596
rect 42295 3556 42340 3584
rect 42334 3544 42340 3556
rect 42392 3544 42398 3596
rect 42978 3584 42984 3596
rect 42939 3556 42984 3584
rect 42978 3544 42984 3556
rect 43036 3544 43042 3596
rect 43625 3587 43683 3593
rect 43625 3553 43637 3587
rect 43671 3553 43683 3587
rect 44818 3584 44824 3596
rect 44779 3556 44824 3584
rect 43625 3547 43683 3553
rect 33008 3488 33732 3516
rect 33008 3476 33014 3488
rect 42150 3476 42156 3528
rect 42208 3516 42214 3528
rect 43640 3516 43668 3547
rect 44818 3544 44824 3556
rect 44876 3544 44882 3596
rect 46290 3584 46296 3596
rect 46251 3556 46296 3584
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 46566 3544 46572 3596
rect 46624 3584 46630 3596
rect 47397 3587 47455 3593
rect 47397 3584 47409 3587
rect 46624 3556 47409 3584
rect 46624 3544 46630 3556
rect 47397 3553 47409 3556
rect 47443 3553 47455 3587
rect 48041 3587 48099 3593
rect 48041 3584 48053 3587
rect 47397 3547 47455 3553
rect 47504 3556 48053 3584
rect 42208 3488 43668 3516
rect 42208 3476 42214 3488
rect 47210 3476 47216 3528
rect 47268 3516 47274 3528
rect 47504 3516 47532 3556
rect 48041 3553 48053 3556
rect 48087 3553 48099 3587
rect 48041 3547 48099 3553
rect 48685 3587 48743 3593
rect 48685 3553 48697 3587
rect 48731 3553 48743 3587
rect 48685 3547 48743 3553
rect 47268 3488 47532 3516
rect 47268 3476 47274 3488
rect 47854 3476 47860 3528
rect 47912 3516 47918 3528
rect 48700 3516 48728 3547
rect 49050 3544 49056 3596
rect 49108 3584 49114 3596
rect 49329 3587 49387 3593
rect 49329 3584 49341 3587
rect 49108 3556 49341 3584
rect 49108 3544 49114 3556
rect 49329 3553 49341 3556
rect 49375 3553 49387 3587
rect 49329 3547 49387 3553
rect 49694 3544 49700 3596
rect 49752 3584 49758 3596
rect 49973 3587 50031 3593
rect 49973 3584 49985 3587
rect 49752 3556 49985 3584
rect 49752 3544 49758 3556
rect 49973 3553 49985 3556
rect 50019 3553 50031 3587
rect 49973 3547 50031 3553
rect 50890 3544 50896 3596
rect 50948 3584 50954 3596
rect 51445 3587 51503 3593
rect 51445 3584 51457 3587
rect 50948 3556 51457 3584
rect 50948 3544 50954 3556
rect 51445 3553 51457 3556
rect 51491 3553 51503 3587
rect 52086 3584 52092 3596
rect 52047 3556 52092 3584
rect 51445 3547 51503 3553
rect 52086 3544 52092 3556
rect 52144 3544 52150 3596
rect 52730 3584 52736 3596
rect 52691 3556 52736 3584
rect 52730 3544 52736 3556
rect 52788 3544 52794 3596
rect 53282 3544 53288 3596
rect 53340 3584 53346 3596
rect 53377 3587 53435 3593
rect 53377 3584 53389 3587
rect 53340 3556 53389 3584
rect 53340 3544 53346 3556
rect 53377 3553 53389 3556
rect 53423 3553 53435 3587
rect 53377 3547 53435 3553
rect 53926 3544 53932 3596
rect 53984 3584 53990 3596
rect 54021 3587 54079 3593
rect 54021 3584 54033 3587
rect 53984 3556 54033 3584
rect 53984 3544 53990 3556
rect 54021 3553 54033 3556
rect 54067 3553 54079 3587
rect 54021 3547 54079 3553
rect 54570 3544 54576 3596
rect 54628 3584 54634 3596
rect 54665 3587 54723 3593
rect 54665 3584 54677 3587
rect 54628 3556 54677 3584
rect 54628 3544 54634 3556
rect 54665 3553 54677 3556
rect 54711 3553 54723 3587
rect 54665 3547 54723 3553
rect 55122 3544 55128 3596
rect 55180 3584 55186 3596
rect 55309 3587 55367 3593
rect 55309 3584 55321 3587
rect 55180 3556 55321 3584
rect 55180 3544 55186 3556
rect 55309 3553 55321 3556
rect 55355 3553 55367 3587
rect 55309 3547 55367 3553
rect 56318 3544 56324 3596
rect 56376 3584 56382 3596
rect 56689 3587 56747 3593
rect 56689 3584 56701 3587
rect 56376 3556 56701 3584
rect 56376 3544 56382 3556
rect 56689 3553 56701 3556
rect 56735 3553 56747 3587
rect 56689 3547 56747 3553
rect 56962 3544 56968 3596
rect 57020 3584 57026 3596
rect 57333 3587 57391 3593
rect 57333 3584 57345 3587
rect 57020 3556 57345 3584
rect 57020 3544 57026 3556
rect 57333 3553 57345 3556
rect 57379 3553 57391 3587
rect 58158 3584 58164 3596
rect 58119 3556 58164 3584
rect 57333 3547 57391 3553
rect 58158 3544 58164 3556
rect 58216 3544 58222 3596
rect 58802 3584 58808 3596
rect 58763 3556 58808 3584
rect 58802 3544 58808 3556
rect 58860 3544 58866 3596
rect 59449 3587 59507 3593
rect 59449 3553 59461 3587
rect 59495 3553 59507 3587
rect 60642 3584 60648 3596
rect 60603 3556 60648 3584
rect 59449 3547 59507 3553
rect 47912 3488 48728 3516
rect 47912 3476 47918 3488
rect 57974 3476 57980 3528
rect 58032 3516 58038 3528
rect 59464 3516 59492 3547
rect 60642 3544 60648 3556
rect 60700 3544 60706 3596
rect 61286 3544 61292 3596
rect 61344 3584 61350 3596
rect 61933 3587 61991 3593
rect 61933 3584 61945 3587
rect 61344 3556 61945 3584
rect 61344 3544 61350 3556
rect 61933 3553 61945 3556
rect 61979 3553 61991 3587
rect 61933 3547 61991 3553
rect 62577 3587 62635 3593
rect 62577 3553 62589 3587
rect 62623 3553 62635 3587
rect 62577 3547 62635 3553
rect 58032 3488 59492 3516
rect 58032 3476 58038 3488
rect 61838 3476 61844 3528
rect 61896 3516 61902 3528
rect 62592 3516 62620 3547
rect 63034 3544 63040 3596
rect 63092 3584 63098 3596
rect 63221 3587 63279 3593
rect 63221 3584 63233 3587
rect 63092 3556 63233 3584
rect 63092 3544 63098 3556
rect 63221 3553 63233 3556
rect 63267 3553 63279 3587
rect 63221 3547 63279 3553
rect 63678 3544 63684 3596
rect 63736 3584 63742 3596
rect 63865 3587 63923 3593
rect 63865 3584 63877 3587
rect 63736 3556 63877 3584
rect 63736 3544 63742 3556
rect 63865 3553 63877 3556
rect 63911 3553 63923 3587
rect 63865 3547 63923 3553
rect 64322 3544 64328 3596
rect 64380 3584 64386 3596
rect 64509 3587 64567 3593
rect 64509 3584 64521 3587
rect 64380 3556 64521 3584
rect 64380 3544 64386 3556
rect 64509 3553 64521 3556
rect 64555 3553 64567 3587
rect 64509 3547 64567 3553
rect 65153 3587 65211 3593
rect 65153 3553 65165 3587
rect 65199 3553 65211 3587
rect 65153 3547 65211 3553
rect 61896 3488 62620 3516
rect 61896 3476 61902 3488
rect 63494 3476 63500 3528
rect 63552 3516 63558 3528
rect 65168 3516 65196 3547
rect 65334 3544 65340 3596
rect 65392 3584 65398 3596
rect 65797 3587 65855 3593
rect 65797 3584 65809 3587
rect 65392 3556 65809 3584
rect 65392 3544 65398 3556
rect 65797 3553 65809 3556
rect 65843 3553 65855 3587
rect 65797 3547 65855 3553
rect 66806 3544 66812 3596
rect 66864 3584 66870 3596
rect 67177 3587 67235 3593
rect 67177 3584 67189 3587
rect 66864 3556 67189 3584
rect 66864 3544 66870 3556
rect 67177 3553 67189 3556
rect 67223 3553 67235 3587
rect 67910 3584 67916 3596
rect 67871 3556 67916 3584
rect 67177 3547 67235 3553
rect 67910 3544 67916 3556
rect 67968 3544 67974 3596
rect 68554 3584 68560 3596
rect 68515 3556 68560 3584
rect 68554 3544 68560 3556
rect 68612 3544 68618 3596
rect 69198 3584 69204 3596
rect 69159 3556 69204 3584
rect 69198 3544 69204 3556
rect 69256 3544 69262 3596
rect 69750 3544 69756 3596
rect 69808 3584 69814 3596
rect 69845 3587 69903 3593
rect 69845 3584 69857 3587
rect 69808 3556 69857 3584
rect 69808 3544 69814 3556
rect 69845 3553 69857 3556
rect 69891 3553 69903 3587
rect 69845 3547 69903 3553
rect 70394 3544 70400 3596
rect 70452 3584 70458 3596
rect 70489 3587 70547 3593
rect 70489 3584 70501 3587
rect 70452 3556 70501 3584
rect 70452 3544 70458 3556
rect 70489 3553 70501 3556
rect 70535 3553 70547 3587
rect 70489 3547 70547 3553
rect 71133 3587 71191 3593
rect 71133 3553 71145 3587
rect 71179 3553 71191 3587
rect 71133 3547 71191 3553
rect 63552 3488 65196 3516
rect 63552 3476 63558 3488
rect 70210 3476 70216 3528
rect 70268 3516 70274 3528
rect 71148 3516 71176 3547
rect 71590 3544 71596 3596
rect 71648 3584 71654 3596
rect 72421 3587 72479 3593
rect 72421 3584 72433 3587
rect 71648 3556 72433 3584
rect 71648 3544 71654 3556
rect 72421 3553 72433 3556
rect 72467 3553 72479 3587
rect 72421 3547 72479 3553
rect 72786 3544 72792 3596
rect 72844 3584 72850 3596
rect 73065 3587 73123 3593
rect 73065 3584 73077 3587
rect 72844 3556 73077 3584
rect 72844 3544 72850 3556
rect 73065 3553 73077 3556
rect 73111 3553 73123 3587
rect 74074 3584 74080 3596
rect 74035 3556 74080 3584
rect 73065 3547 73123 3553
rect 74074 3544 74080 3556
rect 74132 3544 74138 3596
rect 70268 3488 71176 3516
rect 74506 3516 74534 3624
rect 81437 3621 81449 3655
rect 81483 3652 81495 3655
rect 81526 3652 81532 3664
rect 81483 3624 81532 3652
rect 81483 3621 81495 3624
rect 81437 3615 81495 3621
rect 81526 3612 81532 3624
rect 81584 3652 81590 3664
rect 81713 3655 81771 3661
rect 81713 3652 81725 3655
rect 81584 3624 81725 3652
rect 81584 3612 81590 3624
rect 81713 3621 81725 3624
rect 81759 3621 81771 3655
rect 81713 3615 81771 3621
rect 74626 3544 74632 3596
rect 74684 3584 74690 3596
rect 74721 3587 74779 3593
rect 74721 3584 74733 3587
rect 74684 3556 74733 3584
rect 74684 3544 74690 3556
rect 74721 3553 74733 3556
rect 74767 3553 74779 3587
rect 75914 3584 75920 3596
rect 75875 3556 75920 3584
rect 74721 3547 74779 3553
rect 75914 3544 75920 3556
rect 75972 3544 75978 3596
rect 76466 3544 76472 3596
rect 76524 3584 76530 3596
rect 76561 3587 76619 3593
rect 76561 3584 76573 3587
rect 76524 3556 76573 3584
rect 76524 3544 76530 3556
rect 76561 3553 76573 3556
rect 76607 3553 76619 3587
rect 76561 3547 76619 3553
rect 77110 3544 77116 3596
rect 77168 3584 77174 3596
rect 77665 3587 77723 3593
rect 77665 3584 77677 3587
rect 77168 3556 77677 3584
rect 77168 3544 77174 3556
rect 77665 3553 77677 3556
rect 77711 3553 77723 3587
rect 77665 3547 77723 3553
rect 77754 3544 77760 3596
rect 77812 3584 77818 3596
rect 78309 3587 78367 3593
rect 78309 3584 78321 3587
rect 77812 3556 78321 3584
rect 77812 3544 77818 3556
rect 78309 3553 78321 3556
rect 78355 3553 78367 3587
rect 78309 3547 78367 3553
rect 78398 3544 78404 3596
rect 78456 3584 78462 3596
rect 78953 3587 79011 3593
rect 78953 3584 78965 3587
rect 78456 3556 78965 3584
rect 78456 3544 78462 3556
rect 78953 3553 78965 3556
rect 78999 3553 79011 3587
rect 78953 3547 79011 3553
rect 79042 3544 79048 3596
rect 79100 3584 79106 3596
rect 79597 3587 79655 3593
rect 79597 3584 79609 3587
rect 79100 3556 79609 3584
rect 79100 3544 79106 3556
rect 79597 3553 79609 3556
rect 79643 3553 79655 3587
rect 79597 3547 79655 3553
rect 79686 3544 79692 3596
rect 79744 3584 79750 3596
rect 80241 3587 80299 3593
rect 80241 3584 80253 3587
rect 79744 3556 80253 3584
rect 79744 3544 79750 3556
rect 80241 3553 80253 3556
rect 80287 3553 80299 3587
rect 80241 3547 80299 3553
rect 80885 3587 80943 3593
rect 80885 3553 80897 3587
rect 80931 3553 80943 3587
rect 80885 3547 80943 3553
rect 79962 3516 79968 3528
rect 74506 3488 79968 3516
rect 70268 3476 70274 3488
rect 79962 3476 79968 3488
rect 80020 3476 80026 3528
rect 80146 3476 80152 3528
rect 80204 3516 80210 3528
rect 80900 3516 80928 3547
rect 81618 3544 81624 3596
rect 81676 3584 81682 3596
rect 82909 3587 82967 3593
rect 82909 3584 82921 3587
rect 81676 3556 82921 3584
rect 81676 3544 81682 3556
rect 82909 3553 82921 3556
rect 82955 3553 82967 3587
rect 82909 3547 82967 3553
rect 82998 3544 83004 3596
rect 83056 3584 83062 3596
rect 83553 3587 83611 3593
rect 83553 3584 83565 3587
rect 83056 3556 83565 3584
rect 83056 3544 83062 3556
rect 83553 3553 83565 3556
rect 83599 3553 83611 3587
rect 84166 3584 84194 3692
rect 85022 3680 85028 3692
rect 85080 3680 85086 3732
rect 94866 3720 94872 3732
rect 94827 3692 94872 3720
rect 94866 3680 94872 3692
rect 94924 3720 94930 3732
rect 94924 3692 95188 3720
rect 94924 3680 94930 3692
rect 95160 3661 95188 3692
rect 95145 3655 95203 3661
rect 95145 3621 95157 3655
rect 95191 3621 95203 3655
rect 95145 3615 95203 3621
rect 97353 3655 97411 3661
rect 97353 3621 97365 3655
rect 97399 3652 97411 3655
rect 97629 3655 97687 3661
rect 97629 3652 97641 3655
rect 97399 3624 97641 3652
rect 97399 3621 97411 3624
rect 97353 3615 97411 3621
rect 97629 3621 97641 3624
rect 97675 3652 97687 3655
rect 97718 3652 97724 3664
rect 97675 3624 97724 3652
rect 97675 3621 97687 3624
rect 97629 3615 97687 3621
rect 97718 3612 97724 3624
rect 97776 3612 97782 3664
rect 84381 3587 84439 3593
rect 84381 3584 84393 3587
rect 84166 3556 84393 3584
rect 83553 3547 83611 3553
rect 84381 3553 84393 3556
rect 84427 3553 84439 3587
rect 84381 3547 84439 3553
rect 84470 3544 84476 3596
rect 84528 3593 84534 3596
rect 84528 3587 84587 3593
rect 84528 3553 84541 3587
rect 84575 3553 84587 3587
rect 84654 3584 84660 3596
rect 84615 3556 84660 3584
rect 84528 3547 84587 3553
rect 84528 3544 84534 3547
rect 84654 3544 84660 3556
rect 84712 3544 84718 3596
rect 84746 3544 84752 3596
rect 84804 3584 84810 3596
rect 84930 3584 84936 3596
rect 84804 3556 84849 3584
rect 84891 3556 84936 3584
rect 84804 3544 84810 3556
rect 84930 3544 84936 3556
rect 84988 3544 84994 3596
rect 85022 3544 85028 3596
rect 85080 3584 85086 3596
rect 85577 3587 85635 3593
rect 85577 3584 85589 3587
rect 85080 3556 85589 3584
rect 85080 3544 85086 3556
rect 85577 3553 85589 3556
rect 85623 3553 85635 3587
rect 85577 3547 85635 3553
rect 85666 3544 85672 3596
rect 85724 3584 85730 3596
rect 86221 3587 86279 3593
rect 86221 3584 86233 3587
rect 85724 3556 86233 3584
rect 85724 3544 85730 3556
rect 86221 3553 86233 3556
rect 86267 3553 86279 3587
rect 86221 3547 86279 3553
rect 86865 3587 86923 3593
rect 86865 3553 86877 3587
rect 86911 3553 86923 3587
rect 86865 3547 86923 3553
rect 80204 3488 80928 3516
rect 80992 3488 84194 3516
rect 80204 3476 80210 3488
rect 26694 3448 26700 3460
rect 25280 3420 25912 3448
rect 26655 3420 26700 3448
rect 25280 3408 25286 3420
rect 26694 3408 26700 3420
rect 26752 3408 26758 3460
rect 75178 3408 75184 3460
rect 75236 3448 75242 3460
rect 80992 3448 81020 3488
rect 75236 3420 81020 3448
rect 84166 3448 84194 3488
rect 86034 3476 86040 3528
rect 86092 3516 86098 3528
rect 86880 3516 86908 3547
rect 87966 3544 87972 3596
rect 88024 3584 88030 3596
rect 88153 3587 88211 3593
rect 88153 3584 88165 3587
rect 88024 3556 88165 3584
rect 88024 3544 88030 3556
rect 88153 3553 88165 3556
rect 88199 3553 88211 3587
rect 89254 3584 89260 3596
rect 89215 3556 89260 3584
rect 88153 3547 88211 3553
rect 89254 3544 89260 3556
rect 89312 3544 89318 3596
rect 89898 3584 89904 3596
rect 89859 3556 89904 3584
rect 89898 3544 89904 3556
rect 89956 3544 89962 3596
rect 90542 3584 90548 3596
rect 90503 3556 90548 3584
rect 90542 3544 90548 3556
rect 90600 3544 90606 3596
rect 91094 3544 91100 3596
rect 91152 3584 91158 3596
rect 91189 3587 91247 3593
rect 91189 3584 91201 3587
rect 91152 3556 91201 3584
rect 91152 3544 91158 3556
rect 91189 3553 91201 3556
rect 91235 3553 91247 3587
rect 91189 3547 91247 3553
rect 92293 3587 92351 3593
rect 92293 3553 92305 3587
rect 92339 3584 92351 3587
rect 92382 3584 92388 3596
rect 92339 3556 92388 3584
rect 92339 3553 92351 3556
rect 92293 3547 92351 3553
rect 92382 3544 92388 3556
rect 92440 3544 92446 3596
rect 92934 3544 92940 3596
rect 92992 3584 92998 3596
rect 93397 3587 93455 3593
rect 93397 3584 93409 3587
rect 92992 3556 93409 3584
rect 92992 3544 92998 3556
rect 93397 3553 93409 3556
rect 93443 3553 93455 3587
rect 93397 3547 93455 3553
rect 93578 3544 93584 3596
rect 93636 3584 93642 3596
rect 94041 3587 94099 3593
rect 94041 3584 94053 3587
rect 93636 3556 94053 3584
rect 93636 3544 93642 3556
rect 94041 3553 94053 3556
rect 94087 3553 94099 3587
rect 94041 3547 94099 3553
rect 95418 3544 95424 3596
rect 95476 3584 95482 3596
rect 95697 3587 95755 3593
rect 95697 3584 95709 3587
rect 95476 3556 95709 3584
rect 95476 3544 95482 3556
rect 95697 3553 95709 3556
rect 95743 3553 95755 3587
rect 96801 3587 96859 3593
rect 96801 3584 96813 3587
rect 95697 3547 95755 3553
rect 96632 3556 96813 3584
rect 86092 3488 86908 3516
rect 86092 3476 86098 3488
rect 94498 3476 94504 3528
rect 94556 3516 94562 3528
rect 96632 3525 96660 3556
rect 96801 3553 96813 3556
rect 96847 3584 96859 3587
rect 97077 3587 97135 3593
rect 97077 3584 97089 3587
rect 96847 3556 97089 3584
rect 96847 3553 96859 3556
rect 96801 3547 96859 3553
rect 97077 3553 97089 3556
rect 97123 3553 97135 3587
rect 97077 3547 97135 3553
rect 96617 3519 96675 3525
rect 96617 3516 96629 3519
rect 94556 3488 96629 3516
rect 94556 3476 94562 3488
rect 96617 3485 96629 3488
rect 96663 3485 96675 3519
rect 96617 3479 96675 3485
rect 96985 3519 97043 3525
rect 96985 3485 96997 3519
rect 97031 3516 97043 3519
rect 98638 3516 98644 3528
rect 97031 3488 98644 3516
rect 97031 3485 97043 3488
rect 96985 3479 97043 3485
rect 98638 3476 98644 3488
rect 98696 3476 98702 3528
rect 88702 3448 88708 3460
rect 84166 3420 88708 3448
rect 75236 3408 75242 3420
rect 88702 3408 88708 3420
rect 88760 3408 88766 3460
rect 94958 3448 94964 3460
rect 94919 3420 94964 3448
rect 94958 3408 94964 3420
rect 95016 3408 95022 3460
rect 97442 3448 97448 3460
rect 97403 3420 97448 3448
rect 97442 3408 97448 3420
rect 97500 3408 97506 3460
rect 20162 3340 20168 3392
rect 20220 3380 20226 3392
rect 21085 3383 21143 3389
rect 21085 3380 21097 3383
rect 20220 3352 21097 3380
rect 20220 3340 20226 3352
rect 21085 3349 21097 3352
rect 21131 3349 21143 3383
rect 21085 3343 21143 3349
rect 22557 3383 22615 3389
rect 22557 3349 22569 3383
rect 22603 3380 22615 3383
rect 26326 3380 26332 3392
rect 22603 3352 26332 3380
rect 22603 3349 22615 3352
rect 22557 3343 22615 3349
rect 26326 3340 26332 3352
rect 26384 3340 26390 3392
rect 81621 3383 81679 3389
rect 81621 3349 81633 3383
rect 81667 3380 81679 3383
rect 81710 3380 81716 3392
rect 81667 3352 81716 3380
rect 81667 3349 81679 3352
rect 81621 3343 81679 3349
rect 81710 3340 81716 3352
rect 81768 3340 81774 3392
rect 84286 3380 84292 3392
rect 84247 3352 84292 3380
rect 84286 3340 84292 3352
rect 84344 3340 84350 3392
rect 1104 3290 98808 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 65686 3290
rect 65738 3238 65750 3290
rect 65802 3238 65814 3290
rect 65866 3238 65878 3290
rect 65930 3238 96406 3290
rect 96458 3238 96470 3290
rect 96522 3238 96534 3290
rect 96586 3238 96598 3290
rect 96650 3238 98808 3290
rect 1104 3216 98808 3238
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 9306 3176 9312 3188
rect 7239 3148 9312 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 18966 3176 18972 3188
rect 13740 3148 18972 3176
rect 13354 3068 13360 3120
rect 13412 3108 13418 3120
rect 13412 3080 13676 3108
rect 13412 3068 13418 3080
rect 2406 3040 2412 3052
rect 2367 3012 2412 3040
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3040 5319 3043
rect 8754 3040 8760 3052
rect 5307 3012 8760 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 10962 3040 10968 3052
rect 10923 3012 10968 3040
rect 10962 3000 10968 3012
rect 11020 3000 11026 3052
rect 12710 3000 12716 3052
rect 12768 3040 12774 3052
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 12768 3012 12817 3040
rect 12768 3000 12774 3012
rect 12805 3009 12817 3012
rect 12851 3009 12863 3043
rect 12805 3003 12863 3009
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2972 2099 2975
rect 2866 2972 2872 2984
rect 2087 2944 2872 2972
rect 2087 2941 2099 2944
rect 2041 2935 2099 2941
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 3142 2972 3148 2984
rect 3103 2944 3148 2972
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 3694 2932 3700 2984
rect 3752 2972 3758 2984
rect 4709 2975 4767 2981
rect 4709 2972 4721 2975
rect 3752 2944 4721 2972
rect 3752 2932 3758 2944
rect 4709 2941 4721 2944
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2972 7803 2975
rect 8202 2972 8208 2984
rect 7791 2944 8208 2972
rect 7791 2941 7803 2944
rect 7745 2935 7803 2941
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 8444 2944 8493 2972
rect 8444 2932 8450 2944
rect 8481 2941 8493 2944
rect 8527 2941 8539 2975
rect 8481 2935 8539 2941
rect 8662 2932 8668 2984
rect 8720 2972 8726 2984
rect 8849 2975 8907 2981
rect 8849 2972 8861 2975
rect 8720 2944 8861 2972
rect 8720 2932 8726 2944
rect 8849 2941 8861 2944
rect 8895 2941 8907 2975
rect 8849 2935 8907 2941
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2972 9735 2975
rect 9858 2972 9864 2984
rect 9723 2944 9864 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 10870 2972 10876 2984
rect 10551 2944 10876 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 13170 2932 13176 2984
rect 13228 2972 13234 2984
rect 13648 2981 13676 3080
rect 13740 3049 13768 3148
rect 18966 3136 18972 3148
rect 19024 3136 19030 3188
rect 25314 3176 25320 3188
rect 25275 3148 25320 3176
rect 25314 3136 25320 3148
rect 25372 3136 25378 3188
rect 27709 3179 27767 3185
rect 27709 3145 27721 3179
rect 27755 3176 27767 3179
rect 27798 3176 27804 3188
rect 27755 3148 27804 3176
rect 27755 3145 27767 3148
rect 27709 3139 27767 3145
rect 27798 3136 27804 3148
rect 27856 3136 27862 3188
rect 38194 3176 38200 3188
rect 38155 3148 38200 3176
rect 38194 3136 38200 3148
rect 38252 3136 38258 3188
rect 47302 3176 47308 3188
rect 47263 3148 47308 3176
rect 47302 3136 47308 3148
rect 47360 3136 47366 3188
rect 55214 3136 55220 3188
rect 55272 3176 55278 3188
rect 62482 3176 62488 3188
rect 55272 3148 55317 3176
rect 62443 3148 62488 3176
rect 55272 3136 55278 3148
rect 62482 3136 62488 3148
rect 62540 3136 62546 3188
rect 66714 3176 66720 3188
rect 66675 3148 66720 3176
rect 66714 3136 66720 3148
rect 66772 3136 66778 3188
rect 72234 3176 72240 3188
rect 72195 3148 72240 3176
rect 72234 3136 72240 3148
rect 72292 3136 72298 3188
rect 80149 3179 80207 3185
rect 80149 3145 80161 3179
rect 80195 3176 80207 3179
rect 80238 3176 80244 3188
rect 80195 3148 80244 3176
rect 80195 3145 80207 3148
rect 80149 3139 80207 3145
rect 80238 3136 80244 3148
rect 80296 3136 80302 3188
rect 80882 3136 80888 3188
rect 80940 3176 80946 3188
rect 81897 3179 81955 3185
rect 81897 3176 81909 3179
rect 80940 3148 81909 3176
rect 80940 3136 80946 3148
rect 81897 3145 81909 3148
rect 81943 3145 81955 3179
rect 81897 3139 81955 3145
rect 90637 3179 90695 3185
rect 90637 3145 90649 3179
rect 90683 3176 90695 3179
rect 90818 3176 90824 3188
rect 90683 3148 90824 3176
rect 90683 3145 90695 3148
rect 90637 3139 90695 3145
rect 90818 3136 90824 3148
rect 90876 3136 90882 3188
rect 91278 3176 91284 3188
rect 91239 3148 91284 3176
rect 91278 3136 91284 3148
rect 91336 3136 91342 3188
rect 93670 3176 93676 3188
rect 93631 3148 93676 3176
rect 93670 3136 93676 3148
rect 93728 3136 93734 3188
rect 95878 3136 95884 3188
rect 95936 3176 95942 3188
rect 96617 3179 96675 3185
rect 96617 3176 96629 3179
rect 95936 3148 96629 3176
rect 95936 3136 95942 3148
rect 96617 3145 96629 3148
rect 96663 3176 96675 3179
rect 97077 3179 97135 3185
rect 97077 3176 97089 3179
rect 96663 3148 97089 3176
rect 96663 3145 96675 3148
rect 96617 3139 96675 3145
rect 97077 3145 97089 3148
rect 97123 3176 97135 3179
rect 97261 3179 97319 3185
rect 97261 3176 97273 3179
rect 97123 3148 97273 3176
rect 97123 3145 97135 3148
rect 97077 3139 97135 3145
rect 97261 3145 97273 3148
rect 97307 3145 97319 3179
rect 97261 3139 97319 3145
rect 14090 3068 14096 3120
rect 14148 3108 14154 3120
rect 15841 3111 15899 3117
rect 15841 3108 15853 3111
rect 14148 3080 15853 3108
rect 14148 3068 14154 3080
rect 15841 3077 15853 3080
rect 15887 3077 15899 3111
rect 15841 3071 15899 3077
rect 35802 3068 35808 3120
rect 35860 3108 35866 3120
rect 38930 3108 38936 3120
rect 35860 3080 38936 3108
rect 35860 3068 35866 3080
rect 38930 3068 38936 3080
rect 38988 3068 38994 3120
rect 57146 3068 57152 3120
rect 57204 3108 57210 3120
rect 59354 3108 59360 3120
rect 57204 3080 59360 3108
rect 57204 3068 57210 3080
rect 59354 3068 59360 3080
rect 59412 3068 59418 3120
rect 62206 3068 62212 3120
rect 62264 3108 62270 3120
rect 85114 3108 85120 3120
rect 62264 3080 67772 3108
rect 62264 3068 62270 3080
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 13817 3043 13875 3049
rect 13817 3009 13829 3043
rect 13863 3040 13875 3043
rect 13906 3040 13912 3052
rect 13863 3012 13912 3040
rect 13863 3009 13875 3012
rect 13817 3003 13875 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14182 3040 14188 3052
rect 14143 3012 14188 3040
rect 14182 3000 14188 3012
rect 14240 3000 14246 3052
rect 15102 3040 15108 3052
rect 15063 3012 15108 3040
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 17034 3000 17040 3052
rect 17092 3040 17098 3052
rect 17681 3043 17739 3049
rect 17681 3040 17693 3043
rect 17092 3012 17693 3040
rect 17092 3000 17098 3012
rect 17681 3009 17693 3012
rect 17727 3009 17739 3043
rect 19242 3040 19248 3052
rect 19203 3012 19248 3040
rect 17681 3003 17739 3009
rect 19242 3000 19248 3012
rect 19300 3000 19306 3052
rect 20254 3000 20260 3052
rect 20312 3040 20318 3052
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 20312 3012 20361 3040
rect 20312 3000 20318 3012
rect 20349 3009 20361 3012
rect 20395 3009 20407 3043
rect 20349 3003 20407 3009
rect 20622 3000 20628 3052
rect 20680 3000 20686 3052
rect 21450 3040 21456 3052
rect 21411 3012 21456 3040
rect 21450 3000 21456 3012
rect 21508 3000 21514 3052
rect 43530 3000 43536 3052
rect 43588 3040 43594 3052
rect 50617 3043 50675 3049
rect 43588 3012 44312 3040
rect 43588 3000 43594 3012
rect 13449 2975 13507 2981
rect 13449 2972 13461 2975
rect 13228 2944 13461 2972
rect 13228 2932 13234 2944
rect 13449 2941 13461 2944
rect 13495 2941 13507 2975
rect 13449 2935 13507 2941
rect 13632 2975 13690 2981
rect 13632 2941 13644 2975
rect 13678 2941 13690 2975
rect 13998 2972 14004 2984
rect 13959 2944 14004 2972
rect 13632 2935 13690 2941
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 3970 2904 3976 2916
rect 3931 2876 3976 2904
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 5994 2864 6000 2916
rect 6052 2904 6058 2916
rect 6917 2907 6975 2913
rect 6917 2904 6929 2907
rect 6052 2876 6929 2904
rect 6052 2864 6058 2876
rect 6917 2873 6929 2876
rect 6963 2873 6975 2907
rect 6917 2867 6975 2873
rect 11422 2864 11428 2916
rect 11480 2904 11486 2916
rect 12069 2907 12127 2913
rect 12069 2904 12081 2907
rect 11480 2876 12081 2904
rect 11480 2864 11486 2876
rect 12069 2873 12081 2876
rect 12115 2873 12127 2907
rect 12069 2867 12127 2873
rect 13906 2864 13912 2916
rect 13964 2904 13970 2916
rect 14752 2904 14780 2935
rect 15746 2932 15752 2984
rect 15804 2972 15810 2984
rect 17405 2975 17463 2981
rect 17405 2972 17417 2975
rect 15804 2944 17417 2972
rect 15804 2932 15810 2944
rect 17405 2941 17417 2944
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 18782 2932 18788 2984
rect 18840 2972 18846 2984
rect 18877 2975 18935 2981
rect 18877 2972 18889 2975
rect 18840 2944 18889 2972
rect 18840 2932 18846 2944
rect 18877 2941 18889 2944
rect 18923 2941 18935 2975
rect 18877 2935 18935 2941
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 20073 2975 20131 2981
rect 20073 2972 20085 2975
rect 19392 2944 20085 2972
rect 19392 2932 19398 2944
rect 20073 2941 20085 2944
rect 20119 2941 20131 2975
rect 20640 2972 20668 3000
rect 21177 2975 21235 2981
rect 21177 2972 21189 2975
rect 20640 2944 21189 2972
rect 20073 2935 20131 2941
rect 21177 2941 21189 2944
rect 21223 2941 21235 2975
rect 22646 2972 22652 2984
rect 22607 2944 22652 2972
rect 21177 2935 21235 2941
rect 22646 2932 22652 2944
rect 22704 2932 22710 2984
rect 23293 2975 23351 2981
rect 23293 2972 23305 2975
rect 22756 2944 23305 2972
rect 13964 2876 14780 2904
rect 15657 2907 15715 2913
rect 13964 2864 13970 2876
rect 15657 2873 15669 2907
rect 15703 2904 15715 2907
rect 16025 2907 16083 2913
rect 16025 2904 16037 2907
rect 15703 2876 16037 2904
rect 15703 2873 15715 2876
rect 15657 2867 15715 2873
rect 16025 2873 16037 2876
rect 16071 2904 16083 2907
rect 16206 2904 16212 2916
rect 16071 2876 16212 2904
rect 16071 2873 16083 2876
rect 16025 2867 16083 2873
rect 16206 2864 16212 2876
rect 16264 2864 16270 2916
rect 19242 2864 19248 2916
rect 19300 2904 19306 2916
rect 19426 2904 19432 2916
rect 19300 2876 19432 2904
rect 19300 2864 19306 2876
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 21634 2864 21640 2916
rect 21692 2904 21698 2916
rect 22756 2904 22784 2944
rect 23293 2941 23305 2944
rect 23339 2941 23351 2975
rect 23293 2935 23351 2941
rect 23937 2975 23995 2981
rect 23937 2941 23949 2975
rect 23983 2941 23995 2975
rect 23937 2935 23995 2941
rect 21692 2876 22784 2904
rect 21692 2864 21698 2876
rect 22922 2864 22928 2916
rect 22980 2904 22986 2916
rect 23952 2904 23980 2935
rect 24026 2932 24032 2984
rect 24084 2972 24090 2984
rect 24581 2975 24639 2981
rect 24581 2972 24593 2975
rect 24084 2944 24593 2972
rect 24084 2932 24090 2944
rect 24581 2941 24593 2944
rect 24627 2941 24639 2975
rect 24581 2935 24639 2941
rect 25314 2932 25320 2984
rect 25372 2972 25378 2984
rect 25685 2975 25743 2981
rect 25685 2972 25697 2975
rect 25372 2944 25697 2972
rect 25372 2932 25378 2944
rect 25685 2941 25697 2944
rect 25731 2941 25743 2975
rect 26326 2972 26332 2984
rect 26287 2944 26332 2972
rect 25685 2935 25743 2941
rect 26326 2932 26332 2944
rect 26384 2932 26390 2984
rect 27798 2932 27804 2984
rect 27856 2972 27862 2984
rect 27985 2975 28043 2981
rect 27985 2972 27997 2975
rect 27856 2944 27997 2972
rect 27856 2932 27862 2944
rect 27985 2941 27997 2944
rect 28031 2941 28043 2975
rect 27985 2935 28043 2941
rect 28537 2975 28595 2981
rect 28537 2941 28549 2975
rect 28583 2941 28595 2975
rect 28537 2935 28595 2941
rect 29181 2975 29239 2981
rect 29181 2941 29193 2975
rect 29227 2941 29239 2975
rect 29181 2935 29239 2941
rect 25498 2904 25504 2916
rect 22980 2876 23980 2904
rect 25459 2876 25504 2904
rect 22980 2864 22986 2876
rect 25498 2864 25504 2876
rect 25556 2864 25562 2916
rect 27706 2864 27712 2916
rect 27764 2904 27770 2916
rect 28552 2904 28580 2935
rect 27764 2876 28580 2904
rect 27764 2864 27770 2876
rect 9214 2796 9220 2848
rect 9272 2836 9278 2848
rect 9769 2839 9827 2845
rect 9769 2836 9781 2839
rect 9272 2808 9781 2836
rect 9272 2796 9278 2808
rect 9769 2805 9781 2808
rect 9815 2805 9827 2839
rect 9769 2799 9827 2805
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 12526 2836 12532 2848
rect 11296 2808 12532 2836
rect 11296 2796 11302 2808
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 21358 2796 21364 2848
rect 21416 2836 21422 2848
rect 22741 2839 22799 2845
rect 22741 2836 22753 2839
rect 21416 2808 22753 2836
rect 21416 2796 21422 2808
rect 22741 2805 22753 2808
rect 22787 2805 22799 2839
rect 22741 2799 22799 2805
rect 26050 2796 26056 2848
rect 26108 2836 26114 2848
rect 26421 2839 26479 2845
rect 26421 2836 26433 2839
rect 26108 2808 26433 2836
rect 26108 2796 26114 2808
rect 26421 2805 26433 2808
rect 26467 2805 26479 2839
rect 26421 2799 26479 2805
rect 27338 2796 27344 2848
rect 27396 2836 27402 2848
rect 27893 2839 27951 2845
rect 27893 2836 27905 2839
rect 27396 2808 27905 2836
rect 27396 2796 27402 2808
rect 27893 2805 27905 2808
rect 27939 2805 27951 2839
rect 27893 2799 27951 2805
rect 28350 2796 28356 2848
rect 28408 2836 28414 2848
rect 29196 2836 29224 2935
rect 29546 2932 29552 2984
rect 29604 2972 29610 2984
rect 29825 2975 29883 2981
rect 29825 2972 29837 2975
rect 29604 2944 29837 2972
rect 29604 2932 29610 2944
rect 29825 2941 29837 2944
rect 29871 2941 29883 2975
rect 29825 2935 29883 2941
rect 30098 2932 30104 2984
rect 30156 2972 30162 2984
rect 30469 2975 30527 2981
rect 30469 2972 30481 2975
rect 30156 2944 30481 2972
rect 30156 2932 30162 2944
rect 30469 2941 30481 2944
rect 30515 2941 30527 2975
rect 30469 2935 30527 2941
rect 30742 2932 30748 2984
rect 30800 2972 30806 2984
rect 31113 2975 31171 2981
rect 31113 2972 31125 2975
rect 30800 2944 31125 2972
rect 30800 2932 30806 2944
rect 31113 2941 31125 2944
rect 31159 2941 31171 2975
rect 31113 2935 31171 2941
rect 31386 2932 31392 2984
rect 31444 2972 31450 2984
rect 31757 2975 31815 2981
rect 31757 2972 31769 2975
rect 31444 2944 31769 2972
rect 31444 2932 31450 2944
rect 31757 2941 31769 2944
rect 31803 2941 31815 2975
rect 31757 2935 31815 2941
rect 32582 2932 32588 2984
rect 32640 2972 32646 2984
rect 33045 2975 33103 2981
rect 33045 2972 33057 2975
rect 32640 2944 33057 2972
rect 32640 2932 32646 2944
rect 33045 2941 33057 2944
rect 33091 2941 33103 2975
rect 33045 2935 33103 2941
rect 33226 2932 33232 2984
rect 33284 2972 33290 2984
rect 33689 2975 33747 2981
rect 33689 2972 33701 2975
rect 33284 2944 33701 2972
rect 33284 2932 33290 2944
rect 33689 2941 33701 2944
rect 33735 2941 33747 2975
rect 33689 2935 33747 2941
rect 33778 2932 33784 2984
rect 33836 2972 33842 2984
rect 34333 2975 34391 2981
rect 34333 2972 34345 2975
rect 33836 2944 34345 2972
rect 33836 2932 33842 2944
rect 34333 2941 34345 2944
rect 34379 2941 34391 2975
rect 34333 2935 34391 2941
rect 35161 2975 35219 2981
rect 35161 2941 35173 2975
rect 35207 2972 35219 2975
rect 35437 2975 35495 2981
rect 35437 2972 35449 2975
rect 35207 2944 35449 2972
rect 35207 2941 35219 2944
rect 35161 2935 35219 2941
rect 35437 2941 35449 2944
rect 35483 2972 35495 2975
rect 35526 2972 35532 2984
rect 35483 2944 35532 2972
rect 35483 2941 35495 2944
rect 35437 2935 35495 2941
rect 35526 2932 35532 2944
rect 35584 2932 35590 2984
rect 35989 2975 36047 2981
rect 35989 2972 36001 2975
rect 35866 2944 36001 2972
rect 35250 2904 35256 2916
rect 35211 2876 35256 2904
rect 35250 2864 35256 2876
rect 35308 2864 35314 2916
rect 35342 2864 35348 2916
rect 35400 2904 35406 2916
rect 35866 2904 35894 2944
rect 35989 2941 36001 2944
rect 36035 2941 36047 2975
rect 35989 2935 36047 2941
rect 36262 2932 36268 2984
rect 36320 2972 36326 2984
rect 36633 2975 36691 2981
rect 36633 2972 36645 2975
rect 36320 2944 36645 2972
rect 36320 2932 36326 2944
rect 36633 2941 36645 2944
rect 36679 2941 36691 2975
rect 36633 2935 36691 2941
rect 38194 2932 38200 2984
rect 38252 2972 38258 2984
rect 38473 2975 38531 2981
rect 38473 2972 38485 2975
rect 38252 2944 38485 2972
rect 38252 2932 38258 2944
rect 38473 2941 38485 2944
rect 38519 2941 38531 2975
rect 38473 2935 38531 2941
rect 38654 2932 38660 2984
rect 38712 2972 38718 2984
rect 39025 2975 39083 2981
rect 39025 2972 39037 2975
rect 38712 2944 39037 2972
rect 38712 2932 38718 2944
rect 39025 2941 39037 2944
rect 39071 2941 39083 2975
rect 40218 2972 40224 2984
rect 40179 2944 40224 2972
rect 39025 2935 39083 2941
rect 40218 2932 40224 2944
rect 40276 2932 40282 2984
rect 41233 2975 41291 2981
rect 41233 2941 41245 2975
rect 41279 2972 41291 2975
rect 41509 2975 41567 2981
rect 41509 2972 41521 2975
rect 41279 2944 41521 2972
rect 41279 2941 41291 2944
rect 41233 2935 41291 2941
rect 41509 2941 41521 2944
rect 41555 2972 41567 2975
rect 41598 2972 41604 2984
rect 41555 2944 41604 2972
rect 41555 2941 41567 2944
rect 41509 2935 41567 2941
rect 41598 2932 41604 2944
rect 41656 2932 41662 2984
rect 42061 2975 42119 2981
rect 42061 2941 42073 2975
rect 42107 2941 42119 2975
rect 42061 2935 42119 2941
rect 43441 2975 43499 2981
rect 43441 2941 43453 2975
rect 43487 2972 43499 2975
rect 43714 2972 43720 2984
rect 43487 2944 43720 2972
rect 43487 2941 43499 2944
rect 43441 2935 43499 2941
rect 35400 2876 35894 2904
rect 35400 2864 35406 2876
rect 37642 2864 37648 2916
rect 37700 2904 37706 2916
rect 38289 2907 38347 2913
rect 38289 2904 38301 2907
rect 37700 2876 38301 2904
rect 37700 2864 37706 2876
rect 38289 2873 38301 2876
rect 38335 2873 38347 2907
rect 41322 2904 41328 2916
rect 41283 2876 41328 2904
rect 38289 2867 38347 2873
rect 41322 2864 41328 2876
rect 41380 2864 41386 2916
rect 28408 2808 29224 2836
rect 28408 2796 28414 2808
rect 37090 2796 37096 2848
rect 37148 2836 37154 2848
rect 38746 2836 38752 2848
rect 37148 2808 38752 2836
rect 37148 2796 37154 2808
rect 38746 2796 38752 2808
rect 38804 2796 38810 2848
rect 40126 2796 40132 2848
rect 40184 2836 40190 2848
rect 40313 2839 40371 2845
rect 40313 2836 40325 2839
rect 40184 2808 40325 2836
rect 40184 2796 40190 2808
rect 40313 2805 40325 2808
rect 40359 2805 40371 2839
rect 40313 2799 40371 2805
rect 41138 2796 41144 2848
rect 41196 2836 41202 2848
rect 42076 2836 42104 2935
rect 43714 2932 43720 2944
rect 43772 2932 43778 2984
rect 44284 2981 44312 3012
rect 50617 3009 50629 3043
rect 50663 3040 50675 3043
rect 52362 3040 52368 3052
rect 50663 3012 52368 3040
rect 50663 3009 50675 3012
rect 50617 3003 50675 3009
rect 52362 3000 52368 3012
rect 52420 3000 52426 3052
rect 54846 3000 54852 3052
rect 54904 3040 54910 3052
rect 58342 3040 58348 3052
rect 54904 3012 58348 3040
rect 54904 3000 54910 3012
rect 58342 3000 58348 3012
rect 58400 3000 58406 3052
rect 58434 3000 58440 3052
rect 58492 3040 58498 3052
rect 61562 3040 61568 3052
rect 58492 3012 61568 3040
rect 58492 3000 58498 3012
rect 61562 3000 61568 3012
rect 61620 3000 61626 3052
rect 66162 3000 66168 3052
rect 66220 3040 66226 3052
rect 67744 3040 67772 3080
rect 79152 3080 85120 3108
rect 70397 3043 70455 3049
rect 70397 3040 70409 3043
rect 66220 3012 67680 3040
rect 67744 3012 70409 3040
rect 66220 3000 66226 3012
rect 44269 2975 44327 2981
rect 44269 2941 44281 2975
rect 44315 2941 44327 2975
rect 44269 2935 44327 2941
rect 44913 2975 44971 2981
rect 44913 2941 44925 2975
rect 44959 2941 44971 2975
rect 44913 2935 44971 2941
rect 45465 2975 45523 2981
rect 45465 2941 45477 2975
rect 45511 2972 45523 2975
rect 45738 2972 45744 2984
rect 45511 2944 45744 2972
rect 45511 2941 45523 2944
rect 45465 2935 45523 2941
rect 43162 2864 43168 2916
rect 43220 2904 43226 2916
rect 43533 2907 43591 2913
rect 43533 2904 43545 2907
rect 43220 2876 43545 2904
rect 43220 2864 43226 2876
rect 43533 2873 43545 2876
rect 43579 2873 43591 2907
rect 43533 2867 43591 2873
rect 44174 2864 44180 2916
rect 44232 2904 44238 2916
rect 44928 2904 44956 2935
rect 45738 2932 45744 2944
rect 45796 2932 45802 2984
rect 46293 2975 46351 2981
rect 46293 2941 46305 2975
rect 46339 2941 46351 2975
rect 46293 2935 46351 2941
rect 44232 2876 44956 2904
rect 44232 2864 44238 2876
rect 45554 2864 45560 2916
rect 45612 2904 45618 2916
rect 45612 2876 45657 2904
rect 45612 2864 45618 2876
rect 41196 2808 42104 2836
rect 41196 2796 41202 2808
rect 45370 2796 45376 2848
rect 45428 2836 45434 2848
rect 46308 2836 46336 2935
rect 47302 2932 47308 2984
rect 47360 2972 47366 2984
rect 47581 2975 47639 2981
rect 47581 2972 47593 2975
rect 47360 2944 47593 2972
rect 47360 2932 47366 2944
rect 47581 2941 47593 2944
rect 47627 2941 47639 2975
rect 47581 2935 47639 2941
rect 49145 2975 49203 2981
rect 49145 2941 49157 2975
rect 49191 2972 49203 2975
rect 49421 2975 49479 2981
rect 49421 2972 49433 2975
rect 49191 2944 49433 2972
rect 49191 2941 49203 2944
rect 49145 2935 49203 2941
rect 49421 2941 49433 2944
rect 49467 2972 49479 2975
rect 49510 2972 49516 2984
rect 49467 2944 49516 2972
rect 49467 2941 49479 2944
rect 49421 2935 49479 2941
rect 49510 2932 49516 2944
rect 49568 2932 49574 2984
rect 50985 2975 51043 2981
rect 50985 2941 50997 2975
rect 51031 2972 51043 2975
rect 51258 2972 51264 2984
rect 51031 2944 51264 2972
rect 51031 2941 51043 2944
rect 50985 2935 51043 2941
rect 51258 2932 51264 2944
rect 51316 2932 51322 2984
rect 51813 2975 51871 2981
rect 51813 2972 51825 2975
rect 51368 2944 51825 2972
rect 47394 2904 47400 2916
rect 47355 2876 47400 2904
rect 47394 2864 47400 2876
rect 47452 2864 47458 2916
rect 49234 2904 49240 2916
rect 49195 2876 49240 2904
rect 49234 2864 49240 2876
rect 49292 2864 49298 2916
rect 51074 2904 51080 2916
rect 51035 2876 51080 2904
rect 51074 2864 51080 2876
rect 51132 2864 51138 2916
rect 45428 2808 46336 2836
rect 45428 2796 45434 2808
rect 50154 2796 50160 2848
rect 50212 2836 50218 2848
rect 51368 2836 51396 2944
rect 51813 2941 51825 2944
rect 51859 2941 51871 2975
rect 51813 2935 51871 2941
rect 52457 2975 52515 2981
rect 52457 2941 52469 2975
rect 52503 2941 52515 2975
rect 54110 2972 54116 2984
rect 54071 2944 54116 2972
rect 52457 2935 52515 2941
rect 51442 2864 51448 2916
rect 51500 2904 51506 2916
rect 52472 2904 52500 2935
rect 54110 2932 54116 2944
rect 54168 2932 54174 2984
rect 55214 2932 55220 2984
rect 55272 2972 55278 2984
rect 55493 2975 55551 2981
rect 55493 2972 55505 2975
rect 55272 2944 55505 2972
rect 55272 2932 55278 2944
rect 55493 2941 55505 2944
rect 55539 2941 55551 2975
rect 55493 2935 55551 2941
rect 56505 2975 56563 2981
rect 56505 2941 56517 2975
rect 56551 2972 56563 2975
rect 56781 2975 56839 2981
rect 56781 2972 56793 2975
rect 56551 2944 56793 2972
rect 56551 2941 56563 2944
rect 56505 2935 56563 2941
rect 56781 2941 56793 2944
rect 56827 2972 56839 2975
rect 56870 2972 56876 2984
rect 56827 2944 56876 2972
rect 56827 2941 56839 2944
rect 56781 2935 56839 2941
rect 56870 2932 56876 2944
rect 56928 2932 56934 2984
rect 57333 2975 57391 2981
rect 57333 2941 57345 2975
rect 57379 2941 57391 2975
rect 57333 2935 57391 2941
rect 55306 2904 55312 2916
rect 51500 2876 52500 2904
rect 55267 2876 55312 2904
rect 51500 2864 51506 2876
rect 55306 2864 55312 2876
rect 55364 2864 55370 2916
rect 56594 2904 56600 2916
rect 56555 2876 56600 2904
rect 56594 2864 56600 2876
rect 56652 2864 56658 2916
rect 50212 2808 51396 2836
rect 50212 2796 50218 2808
rect 53558 2796 53564 2848
rect 53616 2836 53622 2848
rect 54205 2839 54263 2845
rect 54205 2836 54217 2839
rect 53616 2808 54217 2836
rect 53616 2796 53622 2808
rect 54205 2805 54217 2808
rect 54251 2805 54263 2839
rect 54205 2799 54263 2805
rect 55858 2796 55864 2848
rect 55916 2836 55922 2848
rect 57348 2836 57376 2935
rect 57606 2932 57612 2984
rect 57664 2972 57670 2984
rect 57977 2975 58035 2981
rect 57977 2972 57989 2975
rect 57664 2944 57989 2972
rect 57664 2932 57670 2944
rect 57977 2941 57989 2944
rect 58023 2941 58035 2975
rect 57977 2935 58035 2941
rect 59173 2975 59231 2981
rect 59173 2941 59185 2975
rect 59219 2972 59231 2975
rect 59219 2944 59492 2972
rect 59219 2941 59231 2944
rect 59173 2935 59231 2941
rect 58986 2864 58992 2916
rect 59044 2904 59050 2916
rect 59464 2913 59492 2944
rect 59538 2932 59544 2984
rect 59596 2972 59602 2984
rect 60001 2975 60059 2981
rect 60001 2972 60013 2975
rect 59596 2944 60013 2972
rect 59596 2932 59602 2944
rect 60001 2941 60013 2944
rect 60047 2941 60059 2975
rect 60001 2935 60059 2941
rect 60090 2932 60096 2984
rect 60148 2972 60154 2984
rect 60645 2975 60703 2981
rect 60645 2972 60657 2975
rect 60148 2944 60657 2972
rect 60148 2932 60154 2944
rect 60645 2941 60657 2944
rect 60691 2941 60703 2975
rect 60645 2935 60703 2941
rect 61381 2975 61439 2981
rect 61381 2941 61393 2975
rect 61427 2972 61439 2975
rect 61654 2972 61660 2984
rect 61427 2944 61660 2972
rect 61427 2941 61439 2944
rect 61381 2935 61439 2941
rect 61654 2932 61660 2944
rect 61712 2932 61718 2984
rect 62482 2932 62488 2984
rect 62540 2972 62546 2984
rect 62853 2975 62911 2981
rect 62853 2972 62865 2975
rect 62540 2944 62865 2972
rect 62540 2932 62546 2944
rect 62853 2941 62865 2944
rect 62899 2941 62911 2975
rect 62853 2935 62911 2941
rect 63405 2975 63463 2981
rect 63405 2941 63417 2975
rect 63451 2941 63463 2975
rect 63405 2935 63463 2941
rect 64417 2975 64475 2981
rect 64417 2941 64429 2975
rect 64463 2972 64475 2975
rect 64690 2972 64696 2984
rect 64463 2944 64696 2972
rect 64463 2941 64475 2944
rect 64417 2935 64475 2941
rect 59265 2907 59323 2913
rect 59265 2904 59277 2907
rect 59044 2876 59277 2904
rect 59044 2864 59050 2876
rect 59265 2873 59277 2876
rect 59311 2873 59323 2907
rect 59265 2867 59323 2873
rect 59449 2907 59507 2913
rect 59449 2873 59461 2907
rect 59495 2904 59507 2907
rect 59630 2904 59636 2916
rect 59495 2876 59636 2904
rect 59495 2873 59507 2876
rect 59449 2867 59507 2873
rect 59630 2864 59636 2876
rect 59688 2864 59694 2916
rect 61470 2904 61476 2916
rect 61431 2876 61476 2904
rect 61470 2864 61476 2876
rect 61528 2864 61534 2916
rect 62666 2904 62672 2916
rect 62627 2876 62672 2904
rect 62666 2864 62672 2876
rect 62724 2864 62730 2916
rect 55916 2808 57376 2836
rect 55916 2796 55922 2808
rect 60182 2796 60188 2848
rect 60240 2836 60246 2848
rect 62114 2836 62120 2848
rect 60240 2808 62120 2836
rect 60240 2796 60246 2808
rect 62114 2796 62120 2808
rect 62172 2796 62178 2848
rect 62482 2796 62488 2848
rect 62540 2836 62546 2848
rect 63420 2836 63448 2935
rect 64690 2932 64696 2944
rect 64748 2932 64754 2984
rect 64874 2932 64880 2984
rect 64932 2972 64938 2984
rect 65245 2975 65303 2981
rect 65245 2972 65257 2975
rect 64932 2944 65257 2972
rect 64932 2932 64938 2944
rect 65245 2941 65257 2944
rect 65291 2941 65303 2975
rect 65245 2935 65303 2941
rect 65518 2932 65524 2984
rect 65576 2972 65582 2984
rect 65889 2975 65947 2981
rect 65889 2972 65901 2975
rect 65576 2944 65901 2972
rect 65576 2932 65582 2944
rect 65889 2941 65901 2944
rect 65935 2941 65947 2975
rect 65889 2935 65947 2941
rect 66714 2932 66720 2984
rect 66772 2972 66778 2984
rect 67652 2981 67680 3012
rect 70397 3009 70409 3012
rect 70443 3040 70455 3043
rect 70443 3012 70808 3040
rect 70443 3009 70455 3012
rect 70397 3003 70455 3009
rect 67085 2975 67143 2981
rect 67085 2972 67097 2975
rect 66772 2944 67097 2972
rect 66772 2932 66778 2944
rect 67085 2941 67097 2944
rect 67131 2941 67143 2975
rect 67085 2935 67143 2941
rect 67637 2975 67695 2981
rect 67637 2941 67649 2975
rect 67683 2941 67695 2975
rect 67637 2935 67695 2941
rect 68281 2975 68339 2981
rect 68281 2941 68293 2975
rect 68327 2941 68339 2975
rect 68281 2935 68339 2941
rect 69661 2975 69719 2981
rect 69661 2941 69673 2975
rect 69707 2972 69719 2975
rect 69934 2972 69940 2984
rect 69707 2944 69940 2972
rect 69707 2941 69719 2944
rect 69661 2935 69719 2941
rect 64506 2904 64512 2916
rect 64467 2876 64512 2904
rect 64506 2864 64512 2876
rect 64564 2864 64570 2916
rect 66898 2904 66904 2916
rect 66859 2876 66904 2904
rect 66898 2864 66904 2876
rect 66956 2864 66962 2916
rect 67358 2864 67364 2916
rect 67416 2904 67422 2916
rect 68296 2904 68324 2935
rect 69934 2932 69940 2944
rect 69992 2932 69998 2984
rect 70780 2981 70808 3012
rect 70765 2975 70823 2981
rect 70765 2941 70777 2975
rect 70811 2941 70823 2975
rect 70765 2935 70823 2941
rect 71038 2932 71044 2984
rect 71096 2972 71102 2984
rect 71317 2975 71375 2981
rect 71317 2972 71329 2975
rect 71096 2944 71329 2972
rect 71096 2932 71102 2944
rect 71317 2941 71329 2944
rect 71363 2941 71375 2975
rect 71317 2935 71375 2941
rect 72234 2932 72240 2984
rect 72292 2972 72298 2984
rect 72605 2975 72663 2981
rect 72605 2972 72617 2975
rect 72292 2944 72617 2972
rect 72292 2932 72298 2944
rect 72605 2941 72617 2944
rect 72651 2941 72663 2975
rect 72605 2935 72663 2941
rect 73157 2975 73215 2981
rect 73157 2941 73169 2975
rect 73203 2941 73215 2975
rect 73157 2935 73215 2941
rect 67416 2876 68324 2904
rect 67416 2864 67422 2876
rect 69382 2864 69388 2916
rect 69440 2904 69446 2916
rect 69753 2907 69811 2913
rect 69753 2904 69765 2907
rect 69440 2876 69765 2904
rect 69440 2864 69446 2876
rect 69753 2873 69765 2876
rect 69799 2873 69811 2907
rect 70578 2904 70584 2916
rect 70539 2876 70584 2904
rect 69753 2867 69811 2873
rect 70578 2864 70584 2876
rect 70636 2864 70642 2916
rect 72418 2904 72424 2916
rect 72379 2876 72424 2904
rect 72418 2864 72424 2876
rect 72476 2864 72482 2916
rect 62540 2808 63448 2836
rect 62540 2796 62546 2808
rect 72234 2796 72240 2848
rect 72292 2836 72298 2848
rect 73172 2836 73200 2935
rect 73430 2932 73436 2984
rect 73488 2972 73494 2984
rect 73801 2975 73859 2981
rect 73801 2972 73813 2975
rect 73488 2944 73813 2972
rect 73488 2932 73494 2944
rect 73801 2941 73813 2944
rect 73847 2941 73859 2975
rect 73801 2935 73859 2941
rect 74813 2975 74871 2981
rect 74813 2941 74825 2975
rect 74859 2972 74871 2975
rect 75178 2972 75184 2984
rect 74859 2944 75184 2972
rect 74859 2941 74871 2944
rect 74813 2935 74871 2941
rect 75178 2932 75184 2944
rect 75236 2932 75242 2984
rect 75270 2932 75276 2984
rect 75328 2972 75334 2984
rect 75733 2975 75791 2981
rect 75733 2972 75745 2975
rect 75328 2944 75745 2972
rect 75328 2932 75334 2944
rect 75733 2941 75745 2944
rect 75779 2941 75791 2975
rect 75733 2935 75791 2941
rect 76561 2975 76619 2981
rect 76561 2941 76573 2975
rect 76607 2972 76619 2975
rect 76834 2972 76840 2984
rect 76607 2944 76840 2972
rect 76607 2941 76619 2944
rect 76561 2935 76619 2941
rect 76834 2932 76840 2944
rect 76892 2932 76898 2984
rect 77849 2975 77907 2981
rect 77849 2941 77861 2975
rect 77895 2972 77907 2975
rect 78125 2975 78183 2981
rect 78125 2972 78137 2975
rect 77895 2944 78137 2972
rect 77895 2941 77907 2944
rect 77849 2935 77907 2941
rect 78125 2941 78137 2944
rect 78171 2972 78183 2975
rect 78214 2972 78220 2984
rect 78171 2944 78220 2972
rect 78171 2941 78183 2944
rect 78125 2935 78183 2941
rect 78214 2932 78220 2944
rect 78272 2932 78278 2984
rect 79152 2981 79180 3080
rect 85114 3068 85120 3080
rect 85172 3068 85178 3120
rect 79962 3000 79968 3052
rect 80020 3040 80026 3052
rect 80020 3012 81848 3040
rect 80020 3000 80026 3012
rect 79137 2975 79195 2981
rect 79137 2941 79149 2975
rect 79183 2941 79195 2975
rect 80885 2975 80943 2981
rect 79137 2935 79195 2941
rect 79704 2944 80560 2972
rect 74902 2864 74908 2916
rect 74960 2904 74966 2916
rect 74997 2907 75055 2913
rect 74997 2904 75009 2907
rect 74960 2876 75009 2904
rect 74960 2864 74966 2876
rect 74997 2873 75009 2876
rect 75043 2873 75055 2907
rect 76650 2904 76656 2916
rect 76611 2876 76656 2904
rect 74997 2867 75055 2873
rect 76650 2864 76656 2876
rect 76708 2864 76714 2916
rect 77938 2904 77944 2916
rect 77899 2876 77944 2904
rect 77938 2864 77944 2876
rect 77996 2864 78002 2916
rect 78030 2864 78036 2916
rect 78088 2904 78094 2916
rect 79704 2904 79732 2944
rect 78088 2876 79732 2904
rect 78088 2864 78094 2876
rect 79778 2864 79784 2916
rect 79836 2904 79842 2916
rect 80241 2907 80299 2913
rect 80241 2904 80253 2907
rect 79836 2876 80253 2904
rect 79836 2864 79842 2876
rect 80241 2873 80253 2876
rect 80287 2873 80299 2907
rect 80422 2904 80428 2916
rect 80383 2876 80428 2904
rect 80241 2867 80299 2873
rect 80422 2864 80428 2876
rect 80480 2864 80486 2916
rect 80532 2904 80560 2944
rect 80885 2941 80897 2975
rect 80931 2972 80943 2975
rect 81161 2975 81219 2981
rect 81161 2972 81173 2975
rect 80931 2944 81173 2972
rect 80931 2941 80943 2944
rect 80885 2935 80943 2941
rect 81161 2941 81173 2944
rect 81207 2972 81219 2975
rect 81342 2972 81348 2984
rect 81207 2944 81348 2972
rect 81207 2941 81219 2944
rect 81161 2935 81219 2941
rect 81342 2932 81348 2944
rect 81400 2932 81406 2984
rect 81820 2981 81848 3012
rect 82354 3000 82360 3052
rect 82412 3040 82418 3052
rect 82906 3040 82912 3052
rect 82412 3012 82912 3040
rect 82412 3000 82418 3012
rect 82906 3000 82912 3012
rect 82964 3000 82970 3052
rect 91296 3040 91324 3136
rect 94501 3043 94559 3049
rect 94501 3040 94513 3043
rect 91296 3012 91692 3040
rect 81805 2975 81863 2981
rect 81805 2941 81817 2975
rect 81851 2941 81863 2975
rect 81805 2935 81863 2941
rect 82630 2932 82636 2984
rect 82688 2972 82694 2984
rect 83185 2975 83243 2981
rect 83185 2972 83197 2975
rect 82688 2944 83197 2972
rect 82688 2932 82694 2944
rect 83185 2941 83197 2944
rect 83231 2941 83243 2975
rect 83185 2935 83243 2941
rect 83274 2932 83280 2984
rect 83332 2972 83338 2984
rect 83829 2975 83887 2981
rect 83829 2972 83841 2975
rect 83332 2944 83841 2972
rect 83332 2932 83338 2944
rect 83829 2941 83841 2944
rect 83875 2941 83887 2975
rect 83829 2935 83887 2941
rect 83918 2932 83924 2984
rect 83976 2972 83982 2984
rect 85485 2975 85543 2981
rect 85485 2972 85497 2975
rect 83976 2944 85497 2972
rect 83976 2932 83982 2944
rect 85485 2941 85497 2944
rect 85531 2941 85543 2975
rect 85485 2935 85543 2941
rect 86129 2975 86187 2981
rect 86129 2941 86141 2975
rect 86175 2941 86187 2975
rect 86129 2935 86187 2941
rect 82541 2907 82599 2913
rect 82541 2904 82553 2907
rect 80532 2876 82553 2904
rect 82541 2873 82553 2876
rect 82587 2873 82599 2907
rect 82541 2867 82599 2873
rect 84378 2864 84384 2916
rect 84436 2904 84442 2916
rect 86144 2904 86172 2935
rect 86218 2932 86224 2984
rect 86276 2972 86282 2984
rect 86773 2975 86831 2981
rect 86773 2972 86785 2975
rect 86276 2944 86785 2972
rect 86276 2932 86282 2944
rect 86773 2941 86785 2944
rect 86819 2941 86831 2975
rect 86773 2935 86831 2941
rect 86862 2932 86868 2984
rect 86920 2972 86926 2984
rect 87417 2975 87475 2981
rect 87417 2972 87429 2975
rect 86920 2944 87429 2972
rect 86920 2932 86926 2944
rect 87417 2941 87429 2944
rect 87463 2941 87475 2975
rect 87417 2935 87475 2941
rect 87506 2932 87512 2984
rect 87564 2972 87570 2984
rect 88061 2975 88119 2981
rect 88061 2972 88073 2975
rect 87564 2944 88073 2972
rect 87564 2932 87570 2944
rect 88061 2941 88073 2944
rect 88107 2941 88119 2975
rect 88061 2935 88119 2941
rect 88150 2932 88156 2984
rect 88208 2972 88214 2984
rect 88705 2975 88763 2981
rect 88705 2972 88717 2975
rect 88208 2944 88717 2972
rect 88208 2932 88214 2944
rect 88705 2941 88717 2944
rect 88751 2941 88763 2975
rect 88705 2935 88763 2941
rect 88794 2932 88800 2984
rect 88852 2972 88858 2984
rect 89349 2975 89407 2981
rect 89349 2972 89361 2975
rect 88852 2944 89361 2972
rect 88852 2932 88858 2944
rect 89349 2941 89361 2944
rect 89395 2941 89407 2975
rect 89349 2935 89407 2941
rect 90818 2932 90824 2984
rect 90876 2972 90882 2984
rect 90913 2975 90971 2981
rect 90913 2972 90925 2975
rect 90876 2944 90925 2972
rect 90876 2932 90882 2944
rect 90913 2941 90925 2944
rect 90959 2941 90971 2975
rect 90913 2935 90971 2941
rect 91278 2932 91284 2984
rect 91336 2972 91342 2984
rect 91664 2981 91692 3012
rect 92952 3012 94513 3040
rect 91465 2975 91523 2981
rect 91465 2972 91477 2975
rect 91336 2944 91477 2972
rect 91336 2932 91342 2944
rect 91465 2941 91477 2944
rect 91511 2941 91523 2975
rect 91465 2935 91523 2941
rect 91649 2975 91707 2981
rect 91649 2941 91661 2975
rect 91695 2941 91707 2975
rect 91649 2935 91707 2941
rect 91738 2932 91744 2984
rect 91796 2972 91802 2984
rect 92201 2975 92259 2981
rect 92201 2972 92213 2975
rect 91796 2944 92213 2972
rect 91796 2932 91802 2944
rect 92201 2941 92213 2944
rect 92247 2941 92259 2975
rect 92201 2935 92259 2941
rect 84436 2876 86172 2904
rect 84436 2864 84442 2876
rect 90082 2864 90088 2916
rect 90140 2904 90146 2916
rect 90729 2907 90787 2913
rect 90729 2904 90741 2907
rect 90140 2876 90741 2904
rect 90140 2864 90146 2876
rect 90729 2873 90741 2876
rect 90775 2873 90787 2907
rect 90729 2867 90787 2873
rect 91002 2864 91008 2916
rect 91060 2904 91066 2916
rect 92952 2904 92980 3012
rect 94501 3009 94513 3012
rect 94547 3040 94559 3043
rect 94547 3012 94820 3040
rect 94547 3009 94559 3012
rect 94501 3003 94559 3009
rect 93670 2932 93676 2984
rect 93728 2972 93734 2984
rect 94041 2975 94099 2981
rect 94041 2972 94053 2975
rect 93728 2944 94053 2972
rect 93728 2932 93734 2944
rect 94041 2941 94053 2944
rect 94087 2941 94099 2975
rect 94041 2935 94099 2941
rect 94406 2932 94412 2984
rect 94464 2972 94470 2984
rect 94792 2981 94820 3012
rect 94593 2975 94651 2981
rect 94593 2972 94605 2975
rect 94464 2944 94605 2972
rect 94464 2932 94470 2944
rect 94593 2941 94605 2944
rect 94639 2941 94651 2975
rect 94593 2935 94651 2941
rect 94777 2975 94835 2981
rect 94777 2941 94789 2975
rect 94823 2941 94835 2975
rect 96062 2972 96068 2984
rect 96023 2944 96068 2972
rect 94777 2935 94835 2941
rect 96062 2932 96068 2944
rect 96120 2932 96126 2984
rect 96798 2932 96804 2984
rect 96856 2972 96862 2984
rect 97721 2975 97779 2981
rect 97721 2972 97733 2975
rect 96856 2944 97733 2972
rect 96856 2932 96862 2944
rect 97721 2941 97733 2944
rect 97767 2941 97779 2975
rect 97721 2935 97779 2941
rect 93118 2904 93124 2916
rect 91060 2876 92980 2904
rect 93079 2876 93124 2904
rect 91060 2864 91066 2876
rect 93118 2864 93124 2876
rect 93176 2864 93182 2916
rect 93305 2907 93363 2913
rect 93305 2873 93317 2907
rect 93351 2873 93363 2907
rect 93305 2867 93363 2873
rect 72292 2808 73200 2836
rect 72292 2796 72298 2808
rect 73614 2796 73620 2848
rect 73672 2836 73678 2848
rect 74718 2836 74724 2848
rect 73672 2808 74724 2836
rect 73672 2796 73678 2808
rect 74718 2796 74724 2808
rect 74776 2796 74782 2848
rect 76098 2796 76104 2848
rect 76156 2836 76162 2848
rect 77294 2836 77300 2848
rect 76156 2808 77300 2836
rect 76156 2796 76162 2808
rect 77294 2796 77300 2808
rect 77352 2796 77358 2848
rect 79226 2836 79232 2848
rect 79187 2808 79232 2836
rect 79226 2796 79232 2808
rect 79284 2796 79290 2848
rect 80330 2796 80336 2848
rect 80388 2836 80394 2848
rect 81069 2839 81127 2845
rect 81069 2836 81081 2839
rect 80388 2808 81081 2836
rect 80388 2796 80394 2808
rect 81069 2805 81081 2808
rect 81115 2805 81127 2839
rect 81069 2799 81127 2805
rect 82170 2796 82176 2848
rect 82228 2836 82234 2848
rect 82633 2839 82691 2845
rect 82633 2836 82645 2839
rect 82228 2808 82645 2836
rect 82228 2796 82234 2808
rect 82633 2805 82645 2808
rect 82679 2805 82691 2839
rect 82633 2799 82691 2805
rect 87046 2796 87052 2848
rect 87104 2836 87110 2848
rect 89622 2836 89628 2848
rect 87104 2808 89628 2836
rect 87104 2796 87110 2808
rect 89622 2796 89628 2808
rect 89680 2796 89686 2848
rect 90358 2796 90364 2848
rect 90416 2836 90422 2848
rect 92937 2839 92995 2845
rect 92937 2836 92949 2839
rect 90416 2808 92949 2836
rect 90416 2796 90422 2808
rect 92937 2805 92949 2808
rect 92983 2836 92995 2839
rect 93320 2836 93348 2867
rect 93762 2864 93768 2916
rect 93820 2904 93826 2916
rect 93857 2907 93915 2913
rect 93857 2904 93869 2907
rect 93820 2876 93869 2904
rect 93820 2864 93826 2876
rect 93857 2873 93869 2876
rect 93903 2873 93915 2907
rect 93857 2867 93915 2873
rect 96246 2864 96252 2916
rect 96304 2904 96310 2916
rect 96709 2907 96767 2913
rect 96709 2904 96721 2907
rect 96304 2876 96721 2904
rect 96304 2864 96310 2876
rect 96709 2873 96721 2876
rect 96755 2873 96767 2907
rect 96709 2867 96767 2873
rect 96893 2907 96951 2913
rect 96893 2873 96905 2907
rect 96939 2904 96951 2907
rect 97261 2907 97319 2913
rect 97261 2904 97273 2907
rect 96939 2876 97273 2904
rect 96939 2873 96951 2876
rect 96893 2867 96951 2873
rect 97261 2873 97273 2876
rect 97307 2873 97319 2907
rect 97534 2904 97540 2916
rect 97495 2876 97540 2904
rect 97261 2867 97319 2873
rect 97534 2864 97540 2876
rect 97592 2864 97598 2916
rect 92983 2808 93348 2836
rect 92983 2805 92995 2808
rect 92937 2799 92995 2805
rect 95602 2796 95608 2848
rect 95660 2836 95666 2848
rect 96157 2839 96215 2845
rect 96157 2836 96169 2839
rect 95660 2808 96169 2836
rect 95660 2796 95666 2808
rect 96157 2805 96169 2808
rect 96203 2805 96215 2839
rect 96157 2799 96215 2805
rect 97718 2796 97724 2848
rect 97776 2836 97782 2848
rect 99834 2836 99840 2848
rect 97776 2808 99840 2836
rect 97776 2796 97782 2808
rect 99834 2796 99840 2808
rect 99892 2796 99898 2848
rect 1104 2746 98808 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 50326 2746
rect 50378 2694 50390 2746
rect 50442 2694 50454 2746
rect 50506 2694 50518 2746
rect 50570 2694 81046 2746
rect 81098 2694 81110 2746
rect 81162 2694 81174 2746
rect 81226 2694 81238 2746
rect 81290 2694 98808 2746
rect 1104 2672 98808 2694
rect 8478 2632 8484 2644
rect 8439 2604 8484 2632
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 13449 2635 13507 2641
rect 13449 2601 13461 2635
rect 13495 2632 13507 2635
rect 22738 2632 22744 2644
rect 13495 2604 13860 2632
rect 22699 2604 22744 2632
rect 13495 2601 13507 2604
rect 13449 2595 13507 2601
rect 13832 2576 13860 2604
rect 22738 2592 22744 2604
rect 22796 2632 22802 2644
rect 22796 2604 23152 2632
rect 22796 2592 22802 2604
rect 2130 2524 2136 2576
rect 2188 2564 2194 2576
rect 2225 2567 2283 2573
rect 2225 2564 2237 2567
rect 2188 2536 2237 2564
rect 2188 2524 2194 2536
rect 2225 2533 2237 2536
rect 2271 2533 2283 2567
rect 2225 2527 2283 2533
rect 3145 2567 3203 2573
rect 3145 2533 3157 2567
rect 3191 2564 3203 2567
rect 3234 2564 3240 2576
rect 3191 2536 3240 2564
rect 3191 2533 3203 2536
rect 3145 2527 3203 2533
rect 3234 2524 3240 2536
rect 3292 2524 3298 2576
rect 4982 2564 4988 2576
rect 4943 2536 4988 2564
rect 4982 2524 4988 2536
rect 5040 2524 5046 2576
rect 7650 2564 7656 2576
rect 7611 2536 7656 2564
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 10410 2564 10416 2576
rect 10371 2536 10416 2564
rect 10410 2524 10416 2536
rect 10468 2524 10474 2576
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 11698 2564 11704 2576
rect 11195 2536 11704 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 12250 2564 12256 2576
rect 12211 2536 12256 2564
rect 12250 2524 12256 2536
rect 12308 2524 12314 2576
rect 13081 2567 13139 2573
rect 13081 2533 13093 2567
rect 13127 2564 13139 2567
rect 13538 2564 13544 2576
rect 13127 2536 13544 2564
rect 13127 2533 13139 2536
rect 13081 2527 13139 2533
rect 13538 2524 13544 2536
rect 13596 2524 13602 2576
rect 13814 2564 13820 2576
rect 13775 2536 13820 2564
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 15562 2564 15568 2576
rect 15523 2536 15568 2564
rect 15562 2524 15568 2536
rect 15620 2524 15626 2576
rect 16666 2564 16672 2576
rect 16627 2536 16672 2564
rect 16666 2524 16672 2536
rect 16724 2524 16730 2576
rect 18414 2564 18420 2576
rect 18375 2536 18420 2564
rect 18414 2524 18420 2536
rect 18472 2524 18478 2576
rect 18969 2567 19027 2573
rect 18969 2533 18981 2567
rect 19015 2564 19027 2567
rect 19150 2564 19156 2576
rect 19015 2536 19156 2564
rect 19015 2533 19027 2536
rect 18969 2527 19027 2533
rect 19150 2524 19156 2536
rect 19208 2564 19214 2576
rect 19245 2567 19303 2573
rect 19245 2564 19257 2567
rect 19208 2536 19257 2564
rect 19208 2524 19214 2536
rect 19245 2533 19257 2536
rect 19291 2533 19303 2567
rect 19245 2527 19303 2533
rect 20349 2567 20407 2573
rect 20349 2533 20361 2567
rect 20395 2564 20407 2567
rect 20530 2564 20536 2576
rect 20395 2536 20536 2564
rect 20395 2533 20407 2536
rect 20349 2527 20407 2533
rect 20530 2524 20536 2536
rect 20588 2524 20594 2576
rect 21818 2564 21824 2576
rect 21779 2536 21824 2564
rect 21818 2524 21824 2536
rect 21876 2524 21882 2576
rect 23124 2573 23152 2604
rect 26786 2592 26792 2644
rect 26844 2632 26850 2644
rect 26881 2635 26939 2641
rect 26881 2632 26893 2635
rect 26844 2604 26893 2632
rect 26844 2592 26850 2604
rect 26881 2601 26893 2604
rect 26927 2632 26939 2635
rect 28169 2635 28227 2641
rect 26927 2604 27292 2632
rect 26927 2601 26939 2604
rect 26881 2595 26939 2601
rect 23109 2567 23167 2573
rect 23109 2533 23121 2567
rect 23155 2533 23167 2567
rect 23109 2527 23167 2533
rect 23569 2567 23627 2573
rect 23569 2533 23581 2567
rect 23615 2564 23627 2567
rect 23842 2564 23848 2576
rect 23615 2536 23848 2564
rect 23615 2533 23627 2536
rect 23569 2527 23627 2533
rect 23842 2524 23848 2536
rect 23900 2524 23906 2576
rect 24486 2564 24492 2576
rect 24447 2536 24492 2564
rect 24486 2524 24492 2536
rect 24544 2524 24550 2576
rect 25501 2567 25559 2573
rect 25501 2533 25513 2567
rect 25547 2564 25559 2567
rect 25774 2564 25780 2576
rect 25547 2536 25780 2564
rect 25547 2533 25559 2536
rect 25501 2527 25559 2533
rect 25774 2524 25780 2536
rect 25832 2524 25838 2576
rect 27264 2573 27292 2604
rect 28169 2601 28181 2635
rect 28215 2632 28227 2635
rect 28626 2632 28632 2644
rect 28215 2604 28632 2632
rect 28215 2601 28227 2604
rect 28169 2595 28227 2601
rect 28460 2573 28488 2604
rect 28626 2592 28632 2604
rect 28684 2592 28690 2644
rect 28810 2632 28816 2644
rect 28771 2604 28816 2632
rect 28810 2592 28816 2604
rect 28868 2632 28874 2644
rect 29638 2632 29644 2644
rect 28868 2604 29224 2632
rect 29599 2604 29644 2632
rect 28868 2592 28874 2604
rect 29196 2573 29224 2604
rect 29638 2592 29644 2604
rect 29696 2632 29702 2644
rect 29696 2604 29960 2632
rect 29696 2592 29702 2604
rect 29932 2573 29960 2604
rect 30374 2592 30380 2644
rect 30432 2632 30438 2644
rect 30745 2635 30803 2641
rect 30745 2632 30757 2635
rect 30432 2604 30757 2632
rect 30432 2592 30438 2604
rect 30745 2601 30757 2604
rect 30791 2632 30803 2635
rect 31478 2632 31484 2644
rect 30791 2604 31156 2632
rect 31439 2604 31484 2632
rect 30791 2601 30803 2604
rect 30745 2595 30803 2601
rect 31128 2573 31156 2604
rect 31478 2592 31484 2604
rect 31536 2632 31542 2644
rect 32033 2635 32091 2641
rect 32033 2632 32045 2635
rect 31536 2604 32045 2632
rect 31536 2592 31542 2604
rect 31864 2573 31892 2604
rect 32033 2601 32045 2604
rect 32079 2601 32091 2635
rect 34146 2632 34152 2644
rect 34107 2604 34152 2632
rect 32033 2595 32091 2601
rect 34146 2592 34152 2604
rect 34204 2632 34210 2644
rect 35986 2632 35992 2644
rect 34204 2604 34560 2632
rect 34204 2592 34210 2604
rect 27249 2567 27307 2573
rect 27249 2533 27261 2567
rect 27295 2533 27307 2567
rect 27249 2527 27307 2533
rect 28445 2567 28503 2573
rect 28445 2533 28457 2567
rect 28491 2533 28503 2567
rect 28445 2527 28503 2533
rect 29181 2567 29239 2573
rect 29181 2533 29193 2567
rect 29227 2533 29239 2567
rect 29181 2527 29239 2533
rect 29917 2567 29975 2573
rect 29917 2533 29929 2567
rect 29963 2533 29975 2567
rect 29917 2527 29975 2533
rect 31113 2567 31171 2573
rect 31113 2533 31125 2567
rect 31159 2533 31171 2567
rect 31113 2527 31171 2533
rect 31849 2567 31907 2573
rect 31849 2533 31861 2567
rect 31895 2533 31907 2567
rect 31849 2527 31907 2533
rect 32309 2567 32367 2573
rect 32309 2533 32321 2567
rect 32355 2564 32367 2567
rect 32585 2567 32643 2573
rect 32585 2564 32597 2567
rect 32355 2536 32597 2564
rect 32355 2533 32367 2536
rect 32309 2527 32367 2533
rect 32585 2533 32597 2536
rect 32631 2564 32643 2567
rect 32674 2564 32680 2576
rect 32631 2536 32680 2564
rect 32631 2533 32643 2536
rect 32585 2527 32643 2533
rect 32674 2524 32680 2536
rect 32732 2524 32738 2576
rect 33686 2564 33692 2576
rect 33647 2536 33692 2564
rect 33686 2524 33692 2536
rect 33744 2524 33750 2576
rect 34532 2573 34560 2604
rect 35866 2604 35992 2632
rect 34517 2567 34575 2573
rect 34517 2533 34529 2567
rect 34563 2533 34575 2567
rect 34517 2527 34575 2533
rect 35161 2567 35219 2573
rect 35161 2533 35173 2567
rect 35207 2564 35219 2567
rect 35866 2564 35894 2604
rect 35986 2592 35992 2604
rect 36044 2592 36050 2644
rect 36170 2632 36176 2644
rect 36131 2604 36176 2632
rect 36170 2592 36176 2604
rect 36228 2632 36234 2644
rect 36633 2635 36691 2641
rect 36633 2632 36645 2635
rect 36228 2604 36645 2632
rect 36228 2592 36234 2604
rect 36464 2573 36492 2604
rect 36633 2601 36645 2604
rect 36679 2601 36691 2635
rect 36906 2632 36912 2644
rect 36867 2604 36912 2632
rect 36633 2595 36691 2601
rect 36906 2592 36912 2604
rect 36964 2632 36970 2644
rect 38841 2635 38899 2641
rect 36964 2604 37228 2632
rect 36964 2592 36970 2604
rect 37200 2573 37228 2604
rect 38841 2601 38853 2635
rect 38887 2632 38899 2635
rect 39390 2632 39396 2644
rect 38887 2604 39396 2632
rect 38887 2601 38899 2604
rect 38841 2595 38899 2601
rect 35207 2536 35894 2564
rect 36449 2567 36507 2573
rect 35207 2533 35219 2536
rect 35161 2527 35219 2533
rect 36449 2533 36461 2567
rect 36495 2533 36507 2567
rect 36449 2527 36507 2533
rect 37185 2567 37243 2573
rect 37185 2533 37197 2567
rect 37231 2533 37243 2567
rect 37185 2527 37243 2533
rect 37645 2567 37703 2573
rect 37645 2533 37657 2567
rect 37691 2564 37703 2567
rect 37918 2564 37924 2576
rect 37691 2536 37924 2564
rect 37691 2533 37703 2536
rect 37645 2527 37703 2533
rect 37918 2524 37924 2536
rect 37976 2524 37982 2576
rect 38930 2564 38936 2576
rect 38891 2536 38936 2564
rect 38930 2524 38936 2536
rect 38988 2524 38994 2576
rect 39132 2573 39160 2604
rect 39390 2592 39396 2604
rect 39448 2592 39454 2644
rect 40034 2592 40040 2644
rect 40092 2632 40098 2644
rect 40221 2635 40279 2641
rect 40221 2632 40233 2635
rect 40092 2604 40233 2632
rect 40092 2592 40098 2604
rect 40221 2601 40233 2604
rect 40267 2632 40279 2635
rect 41414 2632 41420 2644
rect 40267 2604 40632 2632
rect 41375 2604 41420 2632
rect 40267 2601 40279 2604
rect 40221 2595 40279 2601
rect 39117 2567 39175 2573
rect 39117 2533 39129 2567
rect 39163 2533 39175 2567
rect 39117 2527 39175 2533
rect 39577 2567 39635 2573
rect 39577 2533 39589 2567
rect 39623 2564 39635 2567
rect 39850 2564 39856 2576
rect 39623 2536 39856 2564
rect 39623 2533 39635 2536
rect 39577 2527 39635 2533
rect 39850 2524 39856 2536
rect 39908 2524 39914 2576
rect 40604 2573 40632 2604
rect 41414 2592 41420 2604
rect 41472 2592 41478 2644
rect 45002 2592 45008 2644
rect 45060 2632 45066 2644
rect 48593 2635 48651 2641
rect 48593 2632 48605 2635
rect 45060 2604 48605 2632
rect 45060 2592 45066 2604
rect 48593 2601 48605 2604
rect 48639 2601 48651 2635
rect 49418 2632 49424 2644
rect 49379 2604 49424 2632
rect 48593 2595 48651 2601
rect 49418 2592 49424 2604
rect 49476 2632 49482 2644
rect 49476 2604 49832 2632
rect 49476 2592 49482 2604
rect 40589 2567 40647 2573
rect 40589 2533 40601 2567
rect 40635 2533 40647 2567
rect 40589 2527 40647 2533
rect 290 2456 296 2508
rect 348 2496 354 2508
rect 1397 2499 1455 2505
rect 1397 2496 1409 2499
rect 348 2468 1409 2496
rect 348 2456 354 2468
rect 1397 2465 1409 2468
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 2884 2428 2912 2459
rect 3878 2456 3884 2508
rect 3936 2496 3942 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 3936 2468 4261 2496
rect 3936 2456 3942 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 5626 2496 5632 2508
rect 5587 2468 5632 2496
rect 4249 2459 4307 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 6546 2456 6552 2508
rect 6604 2496 6610 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6604 2468 6929 2496
rect 6604 2456 6610 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 8297 2499 8355 2505
rect 8297 2496 8309 2499
rect 6917 2459 6975 2465
rect 7576 2468 8309 2496
rect 1360 2400 2912 2428
rect 1360 2388 1366 2400
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 7576 2428 7604 2468
rect 8297 2465 8309 2468
rect 8343 2465 8355 2499
rect 8297 2459 8355 2465
rect 9582 2456 9588 2508
rect 9640 2496 9646 2508
rect 9677 2499 9735 2505
rect 9677 2496 9689 2499
rect 9640 2468 9689 2496
rect 9640 2456 9646 2468
rect 9677 2465 9689 2468
rect 9723 2465 9735 2499
rect 9677 2459 9735 2465
rect 13262 2456 13268 2508
rect 13320 2496 13326 2508
rect 15013 2499 15071 2505
rect 15013 2496 15025 2499
rect 13320 2468 15025 2496
rect 13320 2456 13326 2468
rect 15013 2465 15025 2468
rect 15059 2465 15071 2499
rect 15013 2459 15071 2465
rect 16301 2499 16359 2505
rect 16301 2465 16313 2499
rect 16347 2496 16359 2499
rect 16942 2496 16948 2508
rect 16347 2468 16948 2496
rect 16347 2465 16359 2468
rect 16301 2459 16359 2465
rect 16942 2456 16948 2468
rect 17000 2456 17006 2508
rect 17586 2496 17592 2508
rect 17547 2468 17592 2496
rect 17586 2456 17592 2468
rect 17644 2456 17650 2508
rect 21174 2496 21180 2508
rect 21135 2468 21180 2496
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 24210 2456 24216 2508
rect 24268 2496 24274 2508
rect 26237 2499 26295 2505
rect 24268 2468 25728 2496
rect 24268 2456 24274 2468
rect 5776 2400 7604 2428
rect 5776 2388 5782 2400
rect 14734 2388 14740 2440
rect 14792 2428 14798 2440
rect 19061 2431 19119 2437
rect 19061 2428 19073 2431
rect 14792 2400 19073 2428
rect 14792 2388 14798 2400
rect 19061 2397 19073 2400
rect 19107 2397 19119 2431
rect 19061 2391 19119 2397
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 23716 2400 25605 2428
rect 23716 2388 23722 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25700 2428 25728 2468
rect 26237 2465 26249 2499
rect 26283 2496 26295 2499
rect 26513 2499 26571 2505
rect 26513 2496 26525 2499
rect 26283 2468 26525 2496
rect 26283 2465 26295 2468
rect 26237 2459 26295 2465
rect 26513 2465 26525 2468
rect 26559 2496 26571 2499
rect 27430 2496 27436 2508
rect 26559 2468 27436 2496
rect 26559 2465 26571 2468
rect 26513 2459 26571 2465
rect 27430 2456 27436 2468
rect 27488 2456 27494 2508
rect 33410 2456 33416 2508
rect 33468 2496 33474 2508
rect 36265 2499 36323 2505
rect 36265 2496 36277 2499
rect 33468 2468 36277 2496
rect 33468 2456 33474 2468
rect 36265 2465 36277 2468
rect 36311 2465 36323 2499
rect 36265 2459 36323 2465
rect 38746 2456 38752 2508
rect 38804 2496 38810 2508
rect 40405 2499 40463 2505
rect 40405 2496 40417 2499
rect 38804 2468 40417 2496
rect 38804 2456 38810 2468
rect 40405 2465 40417 2468
rect 40451 2465 40463 2499
rect 41432 2496 41460 2592
rect 42426 2564 42432 2576
rect 42387 2536 42432 2564
rect 42426 2524 42432 2536
rect 42484 2524 42490 2576
rect 42981 2567 43039 2573
rect 42981 2533 42993 2567
rect 43027 2564 43039 2567
rect 43257 2567 43315 2573
rect 43257 2564 43269 2567
rect 43027 2536 43269 2564
rect 43027 2533 43039 2536
rect 42981 2527 43039 2533
rect 43257 2533 43269 2536
rect 43303 2564 43315 2567
rect 43806 2564 43812 2576
rect 43303 2536 43812 2564
rect 43303 2533 43315 2536
rect 43257 2527 43315 2533
rect 43806 2524 43812 2536
rect 43864 2524 43870 2576
rect 44177 2567 44235 2573
rect 44177 2533 44189 2567
rect 44223 2564 44235 2567
rect 44358 2564 44364 2576
rect 44223 2536 44364 2564
rect 44223 2533 44235 2536
rect 44177 2527 44235 2533
rect 44358 2524 44364 2536
rect 44416 2564 44422 2576
rect 44453 2567 44511 2573
rect 44453 2564 44465 2567
rect 44416 2536 44465 2564
rect 44416 2524 44422 2536
rect 44453 2533 44465 2536
rect 44499 2533 44511 2567
rect 45094 2564 45100 2576
rect 45055 2536 45100 2564
rect 44453 2527 44511 2533
rect 45094 2524 45100 2536
rect 45152 2524 45158 2576
rect 45649 2567 45707 2573
rect 45649 2533 45661 2567
rect 45695 2564 45707 2567
rect 45922 2564 45928 2576
rect 45695 2536 45928 2564
rect 45695 2533 45707 2536
rect 45649 2527 45707 2533
rect 45922 2524 45928 2536
rect 45980 2564 45986 2576
rect 46109 2567 46167 2573
rect 46109 2564 46121 2567
rect 45980 2536 46121 2564
rect 45980 2524 45986 2536
rect 46109 2533 46121 2536
rect 46155 2533 46167 2567
rect 46109 2527 46167 2533
rect 47029 2567 47087 2573
rect 47029 2533 47041 2567
rect 47075 2564 47087 2567
rect 48130 2564 48136 2576
rect 47075 2536 48136 2564
rect 47075 2533 47087 2536
rect 47029 2527 47087 2533
rect 48130 2524 48136 2536
rect 48188 2524 48194 2576
rect 48498 2564 48504 2576
rect 48459 2536 48504 2564
rect 48498 2524 48504 2536
rect 48556 2524 48562 2576
rect 49804 2573 49832 2604
rect 50706 2592 50712 2644
rect 50764 2632 50770 2644
rect 50893 2635 50951 2641
rect 50893 2632 50905 2635
rect 50764 2604 50905 2632
rect 50764 2592 50770 2604
rect 50893 2601 50905 2604
rect 50939 2632 50951 2635
rect 54754 2632 54760 2644
rect 50939 2604 51304 2632
rect 54715 2604 54760 2632
rect 50939 2601 50951 2604
rect 50893 2595 50951 2601
rect 49789 2567 49847 2573
rect 49789 2533 49801 2567
rect 49835 2533 49847 2567
rect 49789 2527 49847 2533
rect 50249 2567 50307 2573
rect 50249 2533 50261 2567
rect 50295 2564 50307 2567
rect 50525 2567 50583 2573
rect 50525 2564 50537 2567
rect 50295 2536 50537 2564
rect 50295 2533 50307 2536
rect 50249 2527 50307 2533
rect 50525 2533 50537 2536
rect 50571 2564 50583 2567
rect 50982 2564 50988 2576
rect 50571 2536 50988 2564
rect 50571 2533 50583 2536
rect 50525 2527 50583 2533
rect 50982 2524 50988 2536
rect 51040 2524 51046 2576
rect 51276 2573 51304 2604
rect 54754 2592 54760 2604
rect 54812 2632 54818 2644
rect 54812 2604 55168 2632
rect 54812 2592 54818 2604
rect 51261 2567 51319 2573
rect 51261 2533 51273 2567
rect 51307 2533 51319 2567
rect 52362 2564 52368 2576
rect 52323 2536 52368 2564
rect 51261 2527 51319 2533
rect 52362 2524 52368 2536
rect 52420 2524 52426 2576
rect 52917 2567 52975 2573
rect 52917 2533 52929 2567
rect 52963 2564 52975 2567
rect 53193 2567 53251 2573
rect 53193 2564 53205 2567
rect 52963 2536 53205 2564
rect 52963 2533 52975 2536
rect 52917 2527 52975 2533
rect 53193 2533 53205 2536
rect 53239 2564 53251 2567
rect 53650 2564 53656 2576
rect 53239 2536 53656 2564
rect 53239 2533 53251 2536
rect 53193 2527 53251 2533
rect 53650 2524 53656 2536
rect 53708 2524 53714 2576
rect 53834 2564 53840 2576
rect 53795 2536 53840 2564
rect 53834 2524 53840 2536
rect 53892 2524 53898 2576
rect 55140 2573 55168 2604
rect 58066 2592 58072 2644
rect 58124 2632 58130 2644
rect 58161 2635 58219 2641
rect 58161 2632 58173 2635
rect 58124 2604 58173 2632
rect 58124 2592 58130 2604
rect 58161 2601 58173 2604
rect 58207 2632 58219 2635
rect 60185 2635 60243 2641
rect 58207 2604 58572 2632
rect 58207 2601 58219 2604
rect 58161 2595 58219 2601
rect 55125 2567 55183 2573
rect 55125 2533 55137 2567
rect 55171 2533 55183 2567
rect 55766 2564 55772 2576
rect 55727 2536 55772 2564
rect 55125 2527 55183 2533
rect 55766 2524 55772 2536
rect 55824 2524 55830 2576
rect 56321 2567 56379 2573
rect 56321 2533 56333 2567
rect 56367 2564 56379 2567
rect 56597 2567 56655 2573
rect 56597 2564 56609 2567
rect 56367 2536 56609 2564
rect 56367 2533 56379 2536
rect 56321 2527 56379 2533
rect 56597 2533 56609 2536
rect 56643 2564 56655 2567
rect 56686 2564 56692 2576
rect 56643 2536 56692 2564
rect 56643 2533 56655 2536
rect 56597 2527 56655 2533
rect 56686 2524 56692 2536
rect 56744 2524 56750 2576
rect 57517 2567 57575 2573
rect 57517 2533 57529 2567
rect 57563 2564 57575 2567
rect 57790 2564 57796 2576
rect 57563 2536 57796 2564
rect 57563 2533 57575 2536
rect 57517 2527 57575 2533
rect 57790 2524 57796 2536
rect 57848 2524 57854 2576
rect 58342 2564 58348 2576
rect 58303 2536 58348 2564
rect 58342 2524 58348 2536
rect 58400 2524 58406 2576
rect 58544 2573 58572 2604
rect 60185 2601 60197 2635
rect 60231 2632 60243 2635
rect 60274 2632 60280 2644
rect 60231 2604 60280 2632
rect 60231 2601 60243 2604
rect 60185 2595 60243 2601
rect 60274 2592 60280 2604
rect 60332 2632 60338 2644
rect 61657 2635 61715 2641
rect 60332 2604 60504 2632
rect 60332 2592 60338 2604
rect 58529 2567 58587 2573
rect 58529 2533 58541 2567
rect 58575 2533 58587 2567
rect 58529 2527 58587 2533
rect 58989 2567 59047 2573
rect 58989 2533 59001 2567
rect 59035 2564 59047 2567
rect 59262 2564 59268 2576
rect 59035 2536 59268 2564
rect 59035 2533 59047 2536
rect 58989 2527 59047 2533
rect 59262 2524 59268 2536
rect 59320 2524 59326 2576
rect 60476 2573 60504 2604
rect 61657 2601 61669 2635
rect 61703 2632 61715 2635
rect 61703 2604 61976 2632
rect 61703 2601 61715 2604
rect 61657 2595 61715 2601
rect 61948 2576 61976 2604
rect 62022 2592 62028 2644
rect 62080 2632 62086 2644
rect 65705 2635 65763 2641
rect 65705 2632 65717 2635
rect 62080 2604 65717 2632
rect 62080 2592 62086 2604
rect 65705 2601 65717 2604
rect 65751 2601 65763 2635
rect 66254 2632 66260 2644
rect 66215 2604 66260 2632
rect 65705 2595 65763 2601
rect 66254 2592 66260 2604
rect 66312 2632 66318 2644
rect 68830 2632 68836 2644
rect 66312 2604 66576 2632
rect 68791 2604 68836 2632
rect 66312 2592 66318 2604
rect 60461 2567 60519 2573
rect 60461 2533 60473 2567
rect 60507 2533 60519 2567
rect 60461 2527 60519 2533
rect 60921 2567 60979 2573
rect 60921 2533 60933 2567
rect 60967 2564 60979 2567
rect 61194 2564 61200 2576
rect 60967 2536 61200 2564
rect 60967 2533 60979 2536
rect 60921 2527 60979 2533
rect 61194 2524 61200 2536
rect 61252 2524 61258 2576
rect 61562 2524 61568 2576
rect 61620 2564 61626 2576
rect 61749 2567 61807 2573
rect 61749 2564 61761 2567
rect 61620 2536 61761 2564
rect 61620 2524 61626 2536
rect 61749 2533 61761 2536
rect 61795 2533 61807 2567
rect 61930 2564 61936 2576
rect 61891 2536 61936 2564
rect 61749 2527 61807 2533
rect 61930 2524 61936 2536
rect 61988 2524 61994 2576
rect 62853 2567 62911 2573
rect 62853 2533 62865 2567
rect 62899 2564 62911 2567
rect 63126 2564 63132 2576
rect 62899 2536 63132 2564
rect 62899 2533 62911 2536
rect 62853 2527 62911 2533
rect 63126 2524 63132 2536
rect 63184 2564 63190 2576
rect 63313 2567 63371 2573
rect 63313 2564 63325 2567
rect 63184 2536 63325 2564
rect 63184 2524 63190 2536
rect 63313 2533 63325 2536
rect 63359 2533 63371 2567
rect 63313 2527 63371 2533
rect 63589 2567 63647 2573
rect 63589 2533 63601 2567
rect 63635 2564 63647 2567
rect 63865 2567 63923 2573
rect 63865 2564 63877 2567
rect 63635 2536 63877 2564
rect 63635 2533 63647 2536
rect 63589 2527 63647 2533
rect 63865 2533 63877 2536
rect 63911 2564 63923 2567
rect 64046 2564 64052 2576
rect 63911 2536 64052 2564
rect 63911 2533 63923 2536
rect 63865 2527 63923 2533
rect 64046 2524 64052 2536
rect 64104 2524 64110 2576
rect 65521 2567 65579 2573
rect 65521 2533 65533 2567
rect 65567 2564 65579 2567
rect 65797 2567 65855 2573
rect 65797 2564 65809 2567
rect 65567 2536 65809 2564
rect 65567 2533 65579 2536
rect 65521 2527 65579 2533
rect 65797 2533 65809 2536
rect 65843 2564 65855 2567
rect 66070 2564 66076 2576
rect 65843 2536 66076 2564
rect 65843 2533 65855 2536
rect 65797 2527 65855 2533
rect 66070 2524 66076 2536
rect 66128 2524 66134 2576
rect 66548 2573 66576 2604
rect 68830 2592 68836 2604
rect 68888 2632 68894 2644
rect 68888 2604 69244 2632
rect 68888 2592 68894 2604
rect 66533 2567 66591 2573
rect 66533 2533 66545 2567
rect 66579 2533 66591 2567
rect 66533 2527 66591 2533
rect 67082 2524 67088 2576
rect 67140 2564 67146 2576
rect 67177 2567 67235 2573
rect 67177 2564 67189 2567
rect 67140 2536 67189 2564
rect 67140 2524 67146 2536
rect 67177 2533 67189 2536
rect 67223 2533 67235 2567
rect 68370 2564 68376 2576
rect 68331 2536 68376 2564
rect 67177 2527 67235 2533
rect 68370 2524 68376 2536
rect 68428 2524 68434 2576
rect 69216 2573 69244 2604
rect 69474 2592 69480 2644
rect 69532 2632 69538 2644
rect 69569 2635 69627 2641
rect 69569 2632 69581 2635
rect 69532 2604 69581 2632
rect 69532 2592 69538 2604
rect 69569 2601 69581 2604
rect 69615 2632 69627 2635
rect 70121 2635 70179 2641
rect 70121 2632 70133 2635
rect 69615 2604 70133 2632
rect 69615 2601 69627 2604
rect 69569 2595 69627 2601
rect 69952 2573 69980 2604
rect 70121 2601 70133 2604
rect 70167 2601 70179 2635
rect 70121 2595 70179 2601
rect 70670 2592 70676 2644
rect 70728 2632 70734 2644
rect 70765 2635 70823 2641
rect 70765 2632 70777 2635
rect 70728 2604 70777 2632
rect 70728 2592 70734 2604
rect 70765 2601 70777 2604
rect 70811 2632 70823 2635
rect 71498 2632 71504 2644
rect 70811 2604 71176 2632
rect 71459 2604 71504 2632
rect 70811 2601 70823 2604
rect 70765 2595 70823 2601
rect 71148 2573 71176 2604
rect 71498 2592 71504 2604
rect 71556 2632 71562 2644
rect 74166 2632 74172 2644
rect 71556 2604 71912 2632
rect 74127 2604 74172 2632
rect 71556 2592 71562 2604
rect 71884 2573 71912 2604
rect 74166 2592 74172 2604
rect 74224 2632 74230 2644
rect 74224 2604 74580 2632
rect 74224 2592 74230 2604
rect 69201 2567 69259 2573
rect 69201 2533 69213 2567
rect 69247 2533 69259 2567
rect 69201 2527 69259 2533
rect 69937 2567 69995 2573
rect 69937 2533 69949 2567
rect 69983 2533 69995 2567
rect 69937 2527 69995 2533
rect 71133 2567 71191 2573
rect 71133 2533 71145 2567
rect 71179 2533 71191 2567
rect 71133 2527 71191 2533
rect 71869 2567 71927 2573
rect 71869 2533 71881 2567
rect 71915 2533 71927 2567
rect 71869 2527 71927 2533
rect 72329 2567 72387 2573
rect 72329 2533 72341 2567
rect 72375 2564 72387 2567
rect 72510 2564 72516 2576
rect 72375 2536 72516 2564
rect 72375 2533 72387 2536
rect 72329 2527 72387 2533
rect 72510 2524 72516 2536
rect 72568 2564 72574 2576
rect 74552 2573 74580 2604
rect 74810 2592 74816 2644
rect 74868 2632 74874 2644
rect 74905 2635 74963 2641
rect 74905 2632 74917 2635
rect 74868 2604 74917 2632
rect 74868 2592 74874 2604
rect 74905 2601 74917 2604
rect 74951 2632 74963 2635
rect 74951 2604 75316 2632
rect 74951 2601 74963 2604
rect 74905 2595 74963 2601
rect 75288 2573 75316 2604
rect 77478 2592 77484 2644
rect 77536 2632 77542 2644
rect 77573 2635 77631 2641
rect 77573 2632 77585 2635
rect 77536 2604 77585 2632
rect 77536 2592 77542 2604
rect 77573 2601 77585 2604
rect 77619 2632 77631 2635
rect 78858 2632 78864 2644
rect 77619 2604 77984 2632
rect 78819 2604 78864 2632
rect 77619 2601 77631 2604
rect 77573 2595 77631 2601
rect 72605 2567 72663 2573
rect 72605 2564 72617 2567
rect 72568 2536 72617 2564
rect 72568 2524 72574 2536
rect 72605 2533 72617 2536
rect 72651 2564 72663 2567
rect 72789 2567 72847 2573
rect 72789 2564 72801 2567
rect 72651 2536 72801 2564
rect 72651 2533 72663 2536
rect 72605 2527 72663 2533
rect 72789 2533 72801 2536
rect 72835 2533 72847 2567
rect 74353 2567 74411 2573
rect 74353 2564 74365 2567
rect 72789 2527 72847 2533
rect 72896 2536 74365 2564
rect 41785 2499 41843 2505
rect 41785 2496 41797 2499
rect 41432 2468 41797 2496
rect 40405 2459 40463 2465
rect 41785 2465 41797 2468
rect 41831 2465 41843 2499
rect 44269 2499 44327 2505
rect 44269 2496 44281 2499
rect 41785 2459 41843 2465
rect 41892 2468 44281 2496
rect 26329 2431 26387 2437
rect 26329 2428 26341 2431
rect 25700 2400 26341 2428
rect 25593 2391 25651 2397
rect 26329 2397 26341 2400
rect 26375 2397 26387 2431
rect 26329 2391 26387 2397
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 31665 2431 31723 2437
rect 31665 2428 31677 2431
rect 30432 2400 31677 2428
rect 30432 2388 30438 2400
rect 31665 2397 31677 2400
rect 31711 2397 31723 2431
rect 31665 2391 31723 2397
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 34333 2431 34391 2437
rect 34333 2428 34345 2431
rect 32272 2400 34345 2428
rect 32272 2388 32278 2400
rect 34333 2397 34345 2400
rect 34379 2397 34391 2431
rect 34333 2391 34391 2397
rect 34606 2388 34612 2440
rect 34664 2428 34670 2440
rect 37737 2431 37795 2437
rect 37737 2428 37749 2431
rect 34664 2400 37749 2428
rect 34664 2388 34670 2400
rect 37737 2397 37749 2400
rect 37783 2397 37795 2431
rect 37737 2391 37795 2397
rect 38286 2388 38292 2440
rect 38344 2428 38350 2440
rect 41601 2431 41659 2437
rect 41601 2428 41613 2431
rect 38344 2400 41613 2428
rect 38344 2388 38350 2400
rect 41601 2397 41613 2400
rect 41647 2397 41659 2431
rect 41892 2428 41920 2468
rect 44269 2465 44281 2468
rect 44315 2465 44327 2499
rect 44269 2459 44327 2465
rect 46474 2456 46480 2508
rect 46532 2496 46538 2508
rect 47765 2499 47823 2505
rect 47765 2496 47777 2499
rect 46532 2468 47777 2496
rect 46532 2456 46538 2468
rect 47765 2465 47777 2468
rect 47811 2465 47823 2499
rect 47765 2459 47823 2465
rect 49878 2456 49884 2508
rect 49936 2496 49942 2508
rect 53009 2499 53067 2505
rect 53009 2496 53021 2499
rect 49936 2468 53021 2496
rect 49936 2456 49942 2468
rect 53009 2465 53021 2468
rect 53055 2465 53067 2499
rect 53009 2459 53067 2465
rect 54110 2456 54116 2508
rect 54168 2496 54174 2508
rect 57609 2499 57667 2505
rect 57609 2496 57621 2499
rect 54168 2468 57621 2496
rect 54168 2456 54174 2468
rect 57609 2465 57621 2468
rect 57655 2465 57667 2499
rect 57609 2459 57667 2465
rect 59354 2456 59360 2508
rect 59412 2496 59418 2508
rect 60277 2499 60335 2505
rect 60277 2496 60289 2499
rect 59412 2468 60289 2496
rect 59412 2456 59418 2468
rect 60277 2465 60289 2468
rect 60323 2465 60335 2499
rect 60277 2459 60335 2465
rect 62114 2456 62120 2508
rect 62172 2496 62178 2508
rect 62172 2468 63080 2496
rect 62172 2456 62178 2468
rect 41601 2391 41659 2397
rect 41800 2400 41920 2428
rect 5813 2363 5871 2369
rect 5813 2329 5825 2363
rect 5859 2360 5871 2363
rect 8938 2360 8944 2372
rect 5859 2332 8944 2360
rect 5859 2329 5871 2332
rect 5813 2323 5871 2329
rect 8938 2320 8944 2332
rect 8996 2320 9002 2372
rect 9858 2320 9864 2372
rect 9916 2360 9922 2372
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 9916 2332 13645 2360
rect 9916 2320 9922 2332
rect 13633 2329 13645 2332
rect 13679 2329 13691 2363
rect 13633 2323 13691 2329
rect 15286 2320 15292 2372
rect 15344 2360 15350 2372
rect 20533 2363 20591 2369
rect 20533 2360 20545 2363
rect 15344 2332 20545 2360
rect 15344 2320 15350 2332
rect 20533 2329 20545 2332
rect 20579 2329 20591 2363
rect 20533 2323 20591 2329
rect 21818 2320 21824 2372
rect 21876 2360 21882 2372
rect 22925 2363 22983 2369
rect 22925 2360 22937 2363
rect 21876 2332 22937 2360
rect 21876 2320 21882 2332
rect 22925 2329 22937 2332
rect 22971 2329 22983 2363
rect 22925 2323 22983 2329
rect 23014 2320 23020 2372
rect 23072 2360 23078 2372
rect 24673 2363 24731 2369
rect 24673 2360 24685 2363
rect 23072 2332 24685 2360
rect 23072 2320 23078 2332
rect 24673 2329 24685 2332
rect 24719 2329 24731 2363
rect 24673 2323 24731 2329
rect 24854 2320 24860 2372
rect 24912 2360 24918 2372
rect 27065 2363 27123 2369
rect 27065 2360 27077 2363
rect 24912 2332 27077 2360
rect 24912 2320 24918 2332
rect 27065 2329 27077 2332
rect 27111 2329 27123 2363
rect 27065 2323 27123 2329
rect 27890 2320 27896 2372
rect 27948 2360 27954 2372
rect 28261 2363 28319 2369
rect 28261 2360 28273 2363
rect 27948 2332 28273 2360
rect 27948 2320 27954 2332
rect 28261 2329 28273 2332
rect 28307 2329 28319 2363
rect 28261 2323 28319 2329
rect 28534 2320 28540 2372
rect 28592 2360 28598 2372
rect 28997 2363 29055 2369
rect 28997 2360 29009 2363
rect 28592 2332 29009 2360
rect 28592 2320 28598 2332
rect 28997 2329 29009 2332
rect 29043 2329 29055 2363
rect 28997 2323 29055 2329
rect 29086 2320 29092 2372
rect 29144 2360 29150 2372
rect 29733 2363 29791 2369
rect 29733 2360 29745 2363
rect 29144 2332 29745 2360
rect 29144 2320 29150 2332
rect 29733 2329 29745 2332
rect 29779 2329 29791 2363
rect 29733 2323 29791 2329
rect 29822 2320 29828 2372
rect 29880 2360 29886 2372
rect 30929 2363 30987 2369
rect 30929 2360 30941 2363
rect 29880 2332 30941 2360
rect 29880 2320 29886 2332
rect 30929 2329 30941 2332
rect 30975 2329 30987 2363
rect 30929 2323 30987 2329
rect 31018 2320 31024 2372
rect 31076 2360 31082 2372
rect 32401 2363 32459 2369
rect 32401 2360 32413 2363
rect 31076 2332 32413 2360
rect 31076 2320 31082 2332
rect 32401 2329 32413 2332
rect 32447 2329 32459 2363
rect 32401 2323 32459 2329
rect 32766 2320 32772 2372
rect 32824 2360 32830 2372
rect 32824 2332 33916 2360
rect 32824 2320 32830 2332
rect 8570 2252 8576 2304
rect 8628 2292 8634 2304
rect 11241 2295 11299 2301
rect 11241 2292 11253 2295
rect 8628 2264 11253 2292
rect 8628 2252 8634 2264
rect 11241 2261 11253 2264
rect 11287 2261 11299 2295
rect 11241 2255 11299 2261
rect 22462 2252 22468 2304
rect 22520 2292 22526 2304
rect 23753 2295 23811 2301
rect 23753 2292 23765 2295
rect 22520 2264 23765 2292
rect 22520 2252 22526 2264
rect 23753 2261 23765 2264
rect 23799 2261 23811 2295
rect 23753 2255 23811 2261
rect 31570 2252 31576 2304
rect 31628 2292 31634 2304
rect 33781 2295 33839 2301
rect 33781 2292 33793 2295
rect 31628 2264 33793 2292
rect 31628 2252 31634 2264
rect 33781 2261 33793 2264
rect 33827 2261 33839 2295
rect 33888 2292 33916 2332
rect 33962 2320 33968 2372
rect 34020 2360 34026 2372
rect 37001 2363 37059 2369
rect 37001 2360 37013 2363
rect 34020 2332 37013 2360
rect 34020 2320 34026 2332
rect 37001 2329 37013 2332
rect 37047 2329 37059 2363
rect 37001 2323 37059 2329
rect 38838 2320 38844 2372
rect 38896 2360 38902 2372
rect 38896 2332 40080 2360
rect 38896 2320 38902 2332
rect 35253 2295 35311 2301
rect 35253 2292 35265 2295
rect 33888 2264 35265 2292
rect 33781 2255 33839 2261
rect 35253 2261 35265 2264
rect 35299 2261 35311 2295
rect 35253 2255 35311 2261
rect 36446 2252 36452 2304
rect 36504 2292 36510 2304
rect 39761 2295 39819 2301
rect 39761 2292 39773 2295
rect 36504 2264 39773 2292
rect 36504 2252 36510 2264
rect 39761 2261 39773 2264
rect 39807 2261 39819 2295
rect 40052 2292 40080 2332
rect 40678 2320 40684 2372
rect 40736 2360 40742 2372
rect 41800 2360 41828 2400
rect 42518 2388 42524 2440
rect 42576 2428 42582 2440
rect 43070 2428 43076 2440
rect 42576 2400 42840 2428
rect 43031 2400 43076 2428
rect 42576 2388 42582 2400
rect 42613 2363 42671 2369
rect 42613 2360 42625 2363
rect 40736 2332 41828 2360
rect 41892 2332 42625 2360
rect 40736 2320 40742 2332
rect 41892 2292 41920 2332
rect 42613 2329 42625 2332
rect 42659 2329 42671 2363
rect 42812 2360 42840 2400
rect 43070 2388 43076 2400
rect 43128 2388 43134 2440
rect 43806 2388 43812 2440
rect 43864 2428 43870 2440
rect 47213 2431 47271 2437
rect 47213 2428 47225 2431
rect 43864 2400 47225 2428
rect 43864 2388 43870 2400
rect 47213 2397 47225 2400
rect 47259 2397 47271 2431
rect 47213 2391 47271 2397
rect 48038 2388 48044 2440
rect 48096 2428 48102 2440
rect 51077 2431 51135 2437
rect 51077 2428 51089 2431
rect 48096 2400 51089 2428
rect 48096 2388 48102 2400
rect 51077 2397 51089 2400
rect 51123 2397 51135 2431
rect 51077 2391 51135 2397
rect 51718 2388 51724 2440
rect 51776 2428 51782 2440
rect 54941 2431 54999 2437
rect 54941 2428 54953 2431
rect 51776 2400 54953 2428
rect 51776 2388 51782 2400
rect 54941 2397 54953 2400
rect 54987 2397 54999 2431
rect 54941 2391 54999 2397
rect 55030 2388 55036 2440
rect 55088 2428 55094 2440
rect 55953 2431 56011 2437
rect 55953 2428 55965 2431
rect 55088 2400 55965 2428
rect 55088 2388 55094 2400
rect 55953 2397 55965 2400
rect 55999 2397 56011 2431
rect 55953 2391 56011 2397
rect 59630 2388 59636 2440
rect 59688 2428 59694 2440
rect 62945 2431 63003 2437
rect 62945 2428 62957 2431
rect 59688 2400 62957 2428
rect 59688 2388 59694 2400
rect 62945 2397 62957 2400
rect 62991 2397 63003 2431
rect 63052 2428 63080 2468
rect 63402 2456 63408 2508
rect 63460 2496 63466 2508
rect 64509 2499 64567 2505
rect 64509 2496 64521 2499
rect 63460 2468 64521 2496
rect 63460 2456 63466 2468
rect 64509 2465 64521 2468
rect 64555 2465 64567 2499
rect 64509 2459 64567 2465
rect 66346 2456 66352 2508
rect 66404 2496 66410 2508
rect 69753 2499 69811 2505
rect 69753 2496 69765 2499
rect 66404 2468 69765 2496
rect 66404 2456 66410 2468
rect 69753 2465 69765 2468
rect 69799 2465 69811 2499
rect 69753 2459 69811 2465
rect 69842 2456 69848 2508
rect 69900 2496 69906 2508
rect 69900 2468 71084 2496
rect 69900 2456 69906 2468
rect 63681 2431 63739 2437
rect 63681 2428 63693 2431
rect 63052 2400 63693 2428
rect 62945 2391 63003 2397
rect 63681 2397 63693 2400
rect 63727 2397 63739 2431
rect 63681 2391 63739 2397
rect 63862 2388 63868 2440
rect 63920 2428 63926 2440
rect 67361 2431 67419 2437
rect 67361 2428 67373 2431
rect 63920 2400 67373 2428
rect 63920 2388 63926 2400
rect 67361 2397 67373 2400
rect 67407 2397 67419 2431
rect 67361 2391 67419 2397
rect 67542 2388 67548 2440
rect 67600 2428 67606 2440
rect 70949 2431 71007 2437
rect 70949 2428 70961 2431
rect 67600 2400 70961 2428
rect 67600 2388 67606 2400
rect 70949 2397 70961 2400
rect 70995 2397 71007 2431
rect 71056 2428 71084 2468
rect 71222 2456 71228 2508
rect 71280 2496 71286 2508
rect 72896 2496 72924 2536
rect 74353 2533 74365 2536
rect 74399 2533 74411 2567
rect 74353 2527 74411 2533
rect 74537 2567 74595 2573
rect 74537 2533 74549 2567
rect 74583 2533 74595 2567
rect 74537 2527 74595 2533
rect 75273 2567 75331 2573
rect 75273 2533 75285 2567
rect 75319 2533 75331 2567
rect 75273 2527 75331 2533
rect 76193 2567 76251 2573
rect 76193 2533 76205 2567
rect 76239 2564 76251 2567
rect 76469 2567 76527 2573
rect 76469 2564 76481 2567
rect 76239 2536 76481 2564
rect 76239 2533 76251 2536
rect 76193 2527 76251 2533
rect 76469 2533 76481 2536
rect 76515 2564 76527 2567
rect 76558 2564 76564 2576
rect 76515 2536 76564 2564
rect 76515 2533 76527 2536
rect 76469 2527 76527 2533
rect 76558 2524 76564 2536
rect 76616 2524 76622 2576
rect 76929 2567 76987 2573
rect 76929 2533 76941 2567
rect 76975 2564 76987 2567
rect 77202 2564 77208 2576
rect 76975 2536 77208 2564
rect 76975 2533 76987 2536
rect 76929 2527 76987 2533
rect 77202 2524 77208 2536
rect 77260 2524 77266 2576
rect 77294 2524 77300 2576
rect 77352 2564 77358 2576
rect 77956 2573 77984 2604
rect 78858 2592 78864 2604
rect 78916 2632 78922 2644
rect 79502 2632 79508 2644
rect 78916 2604 79180 2632
rect 79463 2604 79508 2632
rect 78916 2592 78922 2604
rect 79152 2573 79180 2604
rect 79502 2592 79508 2604
rect 79560 2632 79566 2644
rect 81529 2635 81587 2641
rect 79560 2604 79916 2632
rect 79560 2592 79566 2604
rect 79888 2573 79916 2604
rect 81529 2601 81541 2635
rect 81575 2632 81587 2635
rect 82081 2635 82139 2641
rect 82081 2632 82093 2635
rect 81575 2604 82093 2632
rect 81575 2601 81587 2604
rect 81529 2595 81587 2601
rect 77941 2567 77999 2573
rect 77352 2536 77892 2564
rect 77352 2524 77358 2536
rect 73706 2496 73712 2508
rect 71280 2468 72924 2496
rect 73667 2468 73712 2496
rect 71280 2456 71286 2468
rect 73706 2456 73712 2468
rect 73764 2456 73770 2508
rect 74258 2456 74264 2508
rect 74316 2496 74322 2508
rect 77757 2499 77815 2505
rect 77757 2496 77769 2499
rect 74316 2468 77769 2496
rect 74316 2456 74322 2468
rect 77757 2465 77769 2468
rect 77803 2465 77815 2499
rect 77864 2496 77892 2536
rect 77941 2533 77953 2567
rect 77987 2533 77999 2567
rect 77941 2527 77999 2533
rect 79137 2567 79195 2573
rect 79137 2533 79149 2567
rect 79183 2533 79195 2567
rect 79137 2527 79195 2533
rect 79873 2567 79931 2573
rect 79873 2533 79885 2567
rect 79919 2533 79931 2567
rect 79873 2527 79931 2533
rect 80517 2567 80575 2573
rect 80517 2533 80529 2567
rect 80563 2564 80575 2567
rect 80606 2564 80612 2576
rect 80563 2536 80612 2564
rect 80563 2533 80575 2536
rect 80517 2527 80575 2533
rect 80606 2524 80612 2536
rect 80664 2524 80670 2576
rect 81820 2573 81848 2604
rect 82081 2601 82093 2604
rect 82127 2632 82139 2635
rect 82722 2632 82728 2644
rect 82127 2604 82728 2632
rect 82127 2601 82139 2604
rect 82081 2595 82139 2601
rect 82722 2592 82728 2604
rect 82780 2592 82786 2644
rect 84562 2592 84568 2644
rect 84620 2632 84626 2644
rect 84749 2635 84807 2641
rect 84749 2632 84761 2635
rect 84620 2604 84761 2632
rect 84620 2592 84626 2604
rect 84749 2601 84761 2604
rect 84795 2632 84807 2635
rect 84841 2635 84899 2641
rect 84841 2632 84853 2635
rect 84795 2604 84853 2632
rect 84795 2601 84807 2604
rect 84749 2595 84807 2601
rect 84841 2601 84853 2604
rect 84887 2601 84899 2635
rect 88334 2632 88340 2644
rect 88295 2604 88340 2632
rect 84841 2595 84899 2601
rect 88334 2592 88340 2604
rect 88392 2632 88398 2644
rect 89438 2632 89444 2644
rect 88392 2604 88656 2632
rect 89399 2604 89444 2632
rect 88392 2592 88398 2604
rect 81805 2567 81863 2573
rect 81805 2533 81817 2567
rect 81851 2533 81863 2567
rect 81805 2527 81863 2533
rect 82814 2524 82820 2576
rect 82872 2564 82878 2576
rect 82909 2567 82967 2573
rect 82909 2564 82921 2567
rect 82872 2536 82921 2564
rect 82872 2524 82878 2536
rect 82909 2533 82921 2536
rect 82955 2533 82967 2567
rect 82909 2527 82967 2533
rect 84381 2567 84439 2573
rect 84381 2533 84393 2567
rect 84427 2564 84439 2567
rect 85574 2564 85580 2576
rect 84427 2536 85580 2564
rect 84427 2533 84439 2536
rect 84381 2527 84439 2533
rect 85574 2524 85580 2536
rect 85632 2524 85638 2576
rect 85669 2567 85727 2573
rect 85669 2533 85681 2567
rect 85715 2564 85727 2567
rect 85942 2564 85948 2576
rect 85715 2536 85948 2564
rect 85715 2533 85727 2536
rect 85669 2527 85727 2533
rect 85942 2524 85948 2536
rect 86000 2524 86006 2576
rect 86954 2524 86960 2576
rect 87012 2564 87018 2576
rect 87049 2567 87107 2573
rect 87049 2564 87061 2567
rect 87012 2536 87061 2564
rect 87012 2524 87018 2536
rect 87049 2533 87061 2536
rect 87095 2533 87107 2567
rect 87049 2527 87107 2533
rect 87601 2567 87659 2573
rect 87601 2533 87613 2567
rect 87647 2564 87659 2567
rect 87874 2564 87880 2576
rect 87647 2536 87880 2564
rect 87647 2533 87659 2536
rect 87601 2527 87659 2533
rect 87874 2524 87880 2536
rect 87932 2524 87938 2576
rect 88628 2573 88656 2604
rect 89438 2592 89444 2604
rect 89496 2632 89502 2644
rect 89993 2635 90051 2641
rect 89993 2632 90005 2635
rect 89496 2604 90005 2632
rect 89496 2592 89502 2604
rect 88613 2567 88671 2573
rect 88613 2533 88625 2567
rect 88659 2533 88671 2567
rect 89622 2564 89628 2576
rect 89583 2536 89628 2564
rect 88613 2527 88671 2533
rect 89622 2524 89628 2536
rect 89680 2524 89686 2576
rect 89824 2573 89852 2604
rect 89993 2601 90005 2604
rect 90039 2601 90051 2635
rect 90726 2632 90732 2644
rect 90687 2604 90732 2632
rect 89993 2595 90051 2601
rect 90726 2592 90732 2604
rect 90784 2592 90790 2644
rect 91370 2592 91376 2644
rect 91428 2632 91434 2644
rect 92109 2635 92167 2641
rect 92109 2632 92121 2635
rect 91428 2604 92121 2632
rect 91428 2592 91434 2604
rect 92109 2601 92121 2604
rect 92155 2632 92167 2635
rect 92842 2632 92848 2644
rect 92155 2604 92520 2632
rect 92803 2604 92848 2632
rect 92155 2601 92167 2604
rect 92109 2595 92167 2601
rect 89809 2567 89867 2573
rect 89809 2533 89821 2567
rect 89855 2533 89867 2567
rect 89809 2527 89867 2533
rect 90269 2567 90327 2573
rect 90269 2533 90281 2567
rect 90315 2564 90327 2567
rect 90545 2567 90603 2573
rect 90545 2564 90557 2567
rect 90315 2536 90557 2564
rect 90315 2533 90327 2536
rect 90269 2527 90327 2533
rect 90545 2533 90557 2536
rect 90591 2564 90603 2567
rect 90744 2564 90772 2592
rect 90591 2536 90772 2564
rect 91189 2567 91247 2573
rect 90591 2533 90603 2536
rect 90545 2527 90603 2533
rect 91189 2533 91201 2567
rect 91235 2564 91247 2567
rect 91462 2564 91468 2576
rect 91235 2536 91468 2564
rect 91235 2533 91247 2536
rect 91189 2527 91247 2533
rect 91462 2524 91468 2536
rect 91520 2524 91526 2576
rect 92492 2573 92520 2604
rect 92842 2592 92848 2604
rect 92900 2632 92906 2644
rect 92900 2604 93256 2632
rect 92900 2592 92906 2604
rect 93228 2573 93256 2604
rect 94314 2592 94320 2644
rect 94372 2632 94378 2644
rect 94777 2635 94835 2641
rect 94777 2632 94789 2635
rect 94372 2604 94789 2632
rect 94372 2592 94378 2604
rect 94777 2601 94789 2604
rect 94823 2632 94835 2635
rect 95510 2632 95516 2644
rect 94823 2604 95188 2632
rect 95471 2604 95516 2632
rect 94823 2601 94835 2604
rect 94777 2595 94835 2601
rect 92477 2567 92535 2573
rect 92477 2533 92489 2567
rect 92523 2533 92535 2567
rect 92477 2527 92535 2533
rect 93213 2567 93271 2573
rect 93213 2533 93225 2567
rect 93259 2533 93271 2567
rect 93213 2527 93271 2533
rect 93673 2567 93731 2573
rect 93673 2533 93685 2567
rect 93719 2564 93731 2567
rect 93854 2564 93860 2576
rect 93719 2536 93860 2564
rect 93719 2533 93731 2536
rect 93673 2527 93731 2533
rect 93854 2524 93860 2536
rect 93912 2564 93918 2576
rect 95160 2573 95188 2604
rect 95510 2592 95516 2604
rect 95568 2632 95574 2644
rect 95568 2604 95924 2632
rect 95568 2592 95574 2604
rect 95896 2573 95924 2604
rect 96154 2592 96160 2644
rect 96212 2632 96218 2644
rect 96249 2635 96307 2641
rect 96249 2632 96261 2635
rect 96212 2604 96261 2632
rect 96212 2592 96218 2604
rect 96249 2601 96261 2604
rect 96295 2632 96307 2635
rect 96295 2604 96568 2632
rect 96295 2601 96307 2604
rect 96249 2595 96307 2601
rect 96540 2573 96568 2604
rect 93949 2567 94007 2573
rect 93949 2564 93961 2567
rect 93912 2536 93961 2564
rect 93912 2524 93918 2536
rect 93949 2533 93961 2536
rect 93995 2533 94007 2567
rect 93949 2527 94007 2533
rect 95145 2567 95203 2573
rect 95145 2533 95157 2567
rect 95191 2533 95203 2567
rect 95145 2527 95203 2533
rect 95881 2567 95939 2573
rect 95881 2533 95893 2567
rect 95927 2533 95939 2567
rect 95881 2527 95939 2533
rect 96525 2567 96583 2573
rect 96525 2533 96537 2567
rect 96571 2533 96583 2567
rect 96525 2527 96583 2533
rect 96709 2567 96767 2573
rect 96709 2533 96721 2567
rect 96755 2564 96767 2567
rect 97718 2564 97724 2576
rect 96755 2536 97724 2564
rect 96755 2533 96767 2536
rect 96709 2527 96767 2533
rect 97718 2524 97724 2536
rect 97776 2524 97782 2576
rect 79689 2499 79747 2505
rect 79689 2496 79701 2499
rect 77864 2468 79701 2496
rect 77757 2459 77815 2465
rect 79689 2465 79701 2468
rect 79735 2465 79747 2499
rect 79689 2459 79747 2465
rect 84749 2499 84807 2505
rect 84749 2465 84761 2499
rect 84795 2496 84807 2499
rect 85209 2499 85267 2505
rect 85209 2496 85221 2499
rect 84795 2468 85221 2496
rect 84795 2465 84807 2468
rect 84749 2459 84807 2465
rect 85209 2465 85221 2468
rect 85255 2465 85267 2499
rect 85209 2459 85267 2465
rect 95694 2456 95700 2508
rect 95752 2496 95758 2508
rect 97629 2499 97687 2505
rect 97629 2496 97641 2499
rect 95752 2468 97641 2496
rect 95752 2456 95758 2468
rect 97629 2465 97641 2468
rect 97675 2496 97687 2499
rect 97905 2499 97963 2505
rect 97905 2496 97917 2499
rect 97675 2468 97917 2496
rect 97675 2465 97687 2468
rect 97629 2459 97687 2465
rect 97905 2465 97917 2468
rect 97951 2465 97963 2499
rect 97905 2459 97963 2465
rect 72421 2431 72479 2437
rect 72421 2428 72433 2431
rect 71056 2400 72433 2428
rect 70949 2391 71007 2397
rect 72421 2397 72433 2400
rect 72467 2397 72479 2431
rect 72421 2391 72479 2397
rect 73062 2388 73068 2440
rect 73120 2428 73126 2440
rect 76285 2431 76343 2437
rect 76285 2428 76297 2431
rect 73120 2400 76297 2428
rect 73120 2388 73126 2400
rect 76285 2397 76297 2400
rect 76331 2397 76343 2431
rect 76285 2391 76343 2397
rect 77294 2388 77300 2440
rect 77352 2428 77358 2440
rect 80701 2431 80759 2437
rect 80701 2428 80713 2431
rect 77352 2400 80713 2428
rect 77352 2388 77358 2400
rect 80701 2397 80713 2400
rect 80747 2397 80759 2431
rect 80701 2391 80759 2397
rect 81158 2388 81164 2440
rect 81216 2428 81222 2440
rect 81342 2428 81348 2440
rect 81216 2400 81348 2428
rect 81216 2388 81222 2400
rect 81342 2388 81348 2400
rect 81400 2388 81406 2440
rect 84654 2388 84660 2440
rect 84712 2428 84718 2440
rect 85761 2431 85819 2437
rect 85761 2428 85773 2431
rect 84712 2400 85773 2428
rect 84712 2388 84718 2400
rect 85761 2397 85773 2400
rect 85807 2397 85819 2431
rect 85761 2391 85819 2397
rect 86402 2388 86408 2440
rect 86460 2428 86466 2440
rect 88429 2431 88487 2437
rect 88429 2428 88441 2431
rect 86460 2400 88441 2428
rect 86460 2388 86466 2400
rect 88429 2397 88441 2400
rect 88475 2397 88487 2431
rect 90361 2431 90419 2437
rect 90361 2428 90373 2431
rect 88429 2391 88487 2397
rect 89824 2400 90373 2428
rect 45741 2363 45799 2369
rect 45741 2360 45753 2363
rect 42812 2332 45753 2360
rect 42613 2323 42671 2329
rect 45741 2329 45753 2332
rect 45787 2329 45799 2363
rect 45741 2323 45799 2329
rect 46198 2320 46204 2372
rect 46256 2360 46262 2372
rect 49605 2363 49663 2369
rect 49605 2360 49617 2363
rect 46256 2332 49617 2360
rect 46256 2320 46262 2332
rect 49605 2329 49617 2332
rect 49651 2329 49663 2363
rect 49605 2323 49663 2329
rect 51184 2332 52592 2360
rect 40052 2264 41920 2292
rect 39761 2255 39819 2261
rect 41966 2252 41972 2304
rect 42024 2292 42030 2304
rect 45189 2295 45247 2301
rect 45189 2292 45201 2295
rect 42024 2264 45201 2292
rect 42024 2252 42030 2264
rect 45189 2261 45201 2264
rect 45235 2261 45247 2295
rect 45189 2255 45247 2261
rect 46106 2252 46112 2304
rect 46164 2292 46170 2304
rect 47857 2295 47915 2301
rect 47857 2292 47869 2295
rect 46164 2264 47869 2292
rect 46164 2252 46170 2264
rect 47857 2261 47869 2264
rect 47903 2261 47915 2295
rect 47857 2255 47915 2261
rect 47946 2252 47952 2304
rect 48004 2292 48010 2304
rect 50433 2295 50491 2301
rect 50433 2292 50445 2295
rect 48004 2264 50445 2292
rect 48004 2252 48010 2264
rect 50433 2261 50445 2264
rect 50479 2261 50491 2295
rect 50433 2255 50491 2261
rect 50522 2252 50528 2304
rect 50580 2292 50586 2304
rect 51184 2292 51212 2332
rect 50580 2264 51212 2292
rect 50580 2252 50586 2264
rect 51534 2252 51540 2304
rect 51592 2292 51598 2304
rect 52457 2295 52515 2301
rect 52457 2292 52469 2295
rect 51592 2264 52469 2292
rect 51592 2252 51598 2264
rect 52457 2261 52469 2264
rect 52503 2261 52515 2295
rect 52564 2292 52592 2332
rect 52914 2320 52920 2372
rect 52972 2360 52978 2372
rect 56413 2363 56471 2369
rect 56413 2360 56425 2363
rect 52972 2332 56425 2360
rect 52972 2320 52978 2332
rect 56413 2329 56425 2332
rect 56459 2329 56471 2363
rect 56413 2323 56471 2329
rect 57790 2320 57796 2372
rect 57848 2360 57854 2372
rect 61013 2363 61071 2369
rect 61013 2360 61025 2363
rect 57848 2332 61025 2360
rect 57848 2320 57854 2332
rect 61013 2329 61025 2332
rect 61059 2329 61071 2363
rect 61013 2323 61071 2329
rect 61212 2332 62160 2360
rect 53929 2295 53987 2301
rect 53929 2292 53941 2295
rect 52564 2264 53941 2292
rect 52457 2255 52515 2261
rect 53929 2261 53941 2264
rect 53975 2261 53987 2295
rect 53929 2255 53987 2261
rect 55950 2252 55956 2304
rect 56008 2292 56014 2304
rect 59173 2295 59231 2301
rect 59173 2292 59185 2295
rect 56008 2264 59185 2292
rect 56008 2252 56014 2264
rect 59173 2261 59185 2264
rect 59219 2261 59231 2295
rect 59173 2255 59231 2261
rect 60826 2252 60832 2304
rect 60884 2292 60890 2304
rect 61212 2292 61240 2332
rect 60884 2264 61240 2292
rect 62132 2292 62160 2332
rect 63310 2320 63316 2372
rect 63368 2360 63374 2372
rect 66349 2363 66407 2369
rect 66349 2360 66361 2363
rect 63368 2332 66361 2360
rect 63368 2320 63374 2332
rect 66349 2329 66361 2332
rect 66395 2329 66407 2363
rect 66349 2323 66407 2329
rect 66438 2320 66444 2372
rect 66496 2360 66502 2372
rect 69017 2363 69075 2369
rect 69017 2360 69029 2363
rect 66496 2332 69029 2360
rect 66496 2320 66502 2332
rect 69017 2329 69029 2332
rect 69063 2329 69075 2363
rect 69017 2323 69075 2329
rect 69106 2320 69112 2372
rect 69164 2360 69170 2372
rect 71685 2363 71743 2369
rect 71685 2360 71697 2363
rect 69164 2332 71697 2360
rect 69164 2320 69170 2332
rect 71685 2329 71697 2332
rect 71731 2329 71743 2363
rect 71685 2323 71743 2329
rect 71866 2320 71872 2372
rect 71924 2360 71930 2372
rect 75089 2363 75147 2369
rect 75089 2360 75101 2363
rect 71924 2332 75101 2360
rect 71924 2320 71930 2332
rect 75089 2329 75101 2332
rect 75135 2329 75147 2363
rect 75089 2323 75147 2329
rect 75454 2320 75460 2372
rect 75512 2360 75518 2372
rect 75512 2332 77248 2360
rect 75512 2320 75518 2332
rect 64601 2295 64659 2301
rect 64601 2292 64613 2295
rect 62132 2264 64613 2292
rect 60884 2252 60890 2264
rect 64601 2261 64613 2264
rect 64647 2261 64659 2295
rect 64601 2255 64659 2261
rect 65058 2252 65064 2304
rect 65116 2292 65122 2304
rect 68465 2295 68523 2301
rect 68465 2292 68477 2295
rect 65116 2264 68477 2292
rect 65116 2252 65122 2264
rect 68465 2261 68477 2264
rect 68511 2261 68523 2295
rect 68465 2255 68523 2261
rect 70026 2252 70032 2304
rect 70084 2292 70090 2304
rect 73801 2295 73859 2301
rect 73801 2292 73813 2295
rect 70084 2264 73813 2292
rect 70084 2252 70090 2264
rect 73801 2261 73813 2264
rect 73847 2261 73859 2295
rect 73801 2255 73859 2261
rect 74718 2252 74724 2304
rect 74776 2292 74782 2304
rect 77113 2295 77171 2301
rect 77113 2292 77125 2295
rect 74776 2264 77125 2292
rect 74776 2252 74782 2264
rect 77113 2261 77125 2264
rect 77159 2261 77171 2295
rect 77220 2292 77248 2332
rect 78490 2320 78496 2372
rect 78548 2360 78554 2372
rect 81621 2363 81679 2369
rect 81621 2360 81633 2363
rect 78548 2332 81633 2360
rect 78548 2320 78554 2332
rect 81621 2329 81633 2332
rect 81667 2329 81679 2363
rect 81621 2323 81679 2329
rect 84010 2320 84016 2372
rect 84068 2360 84074 2372
rect 85025 2363 85083 2369
rect 85025 2360 85037 2363
rect 84068 2332 85037 2360
rect 84068 2320 84074 2332
rect 85025 2329 85037 2332
rect 85071 2329 85083 2363
rect 85025 2323 85083 2329
rect 85850 2320 85856 2372
rect 85908 2360 85914 2372
rect 87693 2363 87751 2369
rect 87693 2360 87705 2363
rect 85908 2332 87705 2360
rect 85908 2320 85914 2332
rect 87693 2329 87705 2332
rect 87739 2329 87751 2363
rect 87693 2323 87751 2329
rect 87782 2320 87788 2372
rect 87840 2360 87846 2372
rect 89824 2360 89852 2400
rect 90361 2397 90373 2400
rect 90407 2397 90419 2431
rect 91373 2431 91431 2437
rect 91373 2428 91385 2431
rect 90361 2391 90419 2397
rect 90468 2400 91385 2428
rect 87840 2332 89852 2360
rect 87840 2320 87846 2332
rect 79045 2295 79103 2301
rect 79045 2292 79057 2295
rect 77220 2264 79057 2292
rect 77113 2255 77171 2261
rect 79045 2261 79057 2264
rect 79091 2261 79103 2295
rect 79045 2255 79103 2261
rect 82814 2252 82820 2304
rect 82872 2292 82878 2304
rect 83001 2295 83059 2301
rect 83001 2292 83013 2295
rect 82872 2264 83013 2292
rect 82872 2252 82878 2264
rect 83001 2261 83013 2264
rect 83047 2261 83059 2295
rect 83001 2255 83059 2261
rect 83366 2252 83372 2304
rect 83424 2292 83430 2304
rect 84473 2295 84531 2301
rect 84473 2292 84485 2295
rect 83424 2264 84485 2292
rect 83424 2252 83430 2264
rect 84473 2261 84485 2264
rect 84519 2261 84531 2295
rect 84473 2255 84531 2261
rect 85206 2252 85212 2304
rect 85264 2292 85270 2304
rect 87141 2295 87199 2301
rect 87141 2292 87153 2295
rect 85264 2264 87153 2292
rect 85264 2252 85270 2264
rect 87141 2261 87153 2264
rect 87187 2261 87199 2295
rect 87141 2255 87199 2261
rect 88242 2252 88248 2304
rect 88300 2292 88306 2304
rect 90468 2292 90496 2400
rect 91373 2397 91385 2400
rect 91419 2397 91431 2431
rect 91373 2391 91431 2397
rect 91922 2388 91928 2440
rect 91980 2428 91986 2440
rect 94961 2431 95019 2437
rect 94961 2428 94973 2431
rect 91980 2400 94973 2428
rect 91980 2388 91986 2400
rect 94961 2397 94973 2400
rect 95007 2397 95019 2431
rect 94961 2391 95019 2397
rect 91002 2320 91008 2372
rect 91060 2360 91066 2372
rect 92293 2363 92351 2369
rect 92293 2360 92305 2363
rect 91060 2332 92305 2360
rect 91060 2320 91066 2332
rect 92293 2329 92305 2332
rect 92339 2329 92351 2363
rect 93026 2360 93032 2372
rect 92987 2332 93032 2360
rect 92293 2323 92351 2329
rect 93026 2320 93032 2332
rect 93084 2320 93090 2372
rect 93765 2363 93823 2369
rect 93765 2329 93777 2363
rect 93811 2329 93823 2363
rect 93765 2323 93823 2329
rect 88300 2264 90496 2292
rect 88300 2252 88306 2264
rect 90726 2252 90732 2304
rect 90784 2292 90790 2304
rect 93780 2292 93808 2323
rect 94222 2320 94228 2372
rect 94280 2360 94286 2372
rect 95697 2363 95755 2369
rect 95697 2360 95709 2363
rect 94280 2332 95709 2360
rect 94280 2320 94286 2332
rect 95697 2329 95709 2332
rect 95743 2329 95755 2363
rect 95697 2323 95755 2329
rect 98089 2363 98147 2369
rect 98089 2329 98101 2363
rect 98135 2360 98147 2363
rect 99650 2360 99656 2372
rect 98135 2332 99656 2360
rect 98135 2329 98147 2332
rect 98089 2323 98147 2329
rect 99650 2320 99656 2332
rect 99708 2320 99714 2372
rect 90784 2264 93808 2292
rect 90784 2252 90790 2264
rect 1104 2202 98808 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 65686 2202
rect 65738 2150 65750 2202
rect 65802 2150 65814 2202
rect 65866 2150 65878 2202
rect 65930 2150 96406 2202
rect 96458 2150 96470 2202
rect 96522 2150 96534 2202
rect 96586 2150 96598 2202
rect 96650 2150 98808 2202
rect 1104 2128 98808 2150
rect 35986 2048 35992 2100
rect 36044 2088 36050 2100
rect 45646 2088 45652 2100
rect 36044 2060 45652 2088
rect 36044 2048 36050 2060
rect 45646 2048 45652 2060
rect 45704 2048 45710 2100
rect 48682 2048 48688 2100
rect 48740 2088 48746 2100
rect 51534 2088 51540 2100
rect 48740 2060 51540 2088
rect 48740 2048 48746 2060
rect 51534 2048 51540 2060
rect 51592 2048 51598 2100
rect 52270 2048 52276 2100
rect 52328 2088 52334 2100
rect 55030 2088 55036 2100
rect 52328 2060 55036 2088
rect 52328 2048 52334 2060
rect 55030 2048 55036 2060
rect 55088 2048 55094 2100
rect 88886 2048 88892 2100
rect 88944 2088 88950 2100
rect 91002 2088 91008 2100
rect 88944 2060 91008 2088
rect 88944 2048 88950 2060
rect 91002 2048 91008 2060
rect 91060 2048 91066 2100
rect 4338 1844 4344 1896
rect 4396 1884 4402 1896
rect 4798 1884 4804 1896
rect 4396 1856 4804 1884
rect 4396 1844 4402 1856
rect 4798 1844 4804 1856
rect 4856 1844 4862 1896
rect 19794 1844 19800 1896
rect 19852 1884 19858 1896
rect 20070 1884 20076 1896
rect 19852 1856 20076 1884
rect 19852 1844 19858 1856
rect 20070 1844 20076 1856
rect 20128 1844 20134 1896
rect 35066 1504 35072 1556
rect 35124 1544 35130 1556
rect 35342 1544 35348 1556
rect 35124 1516 35348 1544
rect 35124 1504 35130 1516
rect 35342 1504 35348 1516
rect 35400 1504 35406 1556
rect 68738 1436 68744 1488
rect 68796 1476 68802 1488
rect 69842 1476 69848 1488
rect 68796 1448 69848 1476
rect 68796 1436 68802 1448
rect 69842 1436 69848 1448
rect 69900 1436 69906 1488
rect 4522 1368 4528 1420
rect 4580 1408 4586 1420
rect 5626 1408 5632 1420
rect 4580 1380 5632 1408
rect 4580 1368 4586 1380
rect 5626 1368 5632 1380
rect 5684 1368 5690 1420
rect 44358 1368 44364 1420
rect 44416 1408 44422 1420
rect 46106 1408 46112 1420
rect 44416 1380 46112 1408
rect 44416 1368 44422 1380
rect 46106 1368 46112 1380
rect 46164 1368 46170 1420
rect 46842 1368 46848 1420
rect 46900 1408 46906 1420
rect 47946 1408 47952 1420
rect 46900 1380 47952 1408
rect 46900 1368 46906 1380
rect 47946 1368 47952 1380
rect 48004 1368 48010 1420
rect 65702 1368 65708 1420
rect 65760 1408 65766 1420
rect 66438 1408 66444 1420
rect 65760 1380 66444 1408
rect 65760 1368 65766 1380
rect 66438 1368 66444 1380
rect 66496 1368 66502 1420
rect 68186 1368 68192 1420
rect 68244 1408 68250 1420
rect 69106 1408 69112 1420
rect 68244 1380 69112 1408
rect 68244 1368 68250 1380
rect 69106 1368 69112 1380
rect 69164 1368 69170 1420
rect 92566 1368 92572 1420
rect 92624 1408 92630 1420
rect 94222 1408 94228 1420
rect 92624 1380 94228 1408
rect 92624 1368 92630 1380
rect 94222 1368 94228 1380
rect 94280 1368 94286 1420
rect 3970 1300 3976 1352
rect 4028 1340 4034 1352
rect 49786 1340 49792 1352
rect 4028 1312 49792 1340
rect 4028 1300 4034 1312
rect 49786 1300 49792 1312
rect 49844 1340 49850 1352
rect 84286 1340 84292 1352
rect 49844 1312 84292 1340
rect 49844 1300 49850 1312
rect 84286 1300 84292 1312
rect 84344 1300 84350 1352
rect 39482 1164 39488 1216
rect 39540 1204 39546 1216
rect 43070 1204 43076 1216
rect 39540 1176 43076 1204
rect 39540 1164 39546 1176
rect 43070 1164 43076 1176
rect 43128 1164 43134 1216
rect 89530 1164 89536 1216
rect 89588 1204 89594 1216
rect 93026 1204 93032 1216
rect 89588 1176 93032 1204
rect 89588 1164 89594 1176
rect 93026 1164 93032 1176
rect 93084 1164 93090 1216
<< via1 >>
rect 16304 97588 16356 97640
rect 90456 97588 90508 97640
rect 23940 97520 23992 97572
rect 56508 97520 56560 97572
rect 7656 97452 7708 97504
rect 68560 97452 68612 97504
rect 19606 97350 19658 97402
rect 19670 97350 19722 97402
rect 19734 97350 19786 97402
rect 19798 97350 19850 97402
rect 50326 97350 50378 97402
rect 50390 97350 50442 97402
rect 50454 97350 50506 97402
rect 50518 97350 50570 97402
rect 81046 97350 81098 97402
rect 81110 97350 81162 97402
rect 81174 97350 81226 97402
rect 81238 97350 81290 97402
rect 1216 97248 1268 97300
rect 3792 97248 3844 97300
rect 6460 97248 6512 97300
rect 9036 97248 9088 97300
rect 11612 97248 11664 97300
rect 2964 97223 3016 97232
rect 2964 97189 2973 97223
rect 2973 97189 3007 97223
rect 3007 97189 3016 97223
rect 2964 97180 3016 97189
rect 6184 97180 6236 97232
rect 10784 97180 10836 97232
rect 388 97112 440 97164
rect 2504 97112 2556 97164
rect 5540 97155 5592 97164
rect 5540 97121 5549 97155
rect 5549 97121 5583 97155
rect 5583 97121 5592 97155
rect 5540 97112 5592 97121
rect 7012 97155 7064 97164
rect 7012 97121 7021 97155
rect 7021 97121 7055 97155
rect 7055 97121 7064 97155
rect 7012 97112 7064 97121
rect 8208 97155 8260 97164
rect 8208 97121 8217 97155
rect 8217 97121 8251 97155
rect 8251 97121 8260 97155
rect 8208 97112 8260 97121
rect 14280 97180 14332 97232
rect 16028 97180 16080 97232
rect 16856 97248 16908 97300
rect 19432 97248 19484 97300
rect 22100 97248 22152 97300
rect 12348 97155 12400 97164
rect 12348 97121 12357 97155
rect 12357 97121 12391 97155
rect 12391 97121 12400 97155
rect 12348 97112 12400 97121
rect 13360 97155 13412 97164
rect 13360 97121 13369 97155
rect 13369 97121 13403 97155
rect 13403 97121 13412 97155
rect 13360 97112 13412 97121
rect 15016 97155 15068 97164
rect 15016 97121 15025 97155
rect 15025 97121 15059 97155
rect 15059 97121 15068 97155
rect 15016 97112 15068 97121
rect 17684 97155 17736 97164
rect 17684 97121 17693 97155
rect 17693 97121 17727 97155
rect 17727 97121 17736 97155
rect 17684 97112 17736 97121
rect 18604 97180 18656 97232
rect 21456 97180 21508 97232
rect 22836 97180 22888 97232
rect 23940 97180 23992 97232
rect 24676 97223 24728 97232
rect 24676 97189 24685 97223
rect 24685 97189 24719 97223
rect 24719 97189 24728 97223
rect 24676 97180 24728 97189
rect 26424 97180 26476 97232
rect 27344 97248 27396 97300
rect 29920 97291 29972 97300
rect 29920 97257 29929 97291
rect 29929 97257 29963 97291
rect 29963 97257 29972 97291
rect 29920 97248 29972 97257
rect 30748 97248 30800 97300
rect 32496 97248 32548 97300
rect 20352 97155 20404 97164
rect 20352 97121 20361 97155
rect 20361 97121 20395 97155
rect 20395 97121 20404 97155
rect 20352 97112 20404 97121
rect 21180 97155 21232 97164
rect 21180 97121 21189 97155
rect 21189 97121 21223 97155
rect 21223 97121 21232 97155
rect 21180 97112 21232 97121
rect 23112 97112 23164 97164
rect 24492 97155 24544 97164
rect 24492 97121 24501 97155
rect 24501 97121 24535 97155
rect 24535 97121 24544 97155
rect 24492 97112 24544 97121
rect 26056 97112 26108 97164
rect 28264 97112 28316 97164
rect 5724 97087 5776 97096
rect 5724 97053 5733 97087
rect 5733 97053 5767 97087
rect 5767 97053 5776 97087
rect 5724 97044 5776 97053
rect 8760 97044 8812 97096
rect 14832 97044 14884 97096
rect 21364 97087 21416 97096
rect 21364 97053 21373 97087
rect 21373 97053 21407 97087
rect 21407 97053 21416 97087
rect 21364 97044 21416 97053
rect 28172 97044 28224 97096
rect 29000 97180 29052 97232
rect 31760 97223 31812 97232
rect 31760 97189 31769 97223
rect 31769 97189 31803 97223
rect 31803 97189 31812 97223
rect 31760 97180 31812 97189
rect 29828 97155 29880 97164
rect 29828 97121 29837 97155
rect 29837 97121 29871 97155
rect 29871 97121 29880 97155
rect 29828 97112 29880 97121
rect 31024 97155 31076 97164
rect 31024 97121 31033 97155
rect 31033 97121 31067 97155
rect 31067 97121 31076 97155
rect 31024 97112 31076 97121
rect 32496 97155 32548 97164
rect 32496 97121 32505 97155
rect 32505 97121 32539 97155
rect 32539 97121 32548 97155
rect 32496 97112 32548 97121
rect 34244 97155 34296 97164
rect 34244 97121 34253 97155
rect 34253 97121 34287 97155
rect 34287 97121 34296 97155
rect 34244 97112 34296 97121
rect 35164 97248 35216 97300
rect 37740 97248 37792 97300
rect 40316 97248 40368 97300
rect 42984 97248 43036 97300
rect 90456 97291 90508 97300
rect 36820 97180 36872 97232
rect 39488 97180 39540 97232
rect 42064 97180 42116 97232
rect 34796 97112 34848 97164
rect 37832 97155 37884 97164
rect 37832 97121 37841 97155
rect 37841 97121 37875 97155
rect 37875 97121 37884 97155
rect 37832 97112 37884 97121
rect 40500 97155 40552 97164
rect 40500 97121 40509 97155
rect 40509 97121 40543 97155
rect 40543 97121 40552 97155
rect 40500 97112 40552 97121
rect 43076 97155 43128 97164
rect 43076 97121 43085 97155
rect 43085 97121 43119 97155
rect 43119 97121 43128 97155
rect 43076 97112 43128 97121
rect 44732 97180 44784 97232
rect 47308 97180 47360 97232
rect 48136 97180 48188 97232
rect 50804 97180 50856 97232
rect 53380 97180 53432 97232
rect 55956 97180 56008 97232
rect 57704 97180 57756 97232
rect 58624 97180 58676 97232
rect 60372 97180 60424 97232
rect 61200 97180 61252 97232
rect 63868 97180 63920 97232
rect 65524 97180 65576 97232
rect 66444 97180 66496 97232
rect 68560 97223 68612 97232
rect 68560 97189 68569 97223
rect 68569 97189 68603 97223
rect 68603 97189 68612 97223
rect 68560 97180 68612 97189
rect 69020 97180 69072 97232
rect 69940 97180 69992 97232
rect 74264 97180 74316 97232
rect 76012 97180 76064 97232
rect 76840 97180 76892 97232
rect 79508 97180 79560 97232
rect 82084 97180 82136 97232
rect 84660 97223 84712 97232
rect 84660 97189 84669 97223
rect 84669 97189 84703 97223
rect 84703 97189 84712 97223
rect 84660 97180 84712 97189
rect 87328 97223 87380 97232
rect 87328 97189 87337 97223
rect 87337 97189 87371 97223
rect 87371 97189 87380 97223
rect 87328 97180 87380 97189
rect 89904 97223 89956 97232
rect 89904 97189 89913 97223
rect 89913 97189 89947 97223
rect 89947 97189 89956 97223
rect 89904 97180 89956 97189
rect 42064 97044 42116 97096
rect 45468 97112 45520 97164
rect 48320 97155 48372 97164
rect 48320 97121 48329 97155
rect 48329 97121 48363 97155
rect 48363 97121 48372 97155
rect 48320 97112 48372 97121
rect 49884 97155 49936 97164
rect 49884 97121 49893 97155
rect 49893 97121 49927 97155
rect 49927 97121 49936 97155
rect 49884 97112 49936 97121
rect 50896 97155 50948 97164
rect 50896 97121 50905 97155
rect 50905 97121 50939 97155
rect 50939 97121 50948 97155
rect 50896 97112 50948 97121
rect 52552 97155 52604 97164
rect 52552 97121 52561 97155
rect 52561 97121 52595 97155
rect 52595 97121 52604 97155
rect 52552 97112 52604 97121
rect 53472 97155 53524 97164
rect 53472 97121 53481 97155
rect 53481 97121 53515 97155
rect 53515 97121 53524 97155
rect 53472 97112 53524 97121
rect 55128 97155 55180 97164
rect 55128 97121 55137 97155
rect 55137 97121 55171 97155
rect 55171 97121 55180 97155
rect 55128 97112 55180 97121
rect 43444 97044 43496 97096
rect 4896 96976 4948 97028
rect 47584 97019 47636 97028
rect 1584 96951 1636 96960
rect 1584 96917 1593 96951
rect 1593 96917 1627 96951
rect 1627 96917 1636 96951
rect 1584 96908 1636 96917
rect 3056 96951 3108 96960
rect 3056 96917 3065 96951
rect 3065 96917 3099 96951
rect 3099 96917 3108 96951
rect 3056 96908 3108 96917
rect 11060 96908 11112 96960
rect 16212 96951 16264 96960
rect 16212 96917 16221 96951
rect 16221 96917 16255 96951
rect 16255 96917 16264 96951
rect 16212 96908 16264 96917
rect 18788 96951 18840 96960
rect 18788 96917 18797 96951
rect 18797 96917 18831 96951
rect 18831 96917 18840 96951
rect 18788 96908 18840 96917
rect 23572 96908 23624 96960
rect 24492 96908 24544 96960
rect 26608 96951 26660 96960
rect 26608 96917 26617 96951
rect 26617 96917 26651 96951
rect 26651 96917 26660 96951
rect 26608 96908 26660 96917
rect 29184 96951 29236 96960
rect 29184 96917 29193 96951
rect 29193 96917 29227 96951
rect 29227 96917 29236 96951
rect 29184 96908 29236 96917
rect 31852 96951 31904 96960
rect 31852 96917 31861 96951
rect 31861 96917 31895 96951
rect 31895 96917 31904 96951
rect 31852 96908 31904 96917
rect 37096 96908 37148 96960
rect 39672 96951 39724 96960
rect 39672 96917 39681 96951
rect 39681 96917 39715 96951
rect 39715 96917 39724 96951
rect 39672 96908 39724 96917
rect 42248 96951 42300 96960
rect 42248 96917 42257 96951
rect 42257 96917 42291 96951
rect 42291 96917 42300 96951
rect 42248 96908 42300 96917
rect 44916 96951 44968 96960
rect 44916 96917 44925 96951
rect 44925 96917 44959 96951
rect 44959 96917 44968 96951
rect 44916 96908 44968 96917
rect 45560 96908 45612 96960
rect 47584 96985 47593 97019
rect 47593 96985 47627 97019
rect 47627 96985 47636 97019
rect 47584 96976 47636 96985
rect 56416 97112 56468 97164
rect 61384 97155 61436 97164
rect 61384 97121 61393 97155
rect 61393 97121 61427 97155
rect 61427 97121 61436 97155
rect 61384 97112 61436 97121
rect 62948 97155 63000 97164
rect 62948 97121 62957 97155
rect 62957 97121 62991 97155
rect 62991 97121 63000 97155
rect 62948 97112 63000 97121
rect 63960 97155 64012 97164
rect 63960 97121 63969 97155
rect 63969 97121 64003 97155
rect 64003 97121 64012 97155
rect 63960 97112 64012 97121
rect 66536 97155 66588 97164
rect 66536 97121 66545 97155
rect 66545 97121 66579 97155
rect 66579 97121 66588 97155
rect 66536 97112 66588 97121
rect 68192 97112 68244 97164
rect 69296 97155 69348 97164
rect 69296 97121 69305 97155
rect 69305 97121 69339 97155
rect 69339 97121 69348 97155
rect 69296 97112 69348 97121
rect 71044 97155 71096 97164
rect 71044 97121 71053 97155
rect 71053 97121 71087 97155
rect 71087 97121 71096 97155
rect 71044 97112 71096 97121
rect 71872 97112 71924 97164
rect 72332 97112 72384 97164
rect 73344 97112 73396 97164
rect 74448 97155 74500 97164
rect 74448 97121 74457 97155
rect 74457 97121 74491 97155
rect 74491 97121 74500 97155
rect 74448 97112 74500 97121
rect 75184 97155 75236 97164
rect 75184 97121 75193 97155
rect 75193 97121 75227 97155
rect 75227 97121 75236 97155
rect 75184 97112 75236 97121
rect 77300 97155 77352 97164
rect 77300 97121 77309 97155
rect 77309 97121 77343 97155
rect 77343 97121 77352 97155
rect 77300 97112 77352 97121
rect 78680 97112 78732 97164
rect 79968 97155 80020 97164
rect 79968 97121 79977 97155
rect 79977 97121 80011 97155
rect 80011 97121 80020 97155
rect 79968 97112 80020 97121
rect 82176 97155 82228 97164
rect 82176 97121 82185 97155
rect 82185 97121 82219 97155
rect 82219 97121 82228 97155
rect 82176 97112 82228 97121
rect 82912 97155 82964 97164
rect 82912 97121 82921 97155
rect 82921 97121 82955 97155
rect 82955 97121 82964 97155
rect 82912 97112 82964 97121
rect 85028 97112 85080 97164
rect 85488 97155 85540 97164
rect 85488 97121 85497 97155
rect 85497 97121 85531 97155
rect 85531 97121 85540 97155
rect 85488 97112 85540 97121
rect 87512 97155 87564 97164
rect 87512 97121 87521 97155
rect 87521 97121 87555 97155
rect 87555 97121 87564 97155
rect 87512 97112 87564 97121
rect 88156 97155 88208 97164
rect 88156 97121 88165 97155
rect 88165 97121 88199 97155
rect 88199 97121 88208 97155
rect 88156 97112 88208 97121
rect 89720 97112 89772 97164
rect 90456 97257 90465 97291
rect 90465 97257 90499 97291
rect 90499 97257 90508 97291
rect 90456 97248 90508 97257
rect 92480 97223 92532 97232
rect 92480 97189 92489 97223
rect 92489 97189 92523 97223
rect 92523 97189 92532 97223
rect 92480 97180 92532 97189
rect 95148 97223 95200 97232
rect 95148 97189 95157 97223
rect 95157 97189 95191 97223
rect 95191 97189 95200 97223
rect 95148 97180 95200 97189
rect 97724 97223 97776 97232
rect 97724 97189 97733 97223
rect 97733 97189 97767 97223
rect 97767 97189 97776 97223
rect 97724 97180 97776 97189
rect 69664 97044 69716 97096
rect 79140 97087 79192 97096
rect 79140 97053 79149 97087
rect 79149 97053 79183 97087
rect 79183 97053 79192 97087
rect 79140 97044 79192 97053
rect 84108 97044 84160 97096
rect 57980 97019 58032 97028
rect 57980 96985 57989 97019
rect 57989 96985 58023 97019
rect 58023 96985 58032 97019
rect 57980 96976 58032 96985
rect 65984 96976 66036 97028
rect 80704 96976 80756 97028
rect 88340 97019 88392 97028
rect 88340 96985 88349 97019
rect 88349 96985 88383 97019
rect 88383 96985 88392 97019
rect 88340 96976 88392 96985
rect 90640 97019 90692 97028
rect 90640 96985 90649 97019
rect 90649 96985 90683 97019
rect 90683 96985 90692 97019
rect 90640 96976 90692 96985
rect 52736 96951 52788 96960
rect 52736 96917 52745 96951
rect 52745 96917 52779 96951
rect 52779 96917 52788 96951
rect 52736 96908 52788 96917
rect 60740 96951 60792 96960
rect 60740 96917 60749 96951
rect 60749 96917 60783 96951
rect 60783 96917 60792 96951
rect 60740 96908 60792 96917
rect 63132 96951 63184 96960
rect 63132 96917 63141 96951
rect 63141 96917 63175 96951
rect 63175 96917 63184 96951
rect 63132 96908 63184 96917
rect 71136 96951 71188 96960
rect 71136 96917 71145 96951
rect 71145 96917 71179 96951
rect 71179 96917 71188 96951
rect 71136 96908 71188 96917
rect 71780 96908 71832 96960
rect 72516 96908 72568 96960
rect 76380 96908 76432 96960
rect 82820 96908 82872 96960
rect 85028 96951 85080 96960
rect 85028 96917 85037 96951
rect 85037 96917 85071 96951
rect 85071 96917 85080 96951
rect 85028 96908 85080 96917
rect 87512 96908 87564 96960
rect 89720 96951 89772 96960
rect 89720 96917 89729 96951
rect 89729 96917 89763 96951
rect 89763 96917 89772 96951
rect 92296 96951 92348 96960
rect 89720 96908 89772 96917
rect 92296 96917 92305 96951
rect 92305 96917 92339 96951
rect 92339 96917 92348 96951
rect 93308 97112 93360 97164
rect 92756 96976 92808 97028
rect 92296 96908 92348 96917
rect 94964 96951 95016 96960
rect 94964 96917 94973 96951
rect 94973 96917 95007 96951
rect 95007 96917 95016 96951
rect 95884 97019 95936 97028
rect 95884 96985 95893 97019
rect 95893 96985 95927 97019
rect 95927 96985 95936 97019
rect 95884 96976 95936 96985
rect 94964 96908 95016 96917
rect 97540 96951 97592 96960
rect 97540 96917 97549 96951
rect 97549 96917 97583 96951
rect 97583 96917 97592 96951
rect 97540 96908 97592 96917
rect 4246 96806 4298 96858
rect 4310 96806 4362 96858
rect 4374 96806 4426 96858
rect 4438 96806 4490 96858
rect 34966 96806 35018 96858
rect 35030 96806 35082 96858
rect 35094 96806 35146 96858
rect 35158 96806 35210 96858
rect 65686 96806 65738 96858
rect 65750 96806 65802 96858
rect 65814 96806 65866 96858
rect 65878 96806 65930 96858
rect 96406 96806 96458 96858
rect 96470 96806 96522 96858
rect 96534 96806 96586 96858
rect 96598 96806 96650 96858
rect 16304 96747 16356 96756
rect 16304 96713 16313 96747
rect 16313 96713 16347 96747
rect 16347 96713 16356 96747
rect 16304 96704 16356 96713
rect 14464 96636 14516 96688
rect 21364 96704 21416 96756
rect 34612 96704 34664 96756
rect 79140 96704 79192 96756
rect 40684 96636 40736 96688
rect 43444 96636 43496 96688
rect 2044 96568 2096 96620
rect 4712 96568 4764 96620
rect 7288 96611 7340 96620
rect 7288 96577 7297 96611
rect 7297 96577 7331 96611
rect 7331 96577 7340 96611
rect 7288 96568 7340 96577
rect 9864 96568 9916 96620
rect 12532 96568 12584 96620
rect 15108 96568 15160 96620
rect 17776 96568 17828 96620
rect 22928 96568 22980 96620
rect 25596 96568 25648 96620
rect 33416 96568 33468 96620
rect 35992 96568 36044 96620
rect 38568 96568 38620 96620
rect 41236 96568 41288 96620
rect 43812 96568 43864 96620
rect 49056 96568 49108 96620
rect 51632 96568 51684 96620
rect 54300 96568 54352 96620
rect 56876 96568 56928 96620
rect 59452 96568 59504 96620
rect 62120 96568 62172 96620
rect 64696 96568 64748 96620
rect 67272 96568 67324 96620
rect 71136 96568 71188 96620
rect 75092 96568 75144 96620
rect 80336 96568 80388 96620
rect 84108 96568 84160 96620
rect 85580 96568 85632 96620
rect 90640 96568 90692 96620
rect 90824 96568 90876 96620
rect 93400 96611 93452 96620
rect 20444 96500 20496 96552
rect 23572 96500 23624 96552
rect 23848 96543 23900 96552
rect 23848 96509 23857 96543
rect 23857 96509 23891 96543
rect 23891 96509 23900 96543
rect 23848 96500 23900 96509
rect 38752 96500 38804 96552
rect 46112 96500 46164 96552
rect 46480 96500 46532 96552
rect 46756 96543 46808 96552
rect 46756 96509 46765 96543
rect 46765 96509 46799 96543
rect 46799 96509 46808 96543
rect 46756 96500 46808 96509
rect 47032 96543 47084 96552
rect 47032 96509 47041 96543
rect 47041 96509 47075 96543
rect 47075 96509 47084 96543
rect 47032 96500 47084 96509
rect 47216 96543 47268 96552
rect 47216 96509 47225 96543
rect 47225 96509 47259 96543
rect 47259 96509 47268 96543
rect 47216 96500 47268 96509
rect 70768 96543 70820 96552
rect 70768 96509 70777 96543
rect 70777 96509 70811 96543
rect 70811 96509 70820 96543
rect 70768 96500 70820 96509
rect 81348 96500 81400 96552
rect 83832 96543 83884 96552
rect 83832 96509 83841 96543
rect 83841 96509 83875 96543
rect 83875 96509 83884 96543
rect 83832 96500 83884 96509
rect 86408 96543 86460 96552
rect 86408 96509 86417 96543
rect 86417 96509 86451 96543
rect 86451 96509 86460 96543
rect 86408 96500 86460 96509
rect 89076 96543 89128 96552
rect 89076 96509 89085 96543
rect 89085 96509 89119 96543
rect 89119 96509 89128 96543
rect 89076 96500 89128 96509
rect 91652 96543 91704 96552
rect 91652 96509 91661 96543
rect 91661 96509 91695 96543
rect 91695 96509 91704 96543
rect 91652 96500 91704 96509
rect 93400 96577 93409 96611
rect 93409 96577 93443 96611
rect 93443 96577 93452 96611
rect 93400 96568 93452 96577
rect 95884 96568 95936 96620
rect 95976 96568 96028 96620
rect 98644 96568 98696 96620
rect 94228 96543 94280 96552
rect 94228 96509 94237 96543
rect 94237 96509 94271 96543
rect 94271 96509 94280 96543
rect 94228 96500 94280 96509
rect 99472 96500 99524 96552
rect 2136 96475 2188 96484
rect 2136 96441 2145 96475
rect 2145 96441 2179 96475
rect 2179 96441 2188 96475
rect 2136 96432 2188 96441
rect 4804 96475 4856 96484
rect 4804 96441 4813 96475
rect 4813 96441 4847 96475
rect 4847 96441 4856 96475
rect 4804 96432 4856 96441
rect 9956 96475 10008 96484
rect 7104 96407 7156 96416
rect 7104 96373 7113 96407
rect 7113 96373 7147 96407
rect 7147 96373 7156 96407
rect 9956 96441 9965 96475
rect 9965 96441 9999 96475
rect 9999 96441 10008 96475
rect 9956 96432 10008 96441
rect 12624 96475 12676 96484
rect 12624 96441 12633 96475
rect 12633 96441 12667 96475
rect 12667 96441 12676 96475
rect 12624 96432 12676 96441
rect 17868 96475 17920 96484
rect 17868 96441 17877 96475
rect 17877 96441 17911 96475
rect 17911 96441 17920 96475
rect 17868 96432 17920 96441
rect 23020 96475 23072 96484
rect 23020 96441 23029 96475
rect 23029 96441 23063 96475
rect 23063 96441 23072 96475
rect 23020 96432 23072 96441
rect 25688 96475 25740 96484
rect 25688 96441 25697 96475
rect 25697 96441 25731 96475
rect 25731 96441 25740 96475
rect 25688 96432 25740 96441
rect 30380 96432 30432 96484
rect 36084 96475 36136 96484
rect 36084 96441 36093 96475
rect 36093 96441 36127 96475
rect 36127 96441 36136 96475
rect 36084 96432 36136 96441
rect 38660 96475 38712 96484
rect 38660 96441 38669 96475
rect 38669 96441 38703 96475
rect 38703 96441 38712 96475
rect 38660 96432 38712 96441
rect 41328 96475 41380 96484
rect 41328 96441 41337 96475
rect 41337 96441 41371 96475
rect 41371 96441 41380 96475
rect 41328 96432 41380 96441
rect 49148 96475 49200 96484
rect 49148 96441 49157 96475
rect 49157 96441 49191 96475
rect 49191 96441 49200 96475
rect 49148 96432 49200 96441
rect 51724 96475 51776 96484
rect 51724 96441 51733 96475
rect 51733 96441 51767 96475
rect 51767 96441 51776 96475
rect 51724 96432 51776 96441
rect 54392 96475 54444 96484
rect 54392 96441 54401 96475
rect 54401 96441 54435 96475
rect 54435 96441 54444 96475
rect 54392 96432 54444 96441
rect 56968 96475 57020 96484
rect 56968 96441 56977 96475
rect 56977 96441 57011 96475
rect 57011 96441 57020 96475
rect 56968 96432 57020 96441
rect 59544 96475 59596 96484
rect 59544 96441 59553 96475
rect 59553 96441 59587 96475
rect 59587 96441 59596 96475
rect 59544 96432 59596 96441
rect 62212 96475 62264 96484
rect 62212 96441 62221 96475
rect 62221 96441 62255 96475
rect 62255 96441 62264 96475
rect 62212 96432 62264 96441
rect 64788 96475 64840 96484
rect 64788 96441 64797 96475
rect 64797 96441 64831 96475
rect 64831 96441 64840 96475
rect 64788 96432 64840 96441
rect 74540 96432 74592 96484
rect 77760 96432 77812 96484
rect 82820 96432 82872 96484
rect 88248 96432 88300 96484
rect 92756 96432 92808 96484
rect 96068 96475 96120 96484
rect 7104 96364 7156 96373
rect 20444 96364 20496 96416
rect 24032 96407 24084 96416
rect 24032 96373 24041 96407
rect 24041 96373 24075 96407
rect 24075 96373 24084 96407
rect 24032 96364 24084 96373
rect 47492 96407 47544 96416
rect 47492 96373 47501 96407
rect 47501 96373 47535 96407
rect 47535 96373 47544 96407
rect 47492 96364 47544 96373
rect 70860 96364 70912 96416
rect 81440 96407 81492 96416
rect 81440 96373 81449 96407
rect 81449 96373 81483 96407
rect 81483 96373 81492 96407
rect 81440 96364 81492 96373
rect 83004 96364 83056 96416
rect 88340 96364 88392 96416
rect 93216 96407 93268 96416
rect 93216 96373 93225 96407
rect 93225 96373 93259 96407
rect 93259 96373 93268 96407
rect 96068 96441 96077 96475
rect 96077 96441 96111 96475
rect 96111 96441 96120 96475
rect 96068 96432 96120 96441
rect 97908 96475 97960 96484
rect 93216 96364 93268 96373
rect 95884 96364 95936 96416
rect 97908 96441 97917 96475
rect 97917 96441 97951 96475
rect 97951 96441 97960 96475
rect 97908 96432 97960 96441
rect 19606 96262 19658 96314
rect 19670 96262 19722 96314
rect 19734 96262 19786 96314
rect 19798 96262 19850 96314
rect 50326 96262 50378 96314
rect 50390 96262 50442 96314
rect 50454 96262 50506 96314
rect 50518 96262 50570 96314
rect 81046 96262 81098 96314
rect 81110 96262 81162 96314
rect 81174 96262 81226 96314
rect 81238 96262 81290 96314
rect 2136 96160 2188 96212
rect 14556 96160 14608 96212
rect 46388 96160 46440 96212
rect 49148 96160 49200 96212
rect 60096 96160 60148 96212
rect 30288 96024 30340 96076
rect 46848 96024 46900 96076
rect 57428 96067 57480 96076
rect 57428 96033 57437 96067
rect 57437 96033 57471 96067
rect 57471 96033 57480 96067
rect 57428 96024 57480 96033
rect 57796 96067 57848 96076
rect 57796 96033 57805 96067
rect 57805 96033 57839 96067
rect 57839 96033 57848 96067
rect 57796 96024 57848 96033
rect 58164 96067 58216 96076
rect 58164 96033 58173 96067
rect 58173 96033 58207 96067
rect 58207 96033 58216 96067
rect 58164 96024 58216 96033
rect 26884 95956 26936 96008
rect 30380 95956 30432 96008
rect 57612 95999 57664 96008
rect 57612 95965 57621 95999
rect 57621 95965 57655 95999
rect 57655 95965 57664 95999
rect 57612 95956 57664 95965
rect 30656 95888 30708 95940
rect 56508 95888 56560 95940
rect 58532 95931 58584 95940
rect 58532 95897 58541 95931
rect 58541 95897 58575 95931
rect 58575 95897 58584 95931
rect 58532 95888 58584 95897
rect 83464 96024 83516 96076
rect 96896 96067 96948 96076
rect 96896 96033 96905 96067
rect 96905 96033 96939 96067
rect 96939 96033 96948 96067
rect 96896 96024 96948 96033
rect 83832 95999 83884 96008
rect 83832 95965 83841 95999
rect 83841 95965 83875 95999
rect 83875 95965 83884 95999
rect 83832 95956 83884 95965
rect 83924 95888 83976 95940
rect 4246 95718 4298 95770
rect 4310 95718 4362 95770
rect 4374 95718 4426 95770
rect 4438 95718 4490 95770
rect 34966 95718 35018 95770
rect 35030 95718 35082 95770
rect 35094 95718 35146 95770
rect 35158 95718 35210 95770
rect 65686 95718 65738 95770
rect 65750 95718 65802 95770
rect 65814 95718 65866 95770
rect 65878 95718 65930 95770
rect 96406 95718 96458 95770
rect 96470 95718 96522 95770
rect 96534 95718 96586 95770
rect 96598 95718 96650 95770
rect 46756 95616 46808 95668
rect 88984 95616 89036 95668
rect 53840 95591 53892 95600
rect 53840 95557 53849 95591
rect 53849 95557 53883 95591
rect 53883 95557 53892 95591
rect 53840 95548 53892 95557
rect 10876 95387 10928 95396
rect 10876 95353 10885 95387
rect 10885 95353 10919 95387
rect 10919 95353 10928 95387
rect 10876 95344 10928 95353
rect 35348 95455 35400 95464
rect 35348 95421 35357 95455
rect 35357 95421 35391 95455
rect 35391 95421 35400 95455
rect 35348 95412 35400 95421
rect 57980 95480 58032 95532
rect 31392 95344 31444 95396
rect 66904 95412 66956 95464
rect 61660 95344 61712 95396
rect 96160 95276 96212 95328
rect 19606 95174 19658 95226
rect 19670 95174 19722 95226
rect 19734 95174 19786 95226
rect 19798 95174 19850 95226
rect 50326 95174 50378 95226
rect 50390 95174 50442 95226
rect 50454 95174 50506 95226
rect 50518 95174 50570 95226
rect 81046 95174 81098 95226
rect 81110 95174 81162 95226
rect 81174 95174 81226 95226
rect 81238 95174 81290 95226
rect 42248 95004 42300 95056
rect 2596 94936 2648 94988
rect 5448 94936 5500 94988
rect 14924 94979 14976 94988
rect 14924 94945 14933 94979
rect 14933 94945 14967 94979
rect 14967 94945 14976 94979
rect 14924 94936 14976 94945
rect 15384 94979 15436 94988
rect 15384 94945 15387 94979
rect 15387 94945 15436 94979
rect 9864 94868 9916 94920
rect 15384 94936 15436 94945
rect 38752 94868 38804 94920
rect 2596 94800 2648 94852
rect 53932 94843 53984 94852
rect 53932 94809 53941 94843
rect 53941 94809 53975 94843
rect 53975 94809 53984 94843
rect 53932 94800 53984 94809
rect 55404 94936 55456 94988
rect 56416 94936 56468 94988
rect 54576 94911 54628 94920
rect 54576 94877 54585 94911
rect 54585 94877 54619 94911
rect 54619 94877 54628 94911
rect 54576 94868 54628 94877
rect 66076 94800 66128 94852
rect 2044 94775 2096 94784
rect 2044 94741 2053 94775
rect 2053 94741 2087 94775
rect 2087 94741 2096 94775
rect 2044 94732 2096 94741
rect 5172 94775 5224 94784
rect 5172 94741 5181 94775
rect 5181 94741 5215 94775
rect 5215 94741 5224 94775
rect 5172 94732 5224 94741
rect 15476 94775 15528 94784
rect 15476 94741 15485 94775
rect 15485 94741 15519 94775
rect 15519 94741 15528 94775
rect 15476 94732 15528 94741
rect 4246 94630 4298 94682
rect 4310 94630 4362 94682
rect 4374 94630 4426 94682
rect 4438 94630 4490 94682
rect 34966 94630 35018 94682
rect 35030 94630 35082 94682
rect 35094 94630 35146 94682
rect 35158 94630 35210 94682
rect 65686 94630 65738 94682
rect 65750 94630 65802 94682
rect 65814 94630 65866 94682
rect 65878 94630 65930 94682
rect 96406 94630 96458 94682
rect 96470 94630 96522 94682
rect 96534 94630 96586 94682
rect 96598 94630 96650 94682
rect 2596 94528 2648 94580
rect 25872 94324 25924 94376
rect 41880 94367 41932 94376
rect 41880 94333 41889 94367
rect 41889 94333 41923 94367
rect 41923 94333 41932 94367
rect 41880 94324 41932 94333
rect 66168 94392 66220 94444
rect 63224 94367 63276 94376
rect 63224 94333 63233 94367
rect 63233 94333 63267 94367
rect 63267 94333 63276 94367
rect 63224 94324 63276 94333
rect 63408 94299 63460 94308
rect 63408 94265 63417 94299
rect 63417 94265 63451 94299
rect 63451 94265 63460 94299
rect 63408 94256 63460 94265
rect 25504 94188 25556 94240
rect 63040 94231 63092 94240
rect 63040 94197 63049 94231
rect 63049 94197 63083 94231
rect 63083 94197 63092 94231
rect 63040 94188 63092 94197
rect 71872 94188 71924 94240
rect 72424 94188 72476 94240
rect 19606 94086 19658 94138
rect 19670 94086 19722 94138
rect 19734 94086 19786 94138
rect 19798 94086 19850 94138
rect 50326 94086 50378 94138
rect 50390 94086 50442 94138
rect 50454 94086 50506 94138
rect 50518 94086 50570 94138
rect 81046 94086 81098 94138
rect 81110 94086 81162 94138
rect 81174 94086 81226 94138
rect 81238 94086 81290 94138
rect 83832 93984 83884 94036
rect 49884 93916 49936 93968
rect 95608 93916 95660 93968
rect 44824 93848 44876 93900
rect 45468 93848 45520 93900
rect 95976 93891 96028 93900
rect 95976 93857 95985 93891
rect 95985 93857 96019 93891
rect 96019 93857 96028 93891
rect 95976 93848 96028 93857
rect 10692 93780 10744 93832
rect 69296 93780 69348 93832
rect 40500 93712 40552 93764
rect 83464 93712 83516 93764
rect 95608 93644 95660 93696
rect 4246 93542 4298 93594
rect 4310 93542 4362 93594
rect 4374 93542 4426 93594
rect 4438 93542 4490 93594
rect 34966 93542 35018 93594
rect 35030 93542 35082 93594
rect 35094 93542 35146 93594
rect 35158 93542 35210 93594
rect 65686 93542 65738 93594
rect 65750 93542 65802 93594
rect 65814 93542 65866 93594
rect 65878 93542 65930 93594
rect 96406 93542 96458 93594
rect 96470 93542 96522 93594
rect 96534 93542 96586 93594
rect 96598 93542 96650 93594
rect 9864 93304 9916 93356
rect 10692 93304 10744 93356
rect 58072 93236 58124 93288
rect 74448 93236 74500 93288
rect 34520 93168 34572 93220
rect 35348 93168 35400 93220
rect 59544 93168 59596 93220
rect 11704 93100 11756 93152
rect 40500 93100 40552 93152
rect 69296 93100 69348 93152
rect 85856 93100 85908 93152
rect 19606 92998 19658 93050
rect 19670 92998 19722 93050
rect 19734 92998 19786 93050
rect 19798 92998 19850 93050
rect 50326 92998 50378 93050
rect 50390 92998 50442 93050
rect 50454 92998 50506 93050
rect 50518 92998 50570 93050
rect 81046 92998 81098 93050
rect 81110 92998 81162 93050
rect 81174 92998 81226 93050
rect 81238 92998 81290 93050
rect 59544 92556 59596 92608
rect 60556 92556 60608 92608
rect 4246 92454 4298 92506
rect 4310 92454 4362 92506
rect 4374 92454 4426 92506
rect 4438 92454 4490 92506
rect 34966 92454 35018 92506
rect 35030 92454 35082 92506
rect 35094 92454 35146 92506
rect 35158 92454 35210 92506
rect 65686 92454 65738 92506
rect 65750 92454 65802 92506
rect 65814 92454 65866 92506
rect 65878 92454 65930 92506
rect 96406 92454 96458 92506
rect 96470 92454 96522 92506
rect 96534 92454 96586 92506
rect 96598 92454 96650 92506
rect 68928 92284 68980 92336
rect 93768 92327 93820 92336
rect 93768 92293 93777 92327
rect 93777 92293 93811 92327
rect 93811 92293 93820 92327
rect 93768 92284 93820 92293
rect 92664 92259 92716 92268
rect 92664 92225 92673 92259
rect 92673 92225 92707 92259
rect 92707 92225 92716 92259
rect 92664 92216 92716 92225
rect 93860 92259 93912 92268
rect 93860 92225 93869 92259
rect 93869 92225 93903 92259
rect 93903 92225 93912 92259
rect 93860 92216 93912 92225
rect 36360 92191 36412 92200
rect 36360 92157 36369 92191
rect 36369 92157 36403 92191
rect 36403 92157 36412 92191
rect 36360 92148 36412 92157
rect 92480 92191 92532 92200
rect 92480 92157 92486 92191
rect 92486 92157 92532 92191
rect 92480 92148 92532 92157
rect 93676 92191 93728 92200
rect 93676 92157 93682 92191
rect 93682 92157 93728 92191
rect 93676 92148 93728 92157
rect 23480 92123 23532 92132
rect 23480 92089 23489 92123
rect 23489 92089 23523 92123
rect 23523 92089 23532 92123
rect 23480 92080 23532 92089
rect 23664 92123 23716 92132
rect 23664 92089 23673 92123
rect 23673 92089 23707 92123
rect 23707 92089 23716 92123
rect 23664 92080 23716 92089
rect 35440 92080 35492 92132
rect 92204 92080 92256 92132
rect 93492 92123 93544 92132
rect 93492 92089 93501 92123
rect 93501 92089 93535 92123
rect 93535 92089 93544 92123
rect 93492 92080 93544 92089
rect 84292 92012 84344 92064
rect 94136 92055 94188 92064
rect 94136 92021 94145 92055
rect 94145 92021 94179 92055
rect 94179 92021 94188 92055
rect 94136 92012 94188 92021
rect 19606 91910 19658 91962
rect 19670 91910 19722 91962
rect 19734 91910 19786 91962
rect 19798 91910 19850 91962
rect 50326 91910 50378 91962
rect 50390 91910 50442 91962
rect 50454 91910 50506 91962
rect 50518 91910 50570 91962
rect 81046 91910 81098 91962
rect 81110 91910 81162 91962
rect 81174 91910 81226 91962
rect 81238 91910 81290 91962
rect 11796 91740 11848 91792
rect 46480 91740 46532 91792
rect 49056 91808 49108 91860
rect 65248 91808 65300 91860
rect 27068 91604 27120 91656
rect 48964 91740 49016 91792
rect 68468 91672 68520 91724
rect 68928 91672 68980 91724
rect 73620 91715 73672 91724
rect 73620 91681 73629 91715
rect 73629 91681 73663 91715
rect 73663 91681 73672 91715
rect 73620 91672 73672 91681
rect 74172 91715 74224 91724
rect 14740 91468 14792 91520
rect 47952 91511 48004 91520
rect 47952 91477 47961 91511
rect 47961 91477 47995 91511
rect 47995 91477 48004 91511
rect 47952 91468 48004 91477
rect 61568 91536 61620 91588
rect 74172 91681 74181 91715
rect 74181 91681 74215 91715
rect 74215 91681 74224 91715
rect 74172 91672 74224 91681
rect 73988 91647 74040 91656
rect 73988 91613 73997 91647
rect 73997 91613 74031 91647
rect 74031 91613 74040 91647
rect 73988 91604 74040 91613
rect 74356 91579 74408 91588
rect 74356 91545 74365 91579
rect 74365 91545 74399 91579
rect 74399 91545 74408 91579
rect 74356 91536 74408 91545
rect 4246 91366 4298 91418
rect 4310 91366 4362 91418
rect 4374 91366 4426 91418
rect 4438 91366 4490 91418
rect 34966 91366 35018 91418
rect 35030 91366 35082 91418
rect 35094 91366 35146 91418
rect 35158 91366 35210 91418
rect 65686 91366 65738 91418
rect 65750 91366 65802 91418
rect 65814 91366 65866 91418
rect 65878 91366 65930 91418
rect 96406 91366 96458 91418
rect 96470 91366 96522 91418
rect 96534 91366 96586 91418
rect 96598 91366 96650 91418
rect 68560 91264 68612 91316
rect 73988 91264 74040 91316
rect 52460 91128 52512 91180
rect 55036 91060 55088 91112
rect 61476 91060 61528 91112
rect 19606 90822 19658 90874
rect 19670 90822 19722 90874
rect 19734 90822 19786 90874
rect 19798 90822 19850 90874
rect 50326 90822 50378 90874
rect 50390 90822 50442 90874
rect 50454 90822 50506 90874
rect 50518 90822 50570 90874
rect 81046 90822 81098 90874
rect 81110 90822 81162 90874
rect 81174 90822 81226 90874
rect 81238 90822 81290 90874
rect 8300 90584 8352 90636
rect 69848 90627 69900 90636
rect 69848 90593 69857 90627
rect 69857 90593 69891 90627
rect 69891 90593 69900 90627
rect 69848 90584 69900 90593
rect 70308 90559 70360 90568
rect 70308 90525 70317 90559
rect 70317 90525 70351 90559
rect 70351 90525 70360 90559
rect 70308 90516 70360 90525
rect 9680 90423 9732 90432
rect 9680 90389 9689 90423
rect 9689 90389 9723 90423
rect 9723 90389 9732 90423
rect 9680 90380 9732 90389
rect 39396 90380 39448 90432
rect 74356 90380 74408 90432
rect 91744 90380 91796 90432
rect 4246 90278 4298 90330
rect 4310 90278 4362 90330
rect 4374 90278 4426 90330
rect 4438 90278 4490 90330
rect 34966 90278 35018 90330
rect 35030 90278 35082 90330
rect 35094 90278 35146 90330
rect 35158 90278 35210 90330
rect 65686 90278 65738 90330
rect 65750 90278 65802 90330
rect 65814 90278 65866 90330
rect 65878 90278 65930 90330
rect 96406 90278 96458 90330
rect 96470 90278 96522 90330
rect 96534 90278 96586 90330
rect 96598 90278 96650 90330
rect 41052 90176 41104 90228
rect 29276 90015 29328 90024
rect 29276 89981 29285 90015
rect 29285 89981 29319 90015
rect 29319 89981 29328 90015
rect 29276 89972 29328 89981
rect 29460 90015 29512 90024
rect 29460 89981 29468 90015
rect 29468 89981 29502 90015
rect 29502 89981 29512 90015
rect 29460 89972 29512 89981
rect 28264 89904 28316 89956
rect 30288 89972 30340 90024
rect 30748 90015 30800 90024
rect 4068 89836 4120 89888
rect 30748 89981 30757 90015
rect 30757 89981 30791 90015
rect 30791 89981 30800 90015
rect 30748 89972 30800 89981
rect 44456 89972 44508 90024
rect 49976 90108 50028 90160
rect 63040 89972 63092 90024
rect 75276 90015 75328 90024
rect 75276 89981 75280 90015
rect 75280 89981 75314 90015
rect 75314 89981 75328 90015
rect 75276 89972 75328 89981
rect 75828 89972 75880 90024
rect 44180 89947 44232 89956
rect 44180 89913 44214 89947
rect 44214 89913 44232 89947
rect 44180 89904 44232 89913
rect 46848 89904 46900 89956
rect 76196 89947 76248 89956
rect 31944 89836 31996 89888
rect 44916 89836 44968 89888
rect 76196 89913 76205 89947
rect 76205 89913 76239 89947
rect 76239 89913 76248 89947
rect 76196 89904 76248 89913
rect 75736 89879 75788 89888
rect 75736 89845 75745 89879
rect 75745 89845 75779 89879
rect 75779 89845 75788 89879
rect 75736 89836 75788 89845
rect 76288 89879 76340 89888
rect 76288 89845 76297 89879
rect 76297 89845 76331 89879
rect 76331 89845 76340 89879
rect 76288 89836 76340 89845
rect 19606 89734 19658 89786
rect 19670 89734 19722 89786
rect 19734 89734 19786 89786
rect 19798 89734 19850 89786
rect 50326 89734 50378 89786
rect 50390 89734 50442 89786
rect 50454 89734 50506 89786
rect 50518 89734 50570 89786
rect 81046 89734 81098 89786
rect 81110 89734 81162 89786
rect 81174 89734 81226 89786
rect 81238 89734 81290 89786
rect 48964 89564 49016 89616
rect 31116 89496 31168 89548
rect 73804 89539 73856 89548
rect 73804 89505 73813 89539
rect 73813 89505 73847 89539
rect 73847 89505 73856 89539
rect 73804 89496 73856 89505
rect 87972 89564 88024 89616
rect 88156 89564 88208 89616
rect 81440 89496 81492 89548
rect 74632 89471 74684 89480
rect 70768 89360 70820 89412
rect 74632 89437 74641 89471
rect 74641 89437 74675 89471
rect 74675 89437 74684 89471
rect 74632 89428 74684 89437
rect 88248 89471 88300 89480
rect 88248 89437 88257 89471
rect 88257 89437 88291 89471
rect 88291 89437 88300 89471
rect 88248 89428 88300 89437
rect 88616 89471 88668 89480
rect 88616 89437 88625 89471
rect 88625 89437 88659 89471
rect 88659 89437 88668 89471
rect 88616 89428 88668 89437
rect 74908 89403 74960 89412
rect 74908 89369 74917 89403
rect 74917 89369 74951 89403
rect 74951 89369 74960 89403
rect 74908 89360 74960 89369
rect 52460 89292 52512 89344
rect 53196 89292 53248 89344
rect 4246 89190 4298 89242
rect 4310 89190 4362 89242
rect 4374 89190 4426 89242
rect 4438 89190 4490 89242
rect 34966 89190 35018 89242
rect 35030 89190 35082 89242
rect 35094 89190 35146 89242
rect 35158 89190 35210 89242
rect 65686 89190 65738 89242
rect 65750 89190 65802 89242
rect 65814 89190 65866 89242
rect 65878 89190 65930 89242
rect 96406 89190 96458 89242
rect 96470 89190 96522 89242
rect 96534 89190 96586 89242
rect 96598 89190 96650 89242
rect 53748 89088 53800 89140
rect 5080 89020 5132 89072
rect 2596 88884 2648 88936
rect 4068 88884 4120 88936
rect 6920 88791 6972 88800
rect 6920 88757 6929 88791
rect 6929 88757 6963 88791
rect 6963 88757 6972 88791
rect 6920 88748 6972 88757
rect 7564 88927 7616 88936
rect 7564 88893 7573 88927
rect 7573 88893 7607 88927
rect 7607 88893 7616 88927
rect 7564 88884 7616 88893
rect 7748 88884 7800 88936
rect 28172 88952 28224 89004
rect 82176 88952 82228 89004
rect 16304 88884 16356 88936
rect 13820 88816 13872 88868
rect 15108 88816 15160 88868
rect 17960 88927 18012 88936
rect 17960 88893 17969 88927
rect 17969 88893 18003 88927
rect 18003 88893 18012 88927
rect 17960 88884 18012 88893
rect 55036 88927 55088 88936
rect 55036 88893 55045 88927
rect 55045 88893 55079 88927
rect 55079 88893 55088 88927
rect 55036 88884 55088 88893
rect 19064 88791 19116 88800
rect 19064 88757 19073 88791
rect 19073 88757 19107 88791
rect 19107 88757 19116 88791
rect 19064 88748 19116 88757
rect 71136 88816 71188 88868
rect 50068 88748 50120 88800
rect 19606 88646 19658 88698
rect 19670 88646 19722 88698
rect 19734 88646 19786 88698
rect 19798 88646 19850 88698
rect 50326 88646 50378 88698
rect 50390 88646 50442 88698
rect 50454 88646 50506 88698
rect 50518 88646 50570 88698
rect 81046 88646 81098 88698
rect 81110 88646 81162 88698
rect 81174 88646 81226 88698
rect 81238 88646 81290 88698
rect 16120 88544 16172 88596
rect 16304 88544 16356 88596
rect 49700 88544 49752 88596
rect 7748 88476 7800 88528
rect 43812 88476 43864 88528
rect 2596 88408 2648 88460
rect 13820 88408 13872 88460
rect 15844 88451 15896 88460
rect 15844 88417 15853 88451
rect 15853 88417 15887 88451
rect 15887 88417 15896 88451
rect 15844 88408 15896 88417
rect 68284 88340 68336 88392
rect 77484 88204 77536 88256
rect 83832 88204 83884 88256
rect 4246 88102 4298 88154
rect 4310 88102 4362 88154
rect 4374 88102 4426 88154
rect 4438 88102 4490 88154
rect 34966 88102 35018 88154
rect 35030 88102 35082 88154
rect 35094 88102 35146 88154
rect 35158 88102 35210 88154
rect 65686 88102 65738 88154
rect 65750 88102 65802 88154
rect 65814 88102 65866 88154
rect 65878 88102 65930 88154
rect 96406 88102 96458 88154
rect 96470 88102 96522 88154
rect 96534 88102 96586 88154
rect 96598 88102 96650 88154
rect 41052 88000 41104 88052
rect 90272 88000 90324 88052
rect 77668 87932 77720 87984
rect 32496 87864 32548 87916
rect 89628 87864 89680 87916
rect 8300 87839 8352 87848
rect 8300 87805 8309 87839
rect 8309 87805 8343 87839
rect 8343 87805 8352 87839
rect 8300 87796 8352 87805
rect 77484 87796 77536 87848
rect 77576 87796 77628 87848
rect 77760 87796 77812 87848
rect 15752 87728 15804 87780
rect 22100 87728 22152 87780
rect 23388 87728 23440 87780
rect 34796 87728 34848 87780
rect 69756 87728 69808 87780
rect 29276 87660 29328 87712
rect 54484 87660 54536 87712
rect 19606 87558 19658 87610
rect 19670 87558 19722 87610
rect 19734 87558 19786 87610
rect 19798 87558 19850 87610
rect 50326 87558 50378 87610
rect 50390 87558 50442 87610
rect 50454 87558 50506 87610
rect 50518 87558 50570 87610
rect 81046 87558 81098 87610
rect 81110 87558 81162 87610
rect 81174 87558 81226 87610
rect 81238 87558 81290 87610
rect 10784 87388 10836 87440
rect 77576 87456 77628 87508
rect 84568 87456 84620 87508
rect 89628 87456 89680 87508
rect 89812 87456 89864 87508
rect 22100 87388 22152 87440
rect 44456 87388 44508 87440
rect 45100 87388 45152 87440
rect 27896 87363 27948 87372
rect 2320 87295 2372 87304
rect 2320 87261 2329 87295
rect 2329 87261 2363 87295
rect 2363 87261 2372 87295
rect 2320 87252 2372 87261
rect 1952 87159 2004 87168
rect 1952 87125 1961 87159
rect 1961 87125 1995 87159
rect 1995 87125 2004 87159
rect 1952 87116 2004 87125
rect 2412 87184 2464 87236
rect 27896 87329 27905 87363
rect 27905 87329 27939 87363
rect 27939 87329 27948 87363
rect 27896 87320 27948 87329
rect 29276 87320 29328 87372
rect 59912 87320 59964 87372
rect 73528 87363 73580 87372
rect 73528 87329 73537 87363
rect 73537 87329 73571 87363
rect 73571 87329 73580 87363
rect 73528 87320 73580 87329
rect 73896 87363 73948 87372
rect 73896 87329 73905 87363
rect 73905 87329 73939 87363
rect 73939 87329 73948 87363
rect 73896 87320 73948 87329
rect 74540 87320 74592 87372
rect 75368 87320 75420 87372
rect 89904 87363 89956 87372
rect 89904 87329 89913 87363
rect 89913 87329 89947 87363
rect 89947 87329 89956 87363
rect 89904 87320 89956 87329
rect 90272 87363 90324 87372
rect 90272 87329 90281 87363
rect 90281 87329 90315 87363
rect 90315 87329 90324 87363
rect 90272 87320 90324 87329
rect 28448 87295 28500 87304
rect 28448 87261 28457 87295
rect 28457 87261 28491 87295
rect 28491 87261 28500 87295
rect 28448 87252 28500 87261
rect 10140 87184 10192 87236
rect 73712 87252 73764 87304
rect 90088 87295 90140 87304
rect 90088 87261 90097 87295
rect 90097 87261 90131 87295
rect 90131 87261 90140 87295
rect 90088 87252 90140 87261
rect 89812 87227 89864 87236
rect 89812 87193 89821 87227
rect 89821 87193 89855 87227
rect 89855 87193 89864 87227
rect 91008 87227 91060 87236
rect 89812 87184 89864 87193
rect 91008 87193 91017 87227
rect 91017 87193 91051 87227
rect 91051 87193 91060 87227
rect 91008 87184 91060 87193
rect 35256 87116 35308 87168
rect 59912 87116 59964 87168
rect 4246 87014 4298 87066
rect 4310 87014 4362 87066
rect 4374 87014 4426 87066
rect 4438 87014 4490 87066
rect 34966 87014 35018 87066
rect 35030 87014 35082 87066
rect 35094 87014 35146 87066
rect 35158 87014 35210 87066
rect 65686 87014 65738 87066
rect 65750 87014 65802 87066
rect 65814 87014 65866 87066
rect 65878 87014 65930 87066
rect 96406 87014 96458 87066
rect 96470 87014 96522 87066
rect 96534 87014 96586 87066
rect 96598 87014 96650 87066
rect 29368 86912 29420 86964
rect 30196 86912 30248 86964
rect 12532 86844 12584 86896
rect 34520 86776 34572 86828
rect 12072 86751 12124 86760
rect 12072 86717 12081 86751
rect 12081 86717 12115 86751
rect 12115 86717 12124 86751
rect 12072 86708 12124 86717
rect 12808 86751 12860 86760
rect 12808 86717 12817 86751
rect 12817 86717 12851 86751
rect 12851 86717 12860 86751
rect 12808 86708 12860 86717
rect 29368 86708 29420 86760
rect 29736 86751 29788 86760
rect 29736 86717 29745 86751
rect 29745 86717 29779 86751
rect 29779 86717 29788 86751
rect 29736 86708 29788 86717
rect 64144 86708 64196 86760
rect 24216 86640 24268 86692
rect 46848 86640 46900 86692
rect 90548 86572 90600 86624
rect 19606 86470 19658 86522
rect 19670 86470 19722 86522
rect 19734 86470 19786 86522
rect 19798 86470 19850 86522
rect 50326 86470 50378 86522
rect 50390 86470 50442 86522
rect 50454 86470 50506 86522
rect 50518 86470 50570 86522
rect 81046 86470 81098 86522
rect 81110 86470 81162 86522
rect 81174 86470 81226 86522
rect 81238 86470 81290 86522
rect 12072 86300 12124 86352
rect 46296 86300 46348 86352
rect 54668 86300 54720 86352
rect 74632 86300 74684 86352
rect 43536 86275 43588 86284
rect 43536 86241 43545 86275
rect 43545 86241 43579 86275
rect 43579 86241 43588 86275
rect 43536 86232 43588 86241
rect 49056 86232 49108 86284
rect 73804 86232 73856 86284
rect 44916 86164 44968 86216
rect 83096 86164 83148 86216
rect 84568 86207 84620 86216
rect 84568 86173 84577 86207
rect 84577 86173 84611 86207
rect 84611 86173 84620 86207
rect 84568 86164 84620 86173
rect 82820 86028 82872 86080
rect 90272 86028 90324 86080
rect 97632 86028 97684 86080
rect 4246 85926 4298 85978
rect 4310 85926 4362 85978
rect 4374 85926 4426 85978
rect 4438 85926 4490 85978
rect 34966 85926 35018 85978
rect 35030 85926 35082 85978
rect 35094 85926 35146 85978
rect 35158 85926 35210 85978
rect 65686 85926 65738 85978
rect 65750 85926 65802 85978
rect 65814 85926 65866 85978
rect 65878 85926 65930 85978
rect 96406 85926 96458 85978
rect 96470 85926 96522 85978
rect 96534 85926 96586 85978
rect 96598 85926 96650 85978
rect 82084 85620 82136 85672
rect 23664 85595 23716 85604
rect 23664 85561 23673 85595
rect 23673 85561 23707 85595
rect 23707 85561 23716 85595
rect 23664 85552 23716 85561
rect 24400 85595 24452 85604
rect 24400 85561 24409 85595
rect 24409 85561 24443 85595
rect 24443 85561 24452 85595
rect 24400 85552 24452 85561
rect 45008 85552 45060 85604
rect 30380 85484 30432 85536
rect 31300 85484 31352 85536
rect 19606 85382 19658 85434
rect 19670 85382 19722 85434
rect 19734 85382 19786 85434
rect 19798 85382 19850 85434
rect 50326 85382 50378 85434
rect 50390 85382 50442 85434
rect 50454 85382 50506 85434
rect 50518 85382 50570 85434
rect 81046 85382 81098 85434
rect 81110 85382 81162 85434
rect 81174 85382 81226 85434
rect 81238 85382 81290 85434
rect 10508 85280 10560 85332
rect 10600 85212 10652 85264
rect 5080 85187 5132 85196
rect 5080 85153 5089 85187
rect 5089 85153 5123 85187
rect 5123 85153 5132 85187
rect 5080 85144 5132 85153
rect 10048 85144 10100 85196
rect 10508 85187 10560 85196
rect 10508 85153 10517 85187
rect 10517 85153 10551 85187
rect 10551 85153 10560 85187
rect 14648 85280 14700 85332
rect 31852 85280 31904 85332
rect 45468 85280 45520 85332
rect 23664 85212 23716 85264
rect 30012 85212 30064 85264
rect 10508 85144 10560 85153
rect 6460 85076 6512 85128
rect 9588 85119 9640 85128
rect 9588 85085 9597 85119
rect 9597 85085 9631 85119
rect 9631 85085 9640 85119
rect 9588 85076 9640 85085
rect 10232 85119 10284 85128
rect 10232 85085 10241 85119
rect 10241 85085 10275 85119
rect 10275 85085 10284 85119
rect 10232 85076 10284 85085
rect 10324 85076 10376 85128
rect 32588 85144 32640 85196
rect 46296 85187 46348 85196
rect 46296 85153 46305 85187
rect 46305 85153 46339 85187
rect 46339 85153 46348 85187
rect 46296 85144 46348 85153
rect 50160 85280 50212 85332
rect 74908 85280 74960 85332
rect 53932 85212 53984 85264
rect 95700 85212 95752 85264
rect 46756 85144 46808 85196
rect 56968 85144 57020 85196
rect 72516 85187 72568 85196
rect 72516 85153 72525 85187
rect 72525 85153 72559 85187
rect 72559 85153 72568 85187
rect 72516 85144 72568 85153
rect 30380 85076 30432 85128
rect 45192 85076 45244 85128
rect 46572 85119 46624 85128
rect 46572 85085 46581 85119
rect 46581 85085 46615 85119
rect 46615 85085 46624 85119
rect 46572 85076 46624 85085
rect 46940 85076 46992 85128
rect 79508 85076 79560 85128
rect 10600 84940 10652 84992
rect 34152 84940 34204 84992
rect 46480 84940 46532 84992
rect 82636 85008 82688 85060
rect 61108 84940 61160 84992
rect 4246 84838 4298 84890
rect 4310 84838 4362 84890
rect 4374 84838 4426 84890
rect 4438 84838 4490 84890
rect 34966 84838 35018 84890
rect 35030 84838 35082 84890
rect 35094 84838 35146 84890
rect 35158 84838 35210 84890
rect 65686 84838 65738 84890
rect 65750 84838 65802 84890
rect 65814 84838 65866 84890
rect 65878 84838 65930 84890
rect 96406 84838 96458 84890
rect 96470 84838 96522 84890
rect 96534 84838 96586 84890
rect 96598 84838 96650 84890
rect 42064 84736 42116 84788
rect 39856 84668 39908 84720
rect 50160 84668 50212 84720
rect 62304 84575 62356 84584
rect 62304 84541 62313 84575
rect 62313 84541 62347 84575
rect 62347 84541 62356 84575
rect 62304 84532 62356 84541
rect 85764 84575 85816 84584
rect 85764 84541 85773 84575
rect 85773 84541 85807 84575
rect 85807 84541 85816 84575
rect 85764 84532 85816 84541
rect 85948 84439 86000 84448
rect 85948 84405 85957 84439
rect 85957 84405 85991 84439
rect 85991 84405 86000 84439
rect 85948 84396 86000 84405
rect 19606 84294 19658 84346
rect 19670 84294 19722 84346
rect 19734 84294 19786 84346
rect 19798 84294 19850 84346
rect 50326 84294 50378 84346
rect 50390 84294 50442 84346
rect 50454 84294 50506 84346
rect 50518 84294 50570 84346
rect 81046 84294 81098 84346
rect 81110 84294 81162 84346
rect 81174 84294 81226 84346
rect 81238 84294 81290 84346
rect 65984 84124 66036 84176
rect 47584 84056 47636 84108
rect 60372 83988 60424 84040
rect 79324 83988 79376 84040
rect 85304 84031 85356 84040
rect 85304 83997 85313 84031
rect 85313 83997 85347 84031
rect 85347 83997 85356 84031
rect 85304 83988 85356 83997
rect 85672 84031 85724 84040
rect 85672 83997 85681 84031
rect 85681 83997 85715 84031
rect 85715 83997 85724 84031
rect 85672 83988 85724 83997
rect 86224 84099 86276 84108
rect 86224 84065 86233 84099
rect 86233 84065 86267 84099
rect 86267 84065 86276 84099
rect 86224 84056 86276 84065
rect 86132 84031 86184 84040
rect 86132 83997 86141 84031
rect 86141 83997 86175 84031
rect 86175 83997 86184 84031
rect 86132 83988 86184 83997
rect 88524 83988 88576 84040
rect 62028 83920 62080 83972
rect 65524 83852 65576 83904
rect 66904 83852 66956 83904
rect 67548 83852 67600 83904
rect 96896 83852 96948 83904
rect 4246 83750 4298 83802
rect 4310 83750 4362 83802
rect 4374 83750 4426 83802
rect 4438 83750 4490 83802
rect 34966 83750 35018 83802
rect 35030 83750 35082 83802
rect 35094 83750 35146 83802
rect 35158 83750 35210 83802
rect 65686 83750 65738 83802
rect 65750 83750 65802 83802
rect 65814 83750 65866 83802
rect 65878 83750 65930 83802
rect 96406 83750 96458 83802
rect 96470 83750 96522 83802
rect 96534 83750 96586 83802
rect 96598 83750 96650 83802
rect 71044 83648 71096 83700
rect 12808 83580 12860 83632
rect 21088 83580 21140 83632
rect 20352 83512 20404 83564
rect 31208 83512 31260 83564
rect 79324 83648 79376 83700
rect 88524 83648 88576 83700
rect 86224 83512 86276 83564
rect 64328 83444 64380 83496
rect 71136 83444 71188 83496
rect 86132 83444 86184 83496
rect 97172 83376 97224 83428
rect 98000 83351 98052 83360
rect 98000 83317 98009 83351
rect 98009 83317 98043 83351
rect 98043 83317 98052 83351
rect 98000 83308 98052 83317
rect 19606 83206 19658 83258
rect 19670 83206 19722 83258
rect 19734 83206 19786 83258
rect 19798 83206 19850 83258
rect 50326 83206 50378 83258
rect 50390 83206 50442 83258
rect 50454 83206 50506 83258
rect 50518 83206 50570 83258
rect 81046 83206 81098 83258
rect 81110 83206 81162 83258
rect 81174 83206 81226 83258
rect 81238 83206 81290 83258
rect 26608 82968 26660 83020
rect 76564 83011 76616 83020
rect 76564 82977 76573 83011
rect 76573 82977 76607 83011
rect 76607 82977 76616 83011
rect 76564 82968 76616 82977
rect 75644 82943 75696 82952
rect 75644 82909 75653 82943
rect 75653 82909 75687 82943
rect 75687 82909 75696 82943
rect 75644 82900 75696 82909
rect 76012 82943 76064 82952
rect 76012 82909 76021 82943
rect 76021 82909 76055 82943
rect 76055 82909 76064 82943
rect 76012 82900 76064 82909
rect 76472 82943 76524 82952
rect 76472 82909 76481 82943
rect 76481 82909 76515 82943
rect 76515 82909 76524 82943
rect 76472 82900 76524 82909
rect 4246 82662 4298 82714
rect 4310 82662 4362 82714
rect 4374 82662 4426 82714
rect 4438 82662 4490 82714
rect 34966 82662 35018 82714
rect 35030 82662 35082 82714
rect 35094 82662 35146 82714
rect 35158 82662 35210 82714
rect 65686 82662 65738 82714
rect 65750 82662 65802 82714
rect 65814 82662 65866 82714
rect 65878 82662 65930 82714
rect 96406 82662 96458 82714
rect 96470 82662 96522 82714
rect 96534 82662 96586 82714
rect 96598 82662 96650 82714
rect 53840 82424 53892 82476
rect 68836 82424 68888 82476
rect 6920 82288 6972 82340
rect 39488 82288 39540 82340
rect 41880 82288 41932 82340
rect 61200 82356 61252 82408
rect 65984 82356 66036 82408
rect 14648 82220 14700 82272
rect 71044 82220 71096 82272
rect 19606 82118 19658 82170
rect 19670 82118 19722 82170
rect 19734 82118 19786 82170
rect 19798 82118 19850 82170
rect 50326 82118 50378 82170
rect 50390 82118 50442 82170
rect 50454 82118 50506 82170
rect 50518 82118 50570 82170
rect 81046 82118 81098 82170
rect 81110 82118 81162 82170
rect 81174 82118 81226 82170
rect 81238 82118 81290 82170
rect 91744 82016 91796 82068
rect 73804 81948 73856 82000
rect 74080 81923 74132 81932
rect 74080 81889 74089 81923
rect 74089 81889 74123 81923
rect 74123 81889 74132 81923
rect 74080 81880 74132 81889
rect 54300 81812 54352 81864
rect 54484 81812 54536 81864
rect 83004 81923 83056 81932
rect 83004 81889 83013 81923
rect 83013 81889 83047 81923
rect 83047 81889 83056 81923
rect 83004 81880 83056 81889
rect 92572 81812 92624 81864
rect 89904 81744 89956 81796
rect 89720 81676 89772 81728
rect 95240 81719 95292 81728
rect 95240 81685 95249 81719
rect 95249 81685 95283 81719
rect 95283 81685 95292 81719
rect 95240 81676 95292 81685
rect 4246 81574 4298 81626
rect 4310 81574 4362 81626
rect 4374 81574 4426 81626
rect 4438 81574 4490 81626
rect 34966 81574 35018 81626
rect 35030 81574 35082 81626
rect 35094 81574 35146 81626
rect 35158 81574 35210 81626
rect 65686 81574 65738 81626
rect 65750 81574 65802 81626
rect 65814 81574 65866 81626
rect 65878 81574 65930 81626
rect 96406 81574 96458 81626
rect 96470 81574 96522 81626
rect 96534 81574 96586 81626
rect 96598 81574 96650 81626
rect 73804 81472 73856 81524
rect 74172 81472 74224 81524
rect 95240 81472 95292 81524
rect 7012 81336 7064 81388
rect 8208 81336 8260 81388
rect 32496 81200 32548 81252
rect 32588 81200 32640 81252
rect 83004 81200 83056 81252
rect 83648 81200 83700 81252
rect 27620 81175 27672 81184
rect 27620 81141 27629 81175
rect 27629 81141 27663 81175
rect 27663 81141 27672 81175
rect 27620 81132 27672 81141
rect 29920 81175 29972 81184
rect 29920 81141 29929 81175
rect 29929 81141 29963 81175
rect 29963 81141 29972 81175
rect 29920 81132 29972 81141
rect 19606 81030 19658 81082
rect 19670 81030 19722 81082
rect 19734 81030 19786 81082
rect 19798 81030 19850 81082
rect 50326 81030 50378 81082
rect 50390 81030 50442 81082
rect 50454 81030 50506 81082
rect 50518 81030 50570 81082
rect 81046 81030 81098 81082
rect 81110 81030 81162 81082
rect 81174 81030 81226 81082
rect 81238 81030 81290 81082
rect 74080 80903 74132 80912
rect 74080 80869 74089 80903
rect 74089 80869 74123 80903
rect 74123 80869 74132 80903
rect 74080 80860 74132 80869
rect 84292 80903 84344 80912
rect 84292 80869 84301 80903
rect 84301 80869 84335 80903
rect 84335 80869 84344 80903
rect 84292 80860 84344 80869
rect 10232 80588 10284 80640
rect 12900 80588 12952 80640
rect 31392 80588 31444 80640
rect 84384 80724 84436 80776
rect 84660 80767 84712 80776
rect 84660 80733 84669 80767
rect 84669 80733 84703 80767
rect 84703 80733 84712 80767
rect 84660 80724 84712 80733
rect 84476 80631 84528 80640
rect 84476 80597 84500 80631
rect 84500 80597 84528 80631
rect 84476 80588 84528 80597
rect 84752 80631 84804 80640
rect 84752 80597 84761 80631
rect 84761 80597 84795 80631
rect 84795 80597 84804 80631
rect 84752 80588 84804 80597
rect 4246 80486 4298 80538
rect 4310 80486 4362 80538
rect 4374 80486 4426 80538
rect 4438 80486 4490 80538
rect 34966 80486 35018 80538
rect 35030 80486 35082 80538
rect 35094 80486 35146 80538
rect 35158 80486 35210 80538
rect 65686 80486 65738 80538
rect 65750 80486 65802 80538
rect 65814 80486 65866 80538
rect 65878 80486 65930 80538
rect 96406 80486 96458 80538
rect 96470 80486 96522 80538
rect 96534 80486 96586 80538
rect 96598 80486 96650 80538
rect 8208 80248 8260 80300
rect 29644 80180 29696 80232
rect 49608 80223 49660 80232
rect 49608 80189 49617 80223
rect 49617 80189 49651 80223
rect 49651 80189 49660 80223
rect 49608 80180 49660 80189
rect 49792 80223 49844 80232
rect 49792 80189 49801 80223
rect 49801 80189 49835 80223
rect 49835 80189 49844 80223
rect 49792 80180 49844 80189
rect 29368 80044 29420 80096
rect 30840 80112 30892 80164
rect 49700 80112 49752 80164
rect 50068 80180 50120 80232
rect 50160 80180 50212 80232
rect 50712 80112 50764 80164
rect 40776 80044 40828 80096
rect 41328 80044 41380 80096
rect 50804 80087 50856 80096
rect 50804 80053 50813 80087
rect 50813 80053 50847 80087
rect 50847 80053 50856 80087
rect 50804 80044 50856 80053
rect 75644 80044 75696 80096
rect 82176 80044 82228 80096
rect 19606 79942 19658 79994
rect 19670 79942 19722 79994
rect 19734 79942 19786 79994
rect 19798 79942 19850 79994
rect 50326 79942 50378 79994
rect 50390 79942 50442 79994
rect 50454 79942 50506 79994
rect 50518 79942 50570 79994
rect 81046 79942 81098 79994
rect 81110 79942 81162 79994
rect 81174 79942 81226 79994
rect 81238 79942 81290 79994
rect 31024 79840 31076 79892
rect 42892 79815 42944 79824
rect 29184 79704 29236 79756
rect 42616 79747 42668 79756
rect 42616 79713 42625 79747
rect 42625 79713 42659 79747
rect 42659 79713 42668 79747
rect 42616 79704 42668 79713
rect 42892 79781 42901 79815
rect 42901 79781 42935 79815
rect 42935 79781 42944 79815
rect 42892 79772 42944 79781
rect 30472 79636 30524 79688
rect 3976 79500 4028 79552
rect 29184 79500 29236 79552
rect 30380 79500 30432 79552
rect 43168 79747 43220 79756
rect 43168 79713 43194 79747
rect 43194 79713 43220 79747
rect 43168 79704 43220 79713
rect 76472 79704 76524 79756
rect 78128 79636 78180 79688
rect 46296 79568 46348 79620
rect 62120 79568 62172 79620
rect 80796 79568 80848 79620
rect 89168 79704 89220 79756
rect 89628 79747 89680 79756
rect 89628 79713 89637 79747
rect 89637 79713 89671 79747
rect 89671 79713 89680 79747
rect 89628 79704 89680 79713
rect 89352 79679 89404 79688
rect 89352 79645 89361 79679
rect 89361 79645 89395 79679
rect 89395 79645 89404 79679
rect 89352 79636 89404 79645
rect 89812 79611 89864 79620
rect 89812 79577 89821 79611
rect 89821 79577 89855 79611
rect 89855 79577 89864 79611
rect 89812 79568 89864 79577
rect 43444 79543 43496 79552
rect 43444 79509 43453 79543
rect 43453 79509 43487 79543
rect 43487 79509 43496 79543
rect 43444 79500 43496 79509
rect 76012 79500 76064 79552
rect 89168 79500 89220 79552
rect 89352 79500 89404 79552
rect 4246 79398 4298 79450
rect 4310 79398 4362 79450
rect 4374 79398 4426 79450
rect 4438 79398 4490 79450
rect 34966 79398 35018 79450
rect 35030 79398 35082 79450
rect 35094 79398 35146 79450
rect 35158 79398 35210 79450
rect 65686 79398 65738 79450
rect 65750 79398 65802 79450
rect 65814 79398 65866 79450
rect 65878 79398 65930 79450
rect 96406 79398 96458 79450
rect 96470 79398 96522 79450
rect 96534 79398 96586 79450
rect 96598 79398 96650 79450
rect 6828 79296 6880 79348
rect 82820 79296 82872 79348
rect 10324 79228 10376 79280
rect 30380 79228 30432 79280
rect 6276 79160 6328 79212
rect 12900 79160 12952 79212
rect 30472 79160 30524 79212
rect 86224 79160 86276 79212
rect 3976 79135 4028 79144
rect 3976 79101 3985 79135
rect 3985 79101 4019 79135
rect 4019 79101 4028 79135
rect 3976 79092 4028 79101
rect 4528 79092 4580 79144
rect 4712 79135 4764 79144
rect 4712 79101 4721 79135
rect 4721 79101 4755 79135
rect 4755 79101 4764 79135
rect 4712 79092 4764 79101
rect 28540 79092 28592 79144
rect 62120 79092 62172 79144
rect 62856 79092 62908 79144
rect 96896 79135 96948 79144
rect 96896 79101 96905 79135
rect 96905 79101 96939 79135
rect 96939 79101 96948 79135
rect 96896 79092 96948 79101
rect 97080 79135 97132 79144
rect 97080 79101 97089 79135
rect 97089 79101 97123 79135
rect 97123 79101 97132 79135
rect 97080 79092 97132 79101
rect 97448 79135 97500 79144
rect 97448 79101 97457 79135
rect 97457 79101 97491 79135
rect 97491 79101 97500 79135
rect 97448 79092 97500 79101
rect 83096 79024 83148 79076
rect 11612 78956 11664 79008
rect 19606 78854 19658 78906
rect 19670 78854 19722 78906
rect 19734 78854 19786 78906
rect 19798 78854 19850 78906
rect 50326 78854 50378 78906
rect 50390 78854 50442 78906
rect 50454 78854 50506 78906
rect 50518 78854 50570 78906
rect 81046 78854 81098 78906
rect 81110 78854 81162 78906
rect 81174 78854 81226 78906
rect 81238 78854 81290 78906
rect 4712 78752 4764 78804
rect 20720 78752 20772 78804
rect 25780 78752 25832 78804
rect 11520 78659 11572 78668
rect 11520 78625 11529 78659
rect 11529 78625 11563 78659
rect 11563 78625 11572 78659
rect 11520 78616 11572 78625
rect 17040 78616 17092 78668
rect 17132 78616 17184 78668
rect 17592 78684 17644 78736
rect 17776 78616 17828 78668
rect 17408 78548 17460 78600
rect 3884 78480 3936 78532
rect 24032 78616 24084 78668
rect 30472 78659 30524 78668
rect 30472 78625 30481 78659
rect 30481 78625 30515 78659
rect 30515 78625 30524 78659
rect 30472 78616 30524 78625
rect 27896 78548 27948 78600
rect 30380 78591 30432 78600
rect 30380 78557 30389 78591
rect 30389 78557 30423 78591
rect 30423 78557 30432 78591
rect 82728 78616 82780 78668
rect 98000 78616 98052 78668
rect 30380 78548 30432 78557
rect 66076 78548 66128 78600
rect 49056 78480 49108 78532
rect 17040 78455 17092 78464
rect 17040 78421 17049 78455
rect 17049 78421 17083 78455
rect 17083 78421 17092 78455
rect 17040 78412 17092 78421
rect 17224 78455 17276 78464
rect 17224 78421 17233 78455
rect 17233 78421 17267 78455
rect 17267 78421 17276 78455
rect 17224 78412 17276 78421
rect 31116 78412 31168 78464
rect 90364 78412 90416 78464
rect 4246 78310 4298 78362
rect 4310 78310 4362 78362
rect 4374 78310 4426 78362
rect 4438 78310 4490 78362
rect 34966 78310 35018 78362
rect 35030 78310 35082 78362
rect 35094 78310 35146 78362
rect 35158 78310 35210 78362
rect 65686 78310 65738 78362
rect 65750 78310 65802 78362
rect 65814 78310 65866 78362
rect 65878 78310 65930 78362
rect 96406 78310 96458 78362
rect 96470 78310 96522 78362
rect 96534 78310 96586 78362
rect 96598 78310 96650 78362
rect 66168 78208 66220 78260
rect 11520 78140 11572 78192
rect 58624 78140 58676 78192
rect 17040 78072 17092 78124
rect 48964 78072 49016 78124
rect 23664 78047 23716 78056
rect 23664 78013 23673 78047
rect 23673 78013 23707 78047
rect 23707 78013 23716 78047
rect 23664 78004 23716 78013
rect 50896 77868 50948 77920
rect 53656 77868 53708 77920
rect 76748 77868 76800 77920
rect 82728 78047 82780 78056
rect 82268 77979 82320 77988
rect 82268 77945 82277 77979
rect 82277 77945 82311 77979
rect 82311 77945 82320 77979
rect 82268 77936 82320 77945
rect 82728 78013 82737 78047
rect 82737 78013 82771 78047
rect 82771 78013 82780 78047
rect 82728 78004 82780 78013
rect 83096 78047 83148 78056
rect 83096 78013 83105 78047
rect 83105 78013 83139 78047
rect 83139 78013 83148 78047
rect 83096 78004 83148 78013
rect 84200 77936 84252 77988
rect 84568 77936 84620 77988
rect 92572 77936 92624 77988
rect 19606 77766 19658 77818
rect 19670 77766 19722 77818
rect 19734 77766 19786 77818
rect 19798 77766 19850 77818
rect 50326 77766 50378 77818
rect 50390 77766 50442 77818
rect 50454 77766 50506 77818
rect 50518 77766 50570 77818
rect 81046 77766 81098 77818
rect 81110 77766 81162 77818
rect 81174 77766 81226 77818
rect 81238 77766 81290 77818
rect 20720 77639 20772 77648
rect 20720 77605 20729 77639
rect 20729 77605 20763 77639
rect 20763 77605 20772 77639
rect 20720 77596 20772 77605
rect 25964 77571 26016 77580
rect 25964 77537 25973 77571
rect 25973 77537 26007 77571
rect 26007 77537 26016 77571
rect 25964 77528 26016 77537
rect 26148 77571 26200 77580
rect 26148 77537 26156 77571
rect 26156 77537 26190 77571
rect 26190 77537 26200 77571
rect 28448 77664 28500 77716
rect 61384 77664 61436 77716
rect 62764 77664 62816 77716
rect 83096 77664 83148 77716
rect 26148 77528 26200 77537
rect 23388 77460 23440 77512
rect 96804 77596 96856 77648
rect 26516 77571 26568 77580
rect 26516 77537 26525 77571
rect 26525 77537 26559 77571
rect 26559 77537 26568 77571
rect 26516 77528 26568 77537
rect 93768 77528 93820 77580
rect 26424 77324 26476 77376
rect 26608 77367 26660 77376
rect 26608 77333 26617 77367
rect 26617 77333 26651 77367
rect 26651 77333 26660 77367
rect 26608 77324 26660 77333
rect 4246 77222 4298 77274
rect 4310 77222 4362 77274
rect 4374 77222 4426 77274
rect 4438 77222 4490 77274
rect 34966 77222 35018 77274
rect 35030 77222 35082 77274
rect 35094 77222 35146 77274
rect 35158 77222 35210 77274
rect 65686 77222 65738 77274
rect 65750 77222 65802 77274
rect 65814 77222 65866 77274
rect 65878 77222 65930 77274
rect 96406 77222 96458 77274
rect 96470 77222 96522 77274
rect 96534 77222 96586 77274
rect 96598 77222 96650 77274
rect 23388 77120 23440 77172
rect 20720 77095 20772 77104
rect 20720 77061 20729 77095
rect 20729 77061 20763 77095
rect 20763 77061 20772 77095
rect 20720 77052 20772 77061
rect 36360 77120 36412 77172
rect 80796 77052 80848 77104
rect 78128 76984 78180 77036
rect 28816 76959 28868 76968
rect 21364 76848 21416 76900
rect 28816 76925 28825 76959
rect 28825 76925 28859 76959
rect 28859 76925 28868 76959
rect 28816 76916 28868 76925
rect 29184 76959 29236 76968
rect 29184 76925 29193 76959
rect 29193 76925 29227 76959
rect 29227 76925 29236 76959
rect 29184 76916 29236 76925
rect 29368 76959 29420 76968
rect 29368 76925 29377 76959
rect 29377 76925 29411 76959
rect 29411 76925 29420 76959
rect 29368 76916 29420 76925
rect 43812 76959 43864 76968
rect 43812 76925 43821 76959
rect 43821 76925 43855 76959
rect 43855 76925 43864 76959
rect 43812 76916 43864 76925
rect 54484 76959 54536 76968
rect 54484 76925 54493 76959
rect 54493 76925 54527 76959
rect 54527 76925 54536 76959
rect 54484 76916 54536 76925
rect 21272 76780 21324 76832
rect 32588 76848 32640 76900
rect 29644 76823 29696 76832
rect 29644 76789 29653 76823
rect 29653 76789 29687 76823
rect 29687 76789 29696 76823
rect 29644 76780 29696 76789
rect 79416 76780 79468 76832
rect 19606 76678 19658 76730
rect 19670 76678 19722 76730
rect 19734 76678 19786 76730
rect 19798 76678 19850 76730
rect 50326 76678 50378 76730
rect 50390 76678 50442 76730
rect 50454 76678 50506 76730
rect 50518 76678 50570 76730
rect 81046 76678 81098 76730
rect 81110 76678 81162 76730
rect 81174 76678 81226 76730
rect 81238 76678 81290 76730
rect 24492 76576 24544 76628
rect 55588 76576 55640 76628
rect 56232 76576 56284 76628
rect 58072 76619 58124 76628
rect 58072 76585 58081 76619
rect 58081 76585 58115 76619
rect 58115 76585 58124 76619
rect 58072 76576 58124 76585
rect 58348 76576 58400 76628
rect 71780 76508 71832 76560
rect 72516 76508 72568 76560
rect 79784 76508 79836 76560
rect 3332 76440 3384 76492
rect 21364 76440 21416 76492
rect 30564 76483 30616 76492
rect 30564 76449 30573 76483
rect 30573 76449 30607 76483
rect 30607 76449 30616 76483
rect 30564 76440 30616 76449
rect 31392 76440 31444 76492
rect 47676 76440 47728 76492
rect 93584 76440 93636 76492
rect 13820 76372 13872 76424
rect 15108 76372 15160 76424
rect 31116 76415 31168 76424
rect 31116 76381 31125 76415
rect 31125 76381 31159 76415
rect 31159 76381 31168 76415
rect 31116 76372 31168 76381
rect 56692 76415 56744 76424
rect 56692 76381 56701 76415
rect 56701 76381 56735 76415
rect 56735 76381 56744 76415
rect 56692 76372 56744 76381
rect 92572 76372 92624 76424
rect 24124 76304 24176 76356
rect 8944 76236 8996 76288
rect 37556 76279 37608 76288
rect 37556 76245 37565 76279
rect 37565 76245 37599 76279
rect 37599 76245 37608 76279
rect 37556 76236 37608 76245
rect 93584 76279 93636 76288
rect 93584 76245 93593 76279
rect 93593 76245 93627 76279
rect 93627 76245 93636 76279
rect 93584 76236 93636 76245
rect 95148 76279 95200 76288
rect 95148 76245 95157 76279
rect 95157 76245 95191 76279
rect 95191 76245 95200 76279
rect 95148 76236 95200 76245
rect 4246 76134 4298 76186
rect 4310 76134 4362 76186
rect 4374 76134 4426 76186
rect 4438 76134 4490 76186
rect 34966 76134 35018 76186
rect 35030 76134 35082 76186
rect 35094 76134 35146 76186
rect 35158 76134 35210 76186
rect 65686 76134 65738 76186
rect 65750 76134 65802 76186
rect 65814 76134 65866 76186
rect 65878 76134 65930 76186
rect 96406 76134 96458 76186
rect 96470 76134 96522 76186
rect 96534 76134 96586 76186
rect 96598 76134 96650 76186
rect 56232 76032 56284 76084
rect 95148 76032 95200 76084
rect 5356 75964 5408 76016
rect 71780 75896 71832 75948
rect 5080 75871 5132 75880
rect 5080 75837 5089 75871
rect 5089 75837 5123 75871
rect 5123 75837 5132 75871
rect 5080 75828 5132 75837
rect 15016 75828 15068 75880
rect 35440 75828 35492 75880
rect 38016 75828 38068 75880
rect 38660 75828 38712 75880
rect 44088 75871 44140 75880
rect 44088 75837 44097 75871
rect 44097 75837 44131 75871
rect 44131 75837 44140 75871
rect 44088 75828 44140 75837
rect 9680 75760 9732 75812
rect 30564 75760 30616 75812
rect 19606 75590 19658 75642
rect 19670 75590 19722 75642
rect 19734 75590 19786 75642
rect 19798 75590 19850 75642
rect 50326 75590 50378 75642
rect 50390 75590 50442 75642
rect 50454 75590 50506 75642
rect 50518 75590 50570 75642
rect 81046 75590 81098 75642
rect 81110 75590 81162 75642
rect 81174 75590 81226 75642
rect 81238 75590 81290 75642
rect 57520 75420 57572 75472
rect 68560 75420 68612 75472
rect 12440 75352 12492 75404
rect 12624 75352 12676 75404
rect 43444 75352 43496 75404
rect 54484 75352 54536 75404
rect 94504 75352 94556 75404
rect 17776 75284 17828 75336
rect 68376 75284 68428 75336
rect 28540 75216 28592 75268
rect 87880 75216 87932 75268
rect 25872 75148 25924 75200
rect 91100 75148 91152 75200
rect 93952 75148 94004 75200
rect 4246 75046 4298 75098
rect 4310 75046 4362 75098
rect 4374 75046 4426 75098
rect 4438 75046 4490 75098
rect 34966 75046 35018 75098
rect 35030 75046 35082 75098
rect 35094 75046 35146 75098
rect 35158 75046 35210 75098
rect 65686 75046 65738 75098
rect 65750 75046 65802 75098
rect 65814 75046 65866 75098
rect 65878 75046 65930 75098
rect 96406 75046 96458 75098
rect 96470 75046 96522 75098
rect 96534 75046 96586 75098
rect 96598 75046 96650 75098
rect 13728 74808 13780 74860
rect 72424 74808 72476 74860
rect 2872 74783 2924 74792
rect 2872 74749 2881 74783
rect 2881 74749 2915 74783
rect 2915 74749 2924 74783
rect 2872 74740 2924 74749
rect 72240 74740 72292 74792
rect 72700 74740 72752 74792
rect 72884 74783 72936 74792
rect 72884 74749 72893 74783
rect 72893 74749 72927 74783
rect 72927 74749 72936 74783
rect 72884 74740 72936 74749
rect 72976 74783 73028 74792
rect 72976 74749 72985 74783
rect 72985 74749 73019 74783
rect 73019 74749 73028 74783
rect 72976 74740 73028 74749
rect 79324 74672 79376 74724
rect 12440 74604 12492 74656
rect 44180 74604 44232 74656
rect 78312 74604 78364 74656
rect 97080 74604 97132 74656
rect 19606 74502 19658 74554
rect 19670 74502 19722 74554
rect 19734 74502 19786 74554
rect 19798 74502 19850 74554
rect 50326 74502 50378 74554
rect 50390 74502 50442 74554
rect 50454 74502 50506 74554
rect 50518 74502 50570 74554
rect 81046 74502 81098 74554
rect 81110 74502 81162 74554
rect 81174 74502 81226 74554
rect 81238 74502 81290 74554
rect 32496 74400 32548 74452
rect 44088 74400 44140 74452
rect 51448 74307 51500 74316
rect 51448 74273 51457 74307
rect 51457 74273 51491 74307
rect 51491 74273 51500 74307
rect 51448 74264 51500 74273
rect 53288 74400 53340 74452
rect 53380 74332 53432 74384
rect 52000 74307 52052 74316
rect 52000 74273 52009 74307
rect 52009 74273 52043 74307
rect 52043 74273 52052 74307
rect 52000 74264 52052 74273
rect 56692 74307 56744 74316
rect 56692 74273 56701 74307
rect 56701 74273 56735 74307
rect 56735 74273 56744 74307
rect 56692 74264 56744 74273
rect 61936 74264 61988 74316
rect 78312 74307 78364 74316
rect 78312 74273 78321 74307
rect 78321 74273 78355 74307
rect 78355 74273 78364 74307
rect 78312 74264 78364 74273
rect 52460 74196 52512 74248
rect 56968 74239 57020 74248
rect 56968 74205 56977 74239
rect 56977 74205 57011 74239
rect 57011 74205 57020 74239
rect 56968 74196 57020 74205
rect 78496 74239 78548 74248
rect 78496 74205 78505 74239
rect 78505 74205 78539 74239
rect 78539 74205 78548 74239
rect 78496 74196 78548 74205
rect 96068 74196 96120 74248
rect 25044 74060 25096 74112
rect 26792 74060 26844 74112
rect 52092 74103 52144 74112
rect 52092 74069 52101 74103
rect 52101 74069 52135 74103
rect 52135 74069 52144 74103
rect 52092 74060 52144 74069
rect 4246 73958 4298 74010
rect 4310 73958 4362 74010
rect 4374 73958 4426 74010
rect 4438 73958 4490 74010
rect 34966 73958 35018 74010
rect 35030 73958 35082 74010
rect 35094 73958 35146 74010
rect 35158 73958 35210 74010
rect 65686 73958 65738 74010
rect 65750 73958 65802 74010
rect 65814 73958 65866 74010
rect 65878 73958 65930 74010
rect 96406 73958 96458 74010
rect 96470 73958 96522 74010
rect 96534 73958 96586 74010
rect 96598 73958 96650 74010
rect 16304 73856 16356 73908
rect 17868 73856 17920 73908
rect 25044 73856 25096 73908
rect 39580 73856 39632 73908
rect 56968 73856 57020 73908
rect 26056 73788 26108 73840
rect 38844 73788 38896 73840
rect 39948 73788 40000 73840
rect 45284 73788 45336 73840
rect 52092 73788 52144 73840
rect 24216 73720 24268 73772
rect 78496 73720 78548 73772
rect 44088 73584 44140 73636
rect 76840 73627 76892 73636
rect 76840 73593 76849 73627
rect 76849 73593 76883 73627
rect 76883 73593 76892 73627
rect 76840 73584 76892 73593
rect 76932 73559 76984 73568
rect 76932 73525 76941 73559
rect 76941 73525 76975 73559
rect 76975 73525 76984 73559
rect 76932 73516 76984 73525
rect 19606 73414 19658 73466
rect 19670 73414 19722 73466
rect 19734 73414 19786 73466
rect 19798 73414 19850 73466
rect 50326 73414 50378 73466
rect 50390 73414 50442 73466
rect 50454 73414 50506 73466
rect 50518 73414 50570 73466
rect 81046 73414 81098 73466
rect 81110 73414 81162 73466
rect 81174 73414 81226 73466
rect 81238 73414 81290 73466
rect 39948 73244 40000 73296
rect 76564 73244 76616 73296
rect 27896 73176 27948 73228
rect 70216 73176 70268 73228
rect 43812 73108 43864 73160
rect 48780 73108 48832 73160
rect 4246 72870 4298 72922
rect 4310 72870 4362 72922
rect 4374 72870 4426 72922
rect 4438 72870 4490 72922
rect 34966 72870 35018 72922
rect 35030 72870 35082 72922
rect 35094 72870 35146 72922
rect 35158 72870 35210 72922
rect 65686 72870 65738 72922
rect 65750 72870 65802 72922
rect 65814 72870 65866 72922
rect 65878 72870 65930 72922
rect 96406 72870 96458 72922
rect 96470 72870 96522 72922
rect 96534 72870 96586 72922
rect 96598 72870 96650 72922
rect 13728 72632 13780 72684
rect 84200 72768 84252 72820
rect 84568 72768 84620 72820
rect 13544 72607 13596 72616
rect 13544 72573 13553 72607
rect 13553 72573 13587 72607
rect 13587 72573 13596 72607
rect 13544 72564 13596 72573
rect 78588 72564 78640 72616
rect 50068 72496 50120 72548
rect 50620 72496 50672 72548
rect 59912 72496 59964 72548
rect 82912 72496 82964 72548
rect 13636 72428 13688 72480
rect 74540 72428 74592 72480
rect 79968 72428 80020 72480
rect 19606 72326 19658 72378
rect 19670 72326 19722 72378
rect 19734 72326 19786 72378
rect 19798 72326 19850 72378
rect 50326 72326 50378 72378
rect 50390 72326 50442 72378
rect 50454 72326 50506 72378
rect 50518 72326 50570 72378
rect 81046 72326 81098 72378
rect 81110 72326 81162 72378
rect 81174 72326 81226 72378
rect 81238 72326 81290 72378
rect 1952 72224 2004 72276
rect 9496 72088 9548 72140
rect 50712 72224 50764 72276
rect 48780 72156 48832 72208
rect 30840 72020 30892 72072
rect 23204 71952 23256 72004
rect 9680 71927 9732 71936
rect 9680 71893 9689 71927
rect 9689 71893 9723 71927
rect 9723 71893 9732 71927
rect 9680 71884 9732 71893
rect 25320 71884 25372 71936
rect 54852 71927 54904 71936
rect 54852 71893 54861 71927
rect 54861 71893 54895 71927
rect 54895 71893 54904 71927
rect 54852 71884 54904 71893
rect 55312 72131 55364 72140
rect 55312 72097 55321 72131
rect 55321 72097 55355 72131
rect 55355 72097 55364 72131
rect 60004 72156 60056 72208
rect 55312 72088 55364 72097
rect 59912 72131 59964 72140
rect 59912 72097 59922 72131
rect 59922 72097 59956 72131
rect 59956 72097 59964 72131
rect 60096 72131 60148 72140
rect 59912 72088 59964 72097
rect 60096 72097 60105 72131
rect 60105 72097 60139 72131
rect 60139 72097 60148 72131
rect 60096 72088 60148 72097
rect 79968 72224 80020 72276
rect 78680 72088 78732 72140
rect 78864 72063 78916 72072
rect 78864 72029 78873 72063
rect 78873 72029 78907 72063
rect 78907 72029 78916 72063
rect 78864 72020 78916 72029
rect 55220 71952 55272 72004
rect 59544 71952 59596 72004
rect 63224 71952 63276 72004
rect 78588 71884 78640 71936
rect 78680 71927 78732 71936
rect 78680 71893 78689 71927
rect 78689 71893 78723 71927
rect 78723 71893 78732 71927
rect 80244 71927 80296 71936
rect 78680 71884 78732 71893
rect 80244 71893 80253 71927
rect 80253 71893 80287 71927
rect 80287 71893 80296 71927
rect 93676 71952 93728 72004
rect 89260 71927 89312 71936
rect 80244 71884 80296 71893
rect 89260 71893 89269 71927
rect 89269 71893 89303 71927
rect 89303 71893 89312 71927
rect 89260 71884 89312 71893
rect 4246 71782 4298 71834
rect 4310 71782 4362 71834
rect 4374 71782 4426 71834
rect 4438 71782 4490 71834
rect 34966 71782 35018 71834
rect 35030 71782 35082 71834
rect 35094 71782 35146 71834
rect 35158 71782 35210 71834
rect 65686 71782 65738 71834
rect 65750 71782 65802 71834
rect 65814 71782 65866 71834
rect 65878 71782 65930 71834
rect 96406 71782 96458 71834
rect 96470 71782 96522 71834
rect 96534 71782 96586 71834
rect 96598 71782 96650 71834
rect 71228 71655 71280 71664
rect 71228 71621 71237 71655
rect 71237 71621 71271 71655
rect 71271 71621 71280 71655
rect 71228 71612 71280 71621
rect 66168 71544 66220 71596
rect 85672 71544 85724 71596
rect 27160 71476 27212 71528
rect 65432 71476 65484 71528
rect 66628 71476 66680 71528
rect 70676 71519 70728 71528
rect 70676 71485 70685 71519
rect 70685 71485 70719 71519
rect 70719 71485 70728 71519
rect 70676 71476 70728 71485
rect 70860 71519 70912 71528
rect 70860 71485 70869 71519
rect 70869 71485 70903 71519
rect 70903 71485 70912 71519
rect 70860 71476 70912 71485
rect 71136 71519 71188 71528
rect 71136 71485 71139 71519
rect 71139 71485 71188 71519
rect 71136 71476 71188 71485
rect 24032 71340 24084 71392
rect 26976 71340 27028 71392
rect 70124 71408 70176 71460
rect 70952 71451 71004 71460
rect 70952 71417 70961 71451
rect 70961 71417 70995 71451
rect 70995 71417 71004 71451
rect 70952 71408 71004 71417
rect 75184 71408 75236 71460
rect 65432 71340 65484 71392
rect 19606 71238 19658 71290
rect 19670 71238 19722 71290
rect 19734 71238 19786 71290
rect 19798 71238 19850 71290
rect 50326 71238 50378 71290
rect 50390 71238 50442 71290
rect 50454 71238 50506 71290
rect 50518 71238 50570 71290
rect 81046 71238 81098 71290
rect 81110 71238 81162 71290
rect 81174 71238 81226 71290
rect 81238 71238 81290 71290
rect 16212 71136 16264 71188
rect 26424 71136 26476 71188
rect 26976 71136 27028 71188
rect 2136 71068 2188 71120
rect 24032 71068 24084 71120
rect 26792 71111 26844 71120
rect 26792 71077 26801 71111
rect 26801 71077 26835 71111
rect 26835 71077 26844 71111
rect 26792 71068 26844 71077
rect 36360 71068 36412 71120
rect 53288 71068 53340 71120
rect 63592 71068 63644 71120
rect 26332 71000 26384 71052
rect 26700 71043 26752 71052
rect 26700 71009 26709 71043
rect 26709 71009 26743 71043
rect 26743 71009 26752 71043
rect 26700 71000 26752 71009
rect 25688 70839 25740 70848
rect 25688 70805 25697 70839
rect 25697 70805 25731 70839
rect 25731 70805 25740 70839
rect 25688 70796 25740 70805
rect 26792 70932 26844 70984
rect 53380 71000 53432 71052
rect 68100 71000 68152 71052
rect 27160 70932 27212 70984
rect 95608 70932 95660 70984
rect 27068 70907 27120 70916
rect 27068 70873 27077 70907
rect 27077 70873 27111 70907
rect 27111 70873 27120 70907
rect 27068 70864 27120 70873
rect 94780 70864 94832 70916
rect 83464 70796 83516 70848
rect 4246 70694 4298 70746
rect 4310 70694 4362 70746
rect 4374 70694 4426 70746
rect 4438 70694 4490 70746
rect 34966 70694 35018 70746
rect 35030 70694 35082 70746
rect 35094 70694 35146 70746
rect 35158 70694 35210 70746
rect 65686 70694 65738 70746
rect 65750 70694 65802 70746
rect 65814 70694 65866 70746
rect 65878 70694 65930 70746
rect 96406 70694 96458 70746
rect 96470 70694 96522 70746
rect 96534 70694 96586 70746
rect 96598 70694 96650 70746
rect 25688 70592 25740 70644
rect 70032 70592 70084 70644
rect 64236 70456 64288 70508
rect 84568 70456 84620 70508
rect 57244 70388 57296 70440
rect 60004 70388 60056 70440
rect 85212 70388 85264 70440
rect 55220 70320 55272 70372
rect 77300 70320 77352 70372
rect 85580 70295 85632 70304
rect 85580 70261 85589 70295
rect 85589 70261 85623 70295
rect 85623 70261 85632 70295
rect 85580 70252 85632 70261
rect 19606 70150 19658 70202
rect 19670 70150 19722 70202
rect 19734 70150 19786 70202
rect 19798 70150 19850 70202
rect 50326 70150 50378 70202
rect 50390 70150 50442 70202
rect 50454 70150 50506 70202
rect 50518 70150 50570 70202
rect 81046 70150 81098 70202
rect 81110 70150 81162 70202
rect 81174 70150 81226 70202
rect 81238 70150 81290 70202
rect 43536 69912 43588 69964
rect 50160 69912 50212 69964
rect 78680 69912 78732 69964
rect 11336 69844 11388 69896
rect 55220 69844 55272 69896
rect 61568 69844 61620 69896
rect 93032 69844 93084 69896
rect 15936 69819 15988 69828
rect 15936 69785 15945 69819
rect 15945 69785 15979 69819
rect 15979 69785 15988 69819
rect 15936 69776 15988 69785
rect 37924 69776 37976 69828
rect 89260 69776 89312 69828
rect 23664 69708 23716 69760
rect 77208 69708 77260 69760
rect 4246 69606 4298 69658
rect 4310 69606 4362 69658
rect 4374 69606 4426 69658
rect 4438 69606 4490 69658
rect 34966 69606 35018 69658
rect 35030 69606 35082 69658
rect 35094 69606 35146 69658
rect 35158 69606 35210 69658
rect 65686 69606 65738 69658
rect 65750 69606 65802 69658
rect 65814 69606 65866 69658
rect 65878 69606 65930 69658
rect 96406 69606 96458 69658
rect 96470 69606 96522 69658
rect 96534 69606 96586 69658
rect 96598 69606 96650 69658
rect 5080 69436 5132 69488
rect 26792 69300 26844 69352
rect 28264 69300 28316 69352
rect 33876 69300 33928 69352
rect 5264 69232 5316 69284
rect 47584 69164 47636 69216
rect 88708 69164 88760 69216
rect 19606 69062 19658 69114
rect 19670 69062 19722 69114
rect 19734 69062 19786 69114
rect 19798 69062 19850 69114
rect 50326 69062 50378 69114
rect 50390 69062 50442 69114
rect 50454 69062 50506 69114
rect 50518 69062 50570 69114
rect 81046 69062 81098 69114
rect 81110 69062 81162 69114
rect 81174 69062 81226 69114
rect 81238 69062 81290 69114
rect 5356 68960 5408 69012
rect 15936 68867 15988 68876
rect 15936 68833 15945 68867
rect 15945 68833 15979 68867
rect 15979 68833 15988 68867
rect 15936 68824 15988 68833
rect 61384 68824 61436 68876
rect 78312 68960 78364 69012
rect 85856 68960 85908 69012
rect 92388 68960 92440 69012
rect 16488 68799 16540 68808
rect 16488 68765 16497 68799
rect 16497 68765 16531 68799
rect 16531 68765 16540 68799
rect 16488 68756 16540 68765
rect 61936 68799 61988 68808
rect 61936 68765 61945 68799
rect 61945 68765 61979 68799
rect 61979 68765 61988 68799
rect 61936 68756 61988 68765
rect 62396 68756 62448 68808
rect 78220 68824 78272 68876
rect 78496 68824 78548 68876
rect 83556 68824 83608 68876
rect 92388 68824 92440 68876
rect 78312 68799 78364 68808
rect 78312 68765 78321 68799
rect 78321 68765 78355 68799
rect 78355 68765 78364 68799
rect 78312 68756 78364 68765
rect 80796 68756 80848 68808
rect 84568 68799 84620 68808
rect 84568 68765 84577 68799
rect 84577 68765 84611 68799
rect 84611 68765 84620 68799
rect 84568 68756 84620 68765
rect 84844 68799 84896 68808
rect 84844 68765 84853 68799
rect 84853 68765 84887 68799
rect 84887 68765 84896 68799
rect 84844 68756 84896 68765
rect 78772 68731 78824 68740
rect 78772 68697 78781 68731
rect 78781 68697 78815 68731
rect 78815 68697 78824 68731
rect 78772 68688 78824 68697
rect 63684 68620 63736 68672
rect 90180 68663 90232 68672
rect 90180 68629 90189 68663
rect 90189 68629 90223 68663
rect 90223 68629 90232 68663
rect 90180 68620 90232 68629
rect 4246 68518 4298 68570
rect 4310 68518 4362 68570
rect 4374 68518 4426 68570
rect 4438 68518 4490 68570
rect 34966 68518 35018 68570
rect 35030 68518 35082 68570
rect 35094 68518 35146 68570
rect 35158 68518 35210 68570
rect 65686 68518 65738 68570
rect 65750 68518 65802 68570
rect 65814 68518 65866 68570
rect 65878 68518 65930 68570
rect 96406 68518 96458 68570
rect 96470 68518 96522 68570
rect 96534 68518 96586 68570
rect 96598 68518 96650 68570
rect 46204 68416 46256 68468
rect 45560 68348 45612 68400
rect 91192 68416 91244 68468
rect 10048 68323 10100 68332
rect 10048 68289 10057 68323
rect 10057 68289 10091 68323
rect 10091 68289 10100 68323
rect 10048 68280 10100 68289
rect 7012 68255 7064 68264
rect 7012 68221 7021 68255
rect 7021 68221 7055 68255
rect 7055 68221 7064 68255
rect 7012 68212 7064 68221
rect 9772 68255 9824 68264
rect 9772 68221 9781 68255
rect 9781 68221 9815 68255
rect 9815 68221 9824 68255
rect 9772 68212 9824 68221
rect 15936 68280 15988 68332
rect 31392 68280 31444 68332
rect 10692 68255 10744 68264
rect 10692 68221 10701 68255
rect 10701 68221 10735 68255
rect 10735 68221 10744 68255
rect 10692 68212 10744 68221
rect 26884 68212 26936 68264
rect 46388 68280 46440 68332
rect 90088 68348 90140 68400
rect 91836 68348 91888 68400
rect 80704 68280 80756 68332
rect 91928 68280 91980 68332
rect 92112 68280 92164 68332
rect 46848 68255 46900 68264
rect 46848 68221 46857 68255
rect 46857 68221 46891 68255
rect 46891 68221 46900 68255
rect 46848 68212 46900 68221
rect 91744 68212 91796 68264
rect 16120 68144 16172 68196
rect 39764 68076 39816 68128
rect 46204 68076 46256 68128
rect 75460 68144 75512 68196
rect 84844 68076 84896 68128
rect 19606 67974 19658 68026
rect 19670 67974 19722 68026
rect 19734 67974 19786 68026
rect 19798 67974 19850 68026
rect 50326 67974 50378 68026
rect 50390 67974 50442 68026
rect 50454 67974 50506 68026
rect 50518 67974 50570 68026
rect 81046 67974 81098 68026
rect 81110 67974 81162 68026
rect 81174 67974 81226 68026
rect 81238 67974 81290 68026
rect 16120 67779 16172 67788
rect 16120 67745 16129 67779
rect 16129 67745 16163 67779
rect 16163 67745 16172 67779
rect 16120 67736 16172 67745
rect 4712 67668 4764 67720
rect 5172 67668 5224 67720
rect 16948 67711 17000 67720
rect 16948 67677 16957 67711
rect 16957 67677 16991 67711
rect 16991 67677 17000 67711
rect 16948 67668 17000 67677
rect 73528 67600 73580 67652
rect 74080 67600 74132 67652
rect 90916 67643 90968 67652
rect 90916 67609 90925 67643
rect 90925 67609 90959 67643
rect 90959 67609 90968 67643
rect 90916 67600 90968 67609
rect 4988 67532 5040 67584
rect 5264 67532 5316 67584
rect 23480 67532 23532 67584
rect 23756 67532 23808 67584
rect 29276 67532 29328 67584
rect 29920 67532 29972 67584
rect 4246 67430 4298 67482
rect 4310 67430 4362 67482
rect 4374 67430 4426 67482
rect 4438 67430 4490 67482
rect 34966 67430 35018 67482
rect 35030 67430 35082 67482
rect 35094 67430 35146 67482
rect 35158 67430 35210 67482
rect 65686 67430 65738 67482
rect 65750 67430 65802 67482
rect 65814 67430 65866 67482
rect 65878 67430 65930 67482
rect 96406 67430 96458 67482
rect 96470 67430 96522 67482
rect 96534 67430 96586 67482
rect 96598 67430 96650 67482
rect 4068 67328 4120 67380
rect 73896 67328 73948 67380
rect 4252 67260 4304 67312
rect 4712 67260 4764 67312
rect 4160 67235 4212 67244
rect 4160 67201 4194 67235
rect 4194 67201 4212 67235
rect 4160 67192 4212 67201
rect 5172 67192 5224 67244
rect 13636 67192 13688 67244
rect 3976 67124 4028 67176
rect 4068 67167 4120 67176
rect 4068 67133 4077 67167
rect 4077 67133 4111 67167
rect 4111 67133 4120 67167
rect 4068 67124 4120 67133
rect 4436 67167 4488 67176
rect 4436 67133 4441 67167
rect 4441 67133 4475 67167
rect 4475 67133 4488 67167
rect 4160 67056 4212 67108
rect 4436 67124 4488 67133
rect 4528 67124 4580 67176
rect 19432 67192 19484 67244
rect 20628 67235 20680 67244
rect 20628 67201 20637 67235
rect 20637 67201 20671 67235
rect 20671 67201 20680 67235
rect 20628 67192 20680 67201
rect 30840 67260 30892 67312
rect 33968 67260 34020 67312
rect 89168 67260 89220 67312
rect 35256 67192 35308 67244
rect 76840 67192 76892 67244
rect 20260 67167 20312 67176
rect 4344 67056 4396 67108
rect 13544 67056 13596 67108
rect 10508 66988 10560 67040
rect 20260 67133 20269 67167
rect 20269 67133 20303 67167
rect 20303 67133 20312 67167
rect 20260 67124 20312 67133
rect 20444 67167 20496 67176
rect 20444 67133 20453 67167
rect 20453 67133 20487 67167
rect 20487 67133 20496 67167
rect 20444 67124 20496 67133
rect 27528 67124 27580 67176
rect 52368 67167 52420 67176
rect 52368 67133 52377 67167
rect 52377 67133 52411 67167
rect 52411 67133 52420 67167
rect 52368 67124 52420 67133
rect 63592 67124 63644 67176
rect 72700 67167 72752 67176
rect 72700 67133 72709 67167
rect 72709 67133 72743 67167
rect 72743 67133 72752 67167
rect 72700 67124 72752 67133
rect 29276 67056 29328 67108
rect 52644 67099 52696 67108
rect 52644 67065 52653 67099
rect 52653 67065 52687 67099
rect 52687 67065 52696 67099
rect 52644 67056 52696 67065
rect 70216 67056 70268 67108
rect 76196 67056 76248 67108
rect 76656 67056 76708 67108
rect 86592 67056 86644 67108
rect 20076 66988 20128 67040
rect 52552 67031 52604 67040
rect 52552 66997 52561 67031
rect 52561 66997 52595 67031
rect 52595 66997 52604 67031
rect 52552 66988 52604 66997
rect 56968 66988 57020 67040
rect 57888 66988 57940 67040
rect 79324 66988 79376 67040
rect 79600 66988 79652 67040
rect 19606 66886 19658 66938
rect 19670 66886 19722 66938
rect 19734 66886 19786 66938
rect 19798 66886 19850 66938
rect 50326 66886 50378 66938
rect 50390 66886 50442 66938
rect 50454 66886 50506 66938
rect 50518 66886 50570 66938
rect 81046 66886 81098 66938
rect 81110 66886 81162 66938
rect 81174 66886 81226 66938
rect 81238 66886 81290 66938
rect 27252 66784 27304 66836
rect 27528 66784 27580 66836
rect 34152 66827 34204 66836
rect 34152 66793 34161 66827
rect 34161 66793 34195 66827
rect 34195 66793 34204 66827
rect 34152 66784 34204 66793
rect 63592 66784 63644 66836
rect 89444 66784 89496 66836
rect 23756 66648 23808 66700
rect 6368 66580 6420 66632
rect 17684 66512 17736 66564
rect 9404 66444 9456 66496
rect 13728 66444 13780 66496
rect 46940 66580 46992 66632
rect 53288 66444 53340 66496
rect 77944 66487 77996 66496
rect 77944 66453 77953 66487
rect 77953 66453 77987 66487
rect 77987 66453 77996 66487
rect 77944 66444 77996 66453
rect 4246 66342 4298 66394
rect 4310 66342 4362 66394
rect 4374 66342 4426 66394
rect 4438 66342 4490 66394
rect 34966 66342 35018 66394
rect 35030 66342 35082 66394
rect 35094 66342 35146 66394
rect 35158 66342 35210 66394
rect 65686 66342 65738 66394
rect 65750 66342 65802 66394
rect 65814 66342 65866 66394
rect 65878 66342 65930 66394
rect 96406 66342 96458 66394
rect 96470 66342 96522 66394
rect 96534 66342 96586 66394
rect 96598 66342 96650 66394
rect 49516 66036 49568 66088
rect 49884 66036 49936 66088
rect 78864 66036 78916 66088
rect 80520 66079 80572 66088
rect 80520 66045 80529 66079
rect 80529 66045 80563 66079
rect 80563 66045 80572 66079
rect 80520 66036 80572 66045
rect 81992 66036 82044 66088
rect 82544 66079 82596 66088
rect 82544 66045 82553 66079
rect 82553 66045 82587 66079
rect 82587 66045 82596 66079
rect 82544 66036 82596 66045
rect 91192 66104 91244 66156
rect 83096 66079 83148 66088
rect 83096 66045 83105 66079
rect 83105 66045 83139 66079
rect 83139 66045 83148 66079
rect 83096 66036 83148 66045
rect 83280 66079 83332 66088
rect 83280 66045 83289 66079
rect 83289 66045 83323 66079
rect 83323 66045 83332 66079
rect 83280 66036 83332 66045
rect 77300 65900 77352 65952
rect 83556 65943 83608 65952
rect 83556 65909 83565 65943
rect 83565 65909 83599 65943
rect 83599 65909 83608 65943
rect 83556 65900 83608 65909
rect 19606 65798 19658 65850
rect 19670 65798 19722 65850
rect 19734 65798 19786 65850
rect 19798 65798 19850 65850
rect 50326 65798 50378 65850
rect 50390 65798 50442 65850
rect 50454 65798 50506 65850
rect 50518 65798 50570 65850
rect 81046 65798 81098 65850
rect 81110 65798 81162 65850
rect 81174 65798 81226 65850
rect 81238 65798 81290 65850
rect 36544 65696 36596 65748
rect 83556 65696 83608 65748
rect 2320 65628 2372 65680
rect 27344 65628 27396 65680
rect 38200 65628 38252 65680
rect 46756 65628 46808 65680
rect 7380 65603 7432 65612
rect 7380 65569 7389 65603
rect 7389 65569 7423 65603
rect 7423 65569 7432 65603
rect 7380 65560 7432 65569
rect 21456 65560 21508 65612
rect 52552 65560 52604 65612
rect 53564 65560 53616 65612
rect 75000 65560 75052 65612
rect 25964 65492 26016 65544
rect 33784 65492 33836 65544
rect 35440 65492 35492 65544
rect 72700 65492 72752 65544
rect 84568 65424 84620 65476
rect 85396 65424 85448 65476
rect 44272 65356 44324 65408
rect 45468 65356 45520 65408
rect 4246 65254 4298 65306
rect 4310 65254 4362 65306
rect 4374 65254 4426 65306
rect 4438 65254 4490 65306
rect 34966 65254 35018 65306
rect 35030 65254 35082 65306
rect 35094 65254 35146 65306
rect 35158 65254 35210 65306
rect 65686 65254 65738 65306
rect 65750 65254 65802 65306
rect 65814 65254 65866 65306
rect 65878 65254 65930 65306
rect 96406 65254 96458 65306
rect 96470 65254 96522 65306
rect 96534 65254 96586 65306
rect 96598 65254 96650 65306
rect 46756 65016 46808 65068
rect 80336 65152 80388 65204
rect 90548 65195 90600 65204
rect 90548 65161 90557 65195
rect 90557 65161 90591 65195
rect 90591 65161 90600 65195
rect 90548 65152 90600 65161
rect 91192 65152 91244 65204
rect 27344 64948 27396 65000
rect 58900 64948 58952 65000
rect 59452 64991 59504 65000
rect 59452 64957 59461 64991
rect 59461 64957 59495 64991
rect 59495 64957 59504 64991
rect 59452 64948 59504 64957
rect 60280 65016 60332 65068
rect 88340 65084 88392 65136
rect 80888 65016 80940 65068
rect 60188 64991 60240 65000
rect 9772 64880 9824 64932
rect 11888 64880 11940 64932
rect 28632 64923 28684 64932
rect 28632 64889 28641 64923
rect 28641 64889 28675 64923
rect 28675 64889 28684 64923
rect 28632 64880 28684 64889
rect 45468 64880 45520 64932
rect 60188 64957 60197 64991
rect 60197 64957 60231 64991
rect 60231 64957 60240 64991
rect 60188 64948 60240 64957
rect 60556 64880 60608 64932
rect 85396 64880 85448 64932
rect 86960 64880 87012 64932
rect 91192 64880 91244 64932
rect 39672 64812 39724 64864
rect 81716 64812 81768 64864
rect 19606 64710 19658 64762
rect 19670 64710 19722 64762
rect 19734 64710 19786 64762
rect 19798 64710 19850 64762
rect 50326 64710 50378 64762
rect 50390 64710 50442 64762
rect 50454 64710 50506 64762
rect 50518 64710 50570 64762
rect 81046 64710 81098 64762
rect 81110 64710 81162 64762
rect 81174 64710 81226 64762
rect 81238 64710 81290 64762
rect 27344 64651 27396 64660
rect 27344 64617 27353 64651
rect 27353 64617 27387 64651
rect 27387 64617 27396 64651
rect 27344 64608 27396 64617
rect 49700 64608 49752 64660
rect 50988 64608 51040 64660
rect 16028 64472 16080 64524
rect 49424 64515 49476 64524
rect 49424 64481 49433 64515
rect 49433 64481 49467 64515
rect 49467 64481 49476 64515
rect 49424 64472 49476 64481
rect 50068 64540 50120 64592
rect 50344 64540 50396 64592
rect 80244 64540 80296 64592
rect 49516 64404 49568 64456
rect 55312 64472 55364 64524
rect 56048 64472 56100 64524
rect 91744 64515 91796 64524
rect 91744 64481 91753 64515
rect 91753 64481 91787 64515
rect 91787 64481 91796 64515
rect 91744 64472 91796 64481
rect 91836 64515 91888 64524
rect 91836 64481 91845 64515
rect 91845 64481 91879 64515
rect 91879 64481 91888 64515
rect 91836 64472 91888 64481
rect 95056 64515 95108 64524
rect 95056 64481 95065 64515
rect 95065 64481 95099 64515
rect 95099 64481 95108 64515
rect 95056 64472 95108 64481
rect 95792 64515 95844 64524
rect 95792 64481 95801 64515
rect 95801 64481 95835 64515
rect 95835 64481 95844 64515
rect 95792 64472 95844 64481
rect 29552 64336 29604 64388
rect 49884 64336 49936 64388
rect 26424 64311 26476 64320
rect 26424 64277 26433 64311
rect 26433 64277 26467 64311
rect 26467 64277 26476 64311
rect 26424 64268 26476 64277
rect 49976 64268 50028 64320
rect 75368 64404 75420 64456
rect 75828 64404 75880 64456
rect 87696 64404 87748 64456
rect 95240 64447 95292 64456
rect 95240 64413 95249 64447
rect 95249 64413 95283 64447
rect 95283 64413 95292 64447
rect 95240 64404 95292 64413
rect 50252 64336 50304 64388
rect 50160 64268 50212 64320
rect 50896 64268 50948 64320
rect 51448 64268 51500 64320
rect 67088 64268 67140 64320
rect 92756 64336 92808 64388
rect 4246 64166 4298 64218
rect 4310 64166 4362 64218
rect 4374 64166 4426 64218
rect 4438 64166 4490 64218
rect 34966 64166 35018 64218
rect 35030 64166 35082 64218
rect 35094 64166 35146 64218
rect 35158 64166 35210 64218
rect 65686 64166 65738 64218
rect 65750 64166 65802 64218
rect 65814 64166 65866 64218
rect 65878 64166 65930 64218
rect 96406 64166 96458 64218
rect 96470 64166 96522 64218
rect 96534 64166 96586 64218
rect 96598 64166 96650 64218
rect 8944 64107 8996 64116
rect 8300 63903 8352 63912
rect 8300 63869 8309 63903
rect 8309 63869 8343 63903
rect 8343 63869 8352 63903
rect 8300 63860 8352 63869
rect 8668 63996 8720 64048
rect 8944 64073 8953 64107
rect 8953 64073 8987 64107
rect 8987 64073 8996 64107
rect 8944 64064 8996 64073
rect 34152 64064 34204 64116
rect 14280 63996 14332 64048
rect 49424 63996 49476 64048
rect 49700 64064 49752 64116
rect 50896 64064 50948 64116
rect 61936 64064 61988 64116
rect 66352 64107 66404 64116
rect 66352 64073 66361 64107
rect 66361 64073 66395 64107
rect 66395 64073 66404 64107
rect 66352 64064 66404 64073
rect 68468 64107 68520 64116
rect 49976 63996 50028 64048
rect 52460 63996 52512 64048
rect 53012 63996 53064 64048
rect 40776 63928 40828 63980
rect 62672 63928 62724 63980
rect 54852 63860 54904 63912
rect 66996 63996 67048 64048
rect 68468 64073 68477 64107
rect 68477 64073 68511 64107
rect 68511 64073 68520 64107
rect 68468 64064 68520 64073
rect 75000 64064 75052 64116
rect 75276 63996 75328 64048
rect 82452 64039 82504 64048
rect 67272 63928 67324 63980
rect 24124 63792 24176 63844
rect 33784 63792 33836 63844
rect 49700 63792 49752 63844
rect 45376 63724 45428 63776
rect 47952 63724 48004 63776
rect 75368 63860 75420 63912
rect 82452 64005 82461 64039
rect 82461 64005 82495 64039
rect 82495 64005 82504 64039
rect 82452 63996 82504 64005
rect 67456 63724 67508 63776
rect 71688 63792 71740 63844
rect 78864 63792 78916 63844
rect 81716 63792 81768 63844
rect 92756 63792 92808 63844
rect 92940 63767 92992 63776
rect 92940 63733 92949 63767
rect 92949 63733 92983 63767
rect 92983 63733 92992 63767
rect 92940 63724 92992 63733
rect 19606 63622 19658 63674
rect 19670 63622 19722 63674
rect 19734 63622 19786 63674
rect 19798 63622 19850 63674
rect 50326 63622 50378 63674
rect 50390 63622 50442 63674
rect 50454 63622 50506 63674
rect 50518 63622 50570 63674
rect 81046 63622 81098 63674
rect 81110 63622 81162 63674
rect 81174 63622 81226 63674
rect 81238 63622 81290 63674
rect 28356 63520 28408 63572
rect 34152 63520 34204 63572
rect 45468 63520 45520 63572
rect 50988 63520 51040 63572
rect 48964 63452 49016 63504
rect 49516 63452 49568 63504
rect 8392 63384 8444 63436
rect 19340 63384 19392 63436
rect 28356 63384 28408 63436
rect 57060 63316 57112 63368
rect 57796 63316 57848 63368
rect 15476 63248 15528 63300
rect 27252 63291 27304 63300
rect 11980 63180 12032 63232
rect 18696 63180 18748 63232
rect 27252 63257 27261 63291
rect 27261 63257 27295 63291
rect 27295 63257 27304 63291
rect 27252 63248 27304 63257
rect 34244 63180 34296 63232
rect 53104 63180 53156 63232
rect 79692 63223 79744 63232
rect 79692 63189 79701 63223
rect 79701 63189 79735 63223
rect 79735 63189 79744 63223
rect 79692 63180 79744 63189
rect 4246 63078 4298 63130
rect 4310 63078 4362 63130
rect 4374 63078 4426 63130
rect 4438 63078 4490 63130
rect 34966 63078 35018 63130
rect 35030 63078 35082 63130
rect 35094 63078 35146 63130
rect 35158 63078 35210 63130
rect 65686 63078 65738 63130
rect 65750 63078 65802 63130
rect 65814 63078 65866 63130
rect 65878 63078 65930 63130
rect 96406 63078 96458 63130
rect 96470 63078 96522 63130
rect 96534 63078 96586 63130
rect 96598 63078 96650 63130
rect 14740 62908 14792 62960
rect 15660 62840 15712 62892
rect 22100 62976 22152 63028
rect 37832 62976 37884 63028
rect 20628 62908 20680 62960
rect 57336 62908 57388 62960
rect 20444 62840 20496 62892
rect 60924 62840 60976 62892
rect 33784 62815 33836 62824
rect 12992 62704 13044 62756
rect 33784 62781 33793 62815
rect 33793 62781 33827 62815
rect 33827 62781 33836 62815
rect 33784 62772 33836 62781
rect 15476 62704 15528 62756
rect 33692 62679 33744 62688
rect 33692 62645 33701 62679
rect 33701 62645 33735 62679
rect 33735 62645 33744 62679
rect 33692 62636 33744 62645
rect 34152 62815 34204 62824
rect 34152 62781 34161 62815
rect 34161 62781 34195 62815
rect 34195 62781 34204 62815
rect 34152 62772 34204 62781
rect 34520 62772 34572 62824
rect 35808 62772 35860 62824
rect 93492 62772 93544 62824
rect 34244 62704 34296 62756
rect 34152 62636 34204 62688
rect 34336 62636 34388 62688
rect 19606 62534 19658 62586
rect 19670 62534 19722 62586
rect 19734 62534 19786 62586
rect 19798 62534 19850 62586
rect 50326 62534 50378 62586
rect 50390 62534 50442 62586
rect 50454 62534 50506 62586
rect 50518 62534 50570 62586
rect 81046 62534 81098 62586
rect 81110 62534 81162 62586
rect 81174 62534 81226 62586
rect 81238 62534 81290 62586
rect 33692 62432 33744 62484
rect 34520 62432 34572 62484
rect 32404 62364 32456 62416
rect 34152 62364 34204 62416
rect 34796 62364 34848 62416
rect 53564 62364 53616 62416
rect 65708 62364 65760 62416
rect 72424 62364 72476 62416
rect 12992 62339 13044 62348
rect 12992 62305 13001 62339
rect 13001 62305 13035 62339
rect 13035 62305 13044 62339
rect 12992 62296 13044 62305
rect 13176 62339 13228 62348
rect 13176 62305 13185 62339
rect 13185 62305 13219 62339
rect 13219 62305 13228 62339
rect 13176 62296 13228 62305
rect 6460 62228 6512 62280
rect 15844 62296 15896 62348
rect 49608 62296 49660 62348
rect 65616 62296 65668 62348
rect 65800 62296 65852 62348
rect 73988 62339 74040 62348
rect 73988 62305 73997 62339
rect 73997 62305 74031 62339
rect 74031 62305 74040 62339
rect 73988 62296 74040 62305
rect 49516 62228 49568 62280
rect 65708 62228 65760 62280
rect 70308 62228 70360 62280
rect 74448 62296 74500 62348
rect 83464 62339 83516 62348
rect 83464 62305 83473 62339
rect 83473 62305 83507 62339
rect 83507 62305 83516 62339
rect 83464 62296 83516 62305
rect 74264 62271 74316 62280
rect 74264 62237 74273 62271
rect 74273 62237 74307 62271
rect 74307 62237 74316 62271
rect 74264 62228 74316 62237
rect 39948 62160 40000 62212
rect 15108 62092 15160 62144
rect 36636 62092 36688 62144
rect 45468 62092 45520 62144
rect 72424 62092 72476 62144
rect 4246 61990 4298 62042
rect 4310 61990 4362 62042
rect 4374 61990 4426 62042
rect 4438 61990 4490 62042
rect 34966 61990 35018 62042
rect 35030 61990 35082 62042
rect 35094 61990 35146 62042
rect 35158 61990 35210 62042
rect 65686 61990 65738 62042
rect 65750 61990 65802 62042
rect 65814 61990 65866 62042
rect 65878 61990 65930 62042
rect 96406 61990 96458 62042
rect 96470 61990 96522 62042
rect 96534 61990 96586 62042
rect 96598 61990 96650 62042
rect 30656 61795 30708 61804
rect 30656 61761 30665 61795
rect 30665 61761 30699 61795
rect 30699 61761 30708 61795
rect 30656 61752 30708 61761
rect 57520 61888 57572 61940
rect 58624 61888 58676 61940
rect 75000 61931 75052 61940
rect 75000 61897 75009 61931
rect 75009 61897 75043 61931
rect 75043 61897 75052 61931
rect 75000 61888 75052 61897
rect 77944 61820 77996 61872
rect 30840 61727 30892 61736
rect 30840 61693 30849 61727
rect 30849 61693 30883 61727
rect 30883 61693 30892 61727
rect 30840 61684 30892 61693
rect 54208 61752 54260 61804
rect 57428 61752 57480 61804
rect 31392 61727 31444 61736
rect 31392 61693 31401 61727
rect 31401 61693 31435 61727
rect 31435 61693 31444 61727
rect 31392 61684 31444 61693
rect 48780 61727 48832 61736
rect 48780 61693 48789 61727
rect 48789 61693 48823 61727
rect 48823 61693 48832 61727
rect 48780 61684 48832 61693
rect 50988 61727 51040 61736
rect 50988 61693 50997 61727
rect 50997 61693 51031 61727
rect 51031 61693 51040 61727
rect 50988 61684 51040 61693
rect 71320 61684 71372 61736
rect 90824 61684 90876 61736
rect 44548 61616 44600 61668
rect 49608 61659 49660 61668
rect 49608 61625 49617 61659
rect 49617 61625 49651 61659
rect 49651 61625 49660 61659
rect 49608 61616 49660 61625
rect 83464 61616 83516 61668
rect 84936 61616 84988 61668
rect 31668 61591 31720 61600
rect 31668 61557 31677 61591
rect 31677 61557 31711 61591
rect 31711 61557 31720 61591
rect 31668 61548 31720 61557
rect 42708 61548 42760 61600
rect 57428 61548 57480 61600
rect 61936 61548 61988 61600
rect 93400 61591 93452 61600
rect 93400 61557 93409 61591
rect 93409 61557 93443 61591
rect 93443 61557 93452 61591
rect 93400 61548 93452 61557
rect 19606 61446 19658 61498
rect 19670 61446 19722 61498
rect 19734 61446 19786 61498
rect 19798 61446 19850 61498
rect 50326 61446 50378 61498
rect 50390 61446 50442 61498
rect 50454 61446 50506 61498
rect 50518 61446 50570 61498
rect 81046 61446 81098 61498
rect 81110 61446 81162 61498
rect 81174 61446 81226 61498
rect 81238 61446 81290 61498
rect 23112 61344 23164 61396
rect 41604 61344 41656 61396
rect 42708 61344 42760 61396
rect 30840 61276 30892 61328
rect 52920 61344 52972 61396
rect 44548 61276 44600 61328
rect 73620 61344 73672 61396
rect 74816 61344 74868 61396
rect 93400 61344 93452 61396
rect 9404 61208 9456 61260
rect 10140 61208 10192 61260
rect 41144 61251 41196 61260
rect 41144 61217 41153 61251
rect 41153 61217 41187 61251
rect 41187 61217 41196 61251
rect 41144 61208 41196 61217
rect 41420 61251 41472 61260
rect 41420 61217 41429 61251
rect 41429 61217 41463 61251
rect 41463 61217 41472 61251
rect 41696 61251 41748 61260
rect 41420 61208 41472 61217
rect 41696 61217 41705 61251
rect 41705 61217 41739 61251
rect 41739 61217 41748 61251
rect 41696 61208 41748 61217
rect 14740 61140 14792 61192
rect 35440 61140 35492 61192
rect 42892 61208 42944 61260
rect 52552 61208 52604 61260
rect 52920 61208 52972 61260
rect 57428 61208 57480 61260
rect 82452 61276 82504 61328
rect 91928 61208 91980 61260
rect 41880 61140 41932 61192
rect 57934 61140 57986 61192
rect 9036 61004 9088 61056
rect 75460 61072 75512 61124
rect 76656 61072 76708 61124
rect 83740 61072 83792 61124
rect 92020 61072 92072 61124
rect 58992 61047 59044 61056
rect 58992 61013 59001 61047
rect 59001 61013 59035 61047
rect 59035 61013 59044 61047
rect 58992 61004 59044 61013
rect 79324 61004 79376 61056
rect 89076 61004 89128 61056
rect 4246 60902 4298 60954
rect 4310 60902 4362 60954
rect 4374 60902 4426 60954
rect 4438 60902 4490 60954
rect 34966 60902 35018 60954
rect 35030 60902 35082 60954
rect 35094 60902 35146 60954
rect 35158 60902 35210 60954
rect 65686 60902 65738 60954
rect 65750 60902 65802 60954
rect 65814 60902 65866 60954
rect 65878 60902 65930 60954
rect 96406 60902 96458 60954
rect 96470 60902 96522 60954
rect 96534 60902 96586 60954
rect 96598 60902 96650 60954
rect 52552 60800 52604 60852
rect 58992 60800 59044 60852
rect 68100 60843 68152 60852
rect 7380 60732 7432 60784
rect 68100 60809 68109 60843
rect 68109 60809 68143 60843
rect 68143 60809 68152 60843
rect 68100 60800 68152 60809
rect 83740 60800 83792 60852
rect 89904 60800 89956 60852
rect 90824 60800 90876 60852
rect 31760 60596 31812 60648
rect 52736 60596 52788 60648
rect 67548 60639 67600 60648
rect 67548 60605 67557 60639
rect 67557 60605 67591 60639
rect 67591 60605 67600 60639
rect 67548 60596 67600 60605
rect 67824 60639 67876 60648
rect 67824 60605 67833 60639
rect 67833 60605 67867 60639
rect 67867 60605 67876 60639
rect 67824 60596 67876 60605
rect 68008 60596 68060 60648
rect 54852 60528 54904 60580
rect 57060 60528 57112 60580
rect 80152 60664 80204 60716
rect 75920 60596 75972 60648
rect 76932 60596 76984 60648
rect 89996 60664 90048 60716
rect 83188 60639 83240 60648
rect 83188 60605 83197 60639
rect 83197 60605 83231 60639
rect 83231 60605 83240 60639
rect 83188 60596 83240 60605
rect 83372 60639 83424 60648
rect 83372 60605 83381 60639
rect 83381 60605 83415 60639
rect 83415 60605 83424 60639
rect 83372 60596 83424 60605
rect 83648 60639 83700 60648
rect 83648 60605 83657 60639
rect 83657 60605 83691 60639
rect 83691 60605 83700 60639
rect 83648 60596 83700 60605
rect 29736 60460 29788 60512
rect 80888 60528 80940 60580
rect 84844 60596 84896 60648
rect 91928 60596 91980 60648
rect 19606 60358 19658 60410
rect 19670 60358 19722 60410
rect 19734 60358 19786 60410
rect 19798 60358 19850 60410
rect 50326 60358 50378 60410
rect 50390 60358 50442 60410
rect 50454 60358 50506 60410
rect 50518 60358 50570 60410
rect 81046 60358 81098 60410
rect 81110 60358 81162 60410
rect 81174 60358 81226 60410
rect 81238 60358 81290 60410
rect 33968 60188 34020 60240
rect 35900 60188 35952 60240
rect 5080 60120 5132 60172
rect 27712 60120 27764 60172
rect 44272 60256 44324 60308
rect 54392 60256 54444 60308
rect 54760 60256 54812 60308
rect 62028 60256 62080 60308
rect 68008 60256 68060 60308
rect 75736 60256 75788 60308
rect 83648 60256 83700 60308
rect 67640 60188 67692 60240
rect 72700 60188 72752 60240
rect 84844 60188 84896 60240
rect 6000 60095 6052 60104
rect 6000 60061 6009 60095
rect 6009 60061 6043 60095
rect 6043 60061 6052 60095
rect 6000 60052 6052 60061
rect 34152 60052 34204 60104
rect 74816 60163 74868 60172
rect 74816 60129 74825 60163
rect 74825 60129 74859 60163
rect 74859 60129 74868 60163
rect 74816 60120 74868 60129
rect 80428 60120 80480 60172
rect 83372 60120 83424 60172
rect 89904 60120 89956 60172
rect 34520 59984 34572 60036
rect 35256 59984 35308 60036
rect 35900 59984 35952 60036
rect 54484 60052 54536 60104
rect 56968 60052 57020 60104
rect 89996 60095 90048 60104
rect 89996 60061 90005 60095
rect 90005 60061 90039 60095
rect 90039 60061 90048 60095
rect 89996 60052 90048 60061
rect 33784 59916 33836 59968
rect 72332 59984 72384 60036
rect 67180 59959 67232 59968
rect 67180 59925 67189 59959
rect 67189 59925 67223 59959
rect 67223 59925 67232 59959
rect 67180 59916 67232 59925
rect 4246 59814 4298 59866
rect 4310 59814 4362 59866
rect 4374 59814 4426 59866
rect 4438 59814 4490 59866
rect 34966 59814 35018 59866
rect 35030 59814 35082 59866
rect 35094 59814 35146 59866
rect 35158 59814 35210 59866
rect 65686 59814 65738 59866
rect 65750 59814 65802 59866
rect 65814 59814 65866 59866
rect 65878 59814 65930 59866
rect 96406 59814 96458 59866
rect 96470 59814 96522 59866
rect 96534 59814 96586 59866
rect 96598 59814 96650 59866
rect 29460 59712 29512 59764
rect 30288 59712 30340 59764
rect 38292 59644 38344 59696
rect 64880 59644 64932 59696
rect 65432 59644 65484 59696
rect 6460 59508 6512 59560
rect 18144 59508 18196 59560
rect 38292 59551 38344 59560
rect 38292 59517 38301 59551
rect 38301 59517 38335 59551
rect 38335 59517 38344 59551
rect 38292 59508 38344 59517
rect 54852 59576 54904 59628
rect 57152 59576 57204 59628
rect 57796 59576 57848 59628
rect 38844 59551 38896 59560
rect 18604 59372 18656 59424
rect 37740 59372 37792 59424
rect 38844 59517 38853 59551
rect 38853 59517 38887 59551
rect 38887 59517 38896 59551
rect 38844 59508 38896 59517
rect 39028 59483 39080 59492
rect 39028 59449 39037 59483
rect 39037 59449 39071 59483
rect 39071 59449 39080 59483
rect 39028 59440 39080 59449
rect 58164 59508 58216 59560
rect 58716 59508 58768 59560
rect 54484 59440 54536 59492
rect 64880 59508 64932 59560
rect 55772 59372 55824 59424
rect 63684 59372 63736 59424
rect 63960 59372 64012 59424
rect 65340 59372 65392 59424
rect 66076 59372 66128 59424
rect 19606 59270 19658 59322
rect 19670 59270 19722 59322
rect 19734 59270 19786 59322
rect 19798 59270 19850 59322
rect 50326 59270 50378 59322
rect 50390 59270 50442 59322
rect 50454 59270 50506 59322
rect 50518 59270 50570 59322
rect 81046 59270 81098 59322
rect 81110 59270 81162 59322
rect 81174 59270 81226 59322
rect 81238 59270 81290 59322
rect 34796 59168 34848 59220
rect 15660 59100 15712 59152
rect 20996 59032 21048 59084
rect 27712 58964 27764 59016
rect 28172 58964 28224 59016
rect 6552 58896 6604 58948
rect 37740 59032 37792 59084
rect 39028 59168 39080 59220
rect 93676 59168 93728 59220
rect 58900 59100 58952 59152
rect 80152 59100 80204 59152
rect 43076 59032 43128 59084
rect 53564 59032 53616 59084
rect 76564 59032 76616 59084
rect 15476 58828 15528 58880
rect 86868 58964 86920 59016
rect 93676 59007 93728 59016
rect 93676 58973 93685 59007
rect 93685 58973 93719 59007
rect 93719 58973 93728 59007
rect 93676 58964 93728 58973
rect 51448 58896 51500 58948
rect 78588 58896 78640 58948
rect 83924 58828 83976 58880
rect 4246 58726 4298 58778
rect 4310 58726 4362 58778
rect 4374 58726 4426 58778
rect 4438 58726 4490 58778
rect 34966 58726 35018 58778
rect 35030 58726 35082 58778
rect 35094 58726 35146 58778
rect 35158 58726 35210 58778
rect 65686 58726 65738 58778
rect 65750 58726 65802 58778
rect 65814 58726 65866 58778
rect 65878 58726 65930 58778
rect 96406 58726 96458 58778
rect 96470 58726 96522 58778
rect 96534 58726 96586 58778
rect 96598 58726 96650 58778
rect 19340 58624 19392 58676
rect 86224 58624 86276 58676
rect 57060 58488 57112 58540
rect 57428 58488 57480 58540
rect 58164 58420 58216 58472
rect 58624 58420 58676 58472
rect 81348 58284 81400 58336
rect 19606 58182 19658 58234
rect 19670 58182 19722 58234
rect 19734 58182 19786 58234
rect 19798 58182 19850 58234
rect 50326 58182 50378 58234
rect 50390 58182 50442 58234
rect 50454 58182 50506 58234
rect 50518 58182 50570 58234
rect 81046 58182 81098 58234
rect 81110 58182 81162 58234
rect 81174 58182 81226 58234
rect 81238 58182 81290 58234
rect 55864 57876 55916 57928
rect 56508 57876 56560 57928
rect 93676 57740 93728 57792
rect 4246 57638 4298 57690
rect 4310 57638 4362 57690
rect 4374 57638 4426 57690
rect 4438 57638 4490 57690
rect 34966 57638 35018 57690
rect 35030 57638 35082 57690
rect 35094 57638 35146 57690
rect 35158 57638 35210 57690
rect 65686 57638 65738 57690
rect 65750 57638 65802 57690
rect 65814 57638 65866 57690
rect 65878 57638 65930 57690
rect 96406 57638 96458 57690
rect 96470 57638 96522 57690
rect 96534 57638 96586 57690
rect 96598 57638 96650 57690
rect 9220 57536 9272 57588
rect 18788 57468 18840 57520
rect 64052 57468 64104 57520
rect 5356 57400 5408 57452
rect 22744 57400 22796 57452
rect 37556 57400 37608 57452
rect 85948 57400 86000 57452
rect 86868 57400 86920 57452
rect 7196 57332 7248 57384
rect 14004 57375 14056 57384
rect 14004 57341 14013 57375
rect 14013 57341 14047 57375
rect 14047 57341 14056 57375
rect 14004 57332 14056 57341
rect 46940 57332 46992 57384
rect 8484 57264 8536 57316
rect 15016 57264 15068 57316
rect 51908 57264 51960 57316
rect 10692 57239 10744 57248
rect 10692 57205 10701 57239
rect 10701 57205 10735 57239
rect 10735 57205 10744 57239
rect 10692 57196 10744 57205
rect 56508 57264 56560 57316
rect 64512 57264 64564 57316
rect 82360 57239 82412 57248
rect 82360 57205 82369 57239
rect 82369 57205 82403 57239
rect 82403 57205 82412 57239
rect 94320 57332 94372 57384
rect 82360 57196 82412 57205
rect 19606 57094 19658 57146
rect 19670 57094 19722 57146
rect 19734 57094 19786 57146
rect 19798 57094 19850 57146
rect 50326 57094 50378 57146
rect 50390 57094 50442 57146
rect 50454 57094 50506 57146
rect 50518 57094 50570 57146
rect 81046 57094 81098 57146
rect 81110 57094 81162 57146
rect 81174 57094 81226 57146
rect 81238 57094 81290 57146
rect 10692 56992 10744 57044
rect 35440 56992 35492 57044
rect 59268 56992 59320 57044
rect 64052 56967 64104 56976
rect 64052 56933 64061 56967
rect 64061 56933 64095 56967
rect 64095 56933 64104 56967
rect 64512 56967 64564 56976
rect 64052 56924 64104 56933
rect 37464 56899 37516 56908
rect 37464 56865 37473 56899
rect 37473 56865 37507 56899
rect 37507 56865 37516 56899
rect 37464 56856 37516 56865
rect 60648 56856 60700 56908
rect 64512 56933 64521 56967
rect 64521 56933 64555 56967
rect 64555 56933 64564 56967
rect 64512 56924 64564 56933
rect 94044 56924 94096 56976
rect 64604 56899 64656 56908
rect 64604 56865 64613 56899
rect 64613 56865 64647 56899
rect 64647 56865 64656 56899
rect 64604 56856 64656 56865
rect 68744 56899 68796 56908
rect 68744 56865 68753 56899
rect 68753 56865 68787 56899
rect 68787 56865 68796 56899
rect 68744 56856 68796 56865
rect 50436 56788 50488 56840
rect 53748 56788 53800 56840
rect 96068 56856 96120 56908
rect 97172 56899 97224 56908
rect 97172 56865 97181 56899
rect 97181 56865 97215 56899
rect 97215 56865 97224 56899
rect 97172 56856 97224 56865
rect 45560 56720 45612 56772
rect 46848 56720 46900 56772
rect 94964 56652 95016 56704
rect 4246 56550 4298 56602
rect 4310 56550 4362 56602
rect 4374 56550 4426 56602
rect 4438 56550 4490 56602
rect 34966 56550 35018 56602
rect 35030 56550 35082 56602
rect 35094 56550 35146 56602
rect 35158 56550 35210 56602
rect 65686 56550 65738 56602
rect 65750 56550 65802 56602
rect 65814 56550 65866 56602
rect 65878 56550 65930 56602
rect 96406 56550 96458 56602
rect 96470 56550 96522 56602
rect 96534 56550 96586 56602
rect 96598 56550 96650 56602
rect 31760 56448 31812 56500
rect 96252 56448 96304 56500
rect 45744 56380 45796 56432
rect 47584 56380 47636 56432
rect 9496 56244 9548 56296
rect 26332 56176 26384 56228
rect 27160 56244 27212 56296
rect 33968 56287 34020 56296
rect 33968 56253 33977 56287
rect 33977 56253 34011 56287
rect 34011 56253 34020 56287
rect 33968 56244 34020 56253
rect 26608 56176 26660 56228
rect 37464 56312 37516 56364
rect 38108 56312 38160 56364
rect 69848 56312 69900 56364
rect 49976 56244 50028 56296
rect 50436 56287 50488 56296
rect 50436 56253 50445 56287
rect 50445 56253 50479 56287
rect 50479 56253 50488 56287
rect 50436 56244 50488 56253
rect 50712 56287 50764 56296
rect 50712 56253 50721 56287
rect 50721 56253 50755 56287
rect 50755 56253 50764 56287
rect 50712 56244 50764 56253
rect 54208 56287 54260 56296
rect 54208 56253 54217 56287
rect 54217 56253 54251 56287
rect 54251 56253 54260 56287
rect 54208 56244 54260 56253
rect 54484 56287 54536 56296
rect 54484 56253 54493 56287
rect 54493 56253 54527 56287
rect 54527 56253 54536 56287
rect 54484 56244 54536 56253
rect 82912 56244 82964 56296
rect 41880 56219 41932 56228
rect 41880 56185 41889 56219
rect 41889 56185 41923 56219
rect 41923 56185 41932 56219
rect 41880 56176 41932 56185
rect 44640 56176 44692 56228
rect 48780 56176 48832 56228
rect 53380 56176 53432 56228
rect 75828 56176 75880 56228
rect 92664 56176 92716 56228
rect 11152 56108 11204 56160
rect 26516 56108 26568 56160
rect 26976 56108 27028 56160
rect 47768 56108 47820 56160
rect 50068 56108 50120 56160
rect 55496 56108 55548 56160
rect 85488 56108 85540 56160
rect 19606 56006 19658 56058
rect 19670 56006 19722 56058
rect 19734 56006 19786 56058
rect 19798 56006 19850 56058
rect 50326 56006 50378 56058
rect 50390 56006 50442 56058
rect 50454 56006 50506 56058
rect 50518 56006 50570 56058
rect 81046 56006 81098 56058
rect 81110 56006 81162 56058
rect 81174 56006 81226 56058
rect 81238 56006 81290 56058
rect 11612 55904 11664 55956
rect 80520 55904 80572 55956
rect 7012 55836 7064 55888
rect 77484 55836 77536 55888
rect 83740 55836 83792 55888
rect 85672 55836 85724 55888
rect 35256 55768 35308 55820
rect 11060 55632 11112 55684
rect 48780 55632 48832 55684
rect 34336 55564 34388 55616
rect 47768 55564 47820 55616
rect 49148 55768 49200 55820
rect 49516 55768 49568 55820
rect 49700 55768 49752 55820
rect 64052 55768 64104 55820
rect 76656 55768 76708 55820
rect 49056 55632 49108 55684
rect 59268 55700 59320 55752
rect 68744 55700 68796 55752
rect 80612 55700 80664 55752
rect 95056 55836 95108 55888
rect 49700 55564 49752 55616
rect 4246 55462 4298 55514
rect 4310 55462 4362 55514
rect 4374 55462 4426 55514
rect 4438 55462 4490 55514
rect 34966 55462 35018 55514
rect 35030 55462 35082 55514
rect 35094 55462 35146 55514
rect 35158 55462 35210 55514
rect 65686 55462 65738 55514
rect 65750 55462 65802 55514
rect 65814 55462 65866 55514
rect 65878 55462 65930 55514
rect 96406 55462 96458 55514
rect 96470 55462 96522 55514
rect 96534 55462 96586 55514
rect 96598 55462 96650 55514
rect 15108 55360 15160 55412
rect 56600 55360 56652 55412
rect 42708 55292 42760 55344
rect 62028 55292 62080 55344
rect 44272 55267 44324 55276
rect 44272 55233 44281 55267
rect 44281 55233 44315 55267
rect 44315 55233 44324 55267
rect 44272 55224 44324 55233
rect 49700 55224 49752 55276
rect 74816 55224 74868 55276
rect 75828 55224 75880 55276
rect 43628 55199 43680 55208
rect 43628 55165 43637 55199
rect 43637 55165 43671 55199
rect 43671 55165 43680 55199
rect 43628 55156 43680 55165
rect 44180 55199 44232 55208
rect 44180 55165 44189 55199
rect 44189 55165 44223 55199
rect 44223 55165 44232 55199
rect 44180 55156 44232 55165
rect 44456 55199 44508 55208
rect 44456 55165 44465 55199
rect 44465 55165 44499 55199
rect 44499 55165 44508 55199
rect 44456 55156 44508 55165
rect 43536 55088 43588 55140
rect 84108 55156 84160 55208
rect 91744 55156 91796 55208
rect 91928 55199 91980 55208
rect 91928 55165 91937 55199
rect 91937 55165 91971 55199
rect 91971 55165 91980 55199
rect 91928 55156 91980 55165
rect 61292 55131 61344 55140
rect 61292 55097 61301 55131
rect 61301 55097 61335 55131
rect 61335 55097 61344 55131
rect 61292 55088 61344 55097
rect 66352 55088 66404 55140
rect 66628 55088 66680 55140
rect 94044 55088 94096 55140
rect 14832 55020 14884 55072
rect 60464 55020 60516 55072
rect 19606 54918 19658 54970
rect 19670 54918 19722 54970
rect 19734 54918 19786 54970
rect 19798 54918 19850 54970
rect 50326 54918 50378 54970
rect 50390 54918 50442 54970
rect 50454 54918 50506 54970
rect 50518 54918 50570 54970
rect 81046 54918 81098 54970
rect 81110 54918 81162 54970
rect 81174 54918 81226 54970
rect 81238 54918 81290 54970
rect 1768 54816 1820 54868
rect 44456 54816 44508 54868
rect 46940 54816 46992 54868
rect 95424 54816 95476 54868
rect 84108 54791 84160 54800
rect 36544 54723 36596 54732
rect 36544 54689 36553 54723
rect 36553 54689 36587 54723
rect 36587 54689 36596 54723
rect 36544 54680 36596 54689
rect 33968 54612 34020 54664
rect 34428 54612 34480 54664
rect 79692 54680 79744 54732
rect 43444 54612 43496 54664
rect 53840 54612 53892 54664
rect 58256 54612 58308 54664
rect 76748 54612 76800 54664
rect 78128 54612 78180 54664
rect 84108 54757 84117 54791
rect 84117 54757 84151 54791
rect 84151 54757 84160 54791
rect 84108 54748 84160 54757
rect 83648 54723 83700 54732
rect 83648 54689 83657 54723
rect 83657 54689 83691 54723
rect 83691 54689 83700 54723
rect 83648 54680 83700 54689
rect 88616 54680 88668 54732
rect 32588 54476 32640 54528
rect 53012 54544 53064 54596
rect 78956 54544 79008 54596
rect 37832 54519 37884 54528
rect 37832 54485 37841 54519
rect 37841 54485 37875 54519
rect 37875 54485 37884 54519
rect 37832 54476 37884 54485
rect 69940 54476 69992 54528
rect 84568 54519 84620 54528
rect 84568 54485 84577 54519
rect 84577 54485 84611 54519
rect 84611 54485 84620 54519
rect 84568 54476 84620 54485
rect 84844 54519 84896 54528
rect 84844 54485 84853 54519
rect 84853 54485 84887 54519
rect 84887 54485 84896 54519
rect 84844 54476 84896 54485
rect 85948 54476 86000 54528
rect 4246 54374 4298 54426
rect 4310 54374 4362 54426
rect 4374 54374 4426 54426
rect 4438 54374 4490 54426
rect 34966 54374 35018 54426
rect 35030 54374 35082 54426
rect 35094 54374 35146 54426
rect 35158 54374 35210 54426
rect 65686 54374 65738 54426
rect 65750 54374 65802 54426
rect 65814 54374 65866 54426
rect 65878 54374 65930 54426
rect 96406 54374 96458 54426
rect 96470 54374 96522 54426
rect 96534 54374 96586 54426
rect 96598 54374 96650 54426
rect 1584 54136 1636 54188
rect 15936 54204 15988 54256
rect 6184 54068 6236 54120
rect 8944 54068 8996 54120
rect 25596 54111 25648 54120
rect 25596 54077 25605 54111
rect 25605 54077 25639 54111
rect 25639 54077 25648 54111
rect 25596 54068 25648 54077
rect 44916 54000 44968 54052
rect 46756 54000 46808 54052
rect 32404 53932 32456 53984
rect 45192 53932 45244 53984
rect 46848 53932 46900 53984
rect 19606 53830 19658 53882
rect 19670 53830 19722 53882
rect 19734 53830 19786 53882
rect 19798 53830 19850 53882
rect 50326 53830 50378 53882
rect 50390 53830 50442 53882
rect 50454 53830 50506 53882
rect 50518 53830 50570 53882
rect 81046 53830 81098 53882
rect 81110 53830 81162 53882
rect 81174 53830 81226 53882
rect 81238 53830 81290 53882
rect 14740 53635 14792 53644
rect 14740 53601 14749 53635
rect 14749 53601 14783 53635
rect 14783 53601 14792 53635
rect 14740 53592 14792 53601
rect 62856 53728 62908 53780
rect 15016 53567 15068 53576
rect 15016 53533 15025 53567
rect 15025 53533 15059 53567
rect 15059 53533 15068 53567
rect 15016 53524 15068 53533
rect 23940 53660 23992 53712
rect 24216 53660 24268 53712
rect 27712 53660 27764 53712
rect 28264 53660 28316 53712
rect 53380 53703 53432 53712
rect 53380 53669 53389 53703
rect 53389 53669 53423 53703
rect 53423 53669 53432 53703
rect 53380 53660 53432 53669
rect 53840 53703 53892 53712
rect 53840 53669 53849 53703
rect 53849 53669 53883 53703
rect 53883 53669 53892 53703
rect 53840 53660 53892 53669
rect 58716 53660 58768 53712
rect 21180 53635 21232 53644
rect 21180 53601 21188 53635
rect 21188 53601 21222 53635
rect 21222 53601 21232 53635
rect 21548 53635 21600 53644
rect 21180 53592 21232 53601
rect 21548 53601 21557 53635
rect 21557 53601 21591 53635
rect 21591 53601 21600 53635
rect 21548 53592 21600 53601
rect 54024 53635 54076 53644
rect 54024 53601 54027 53635
rect 54027 53601 54076 53635
rect 21364 53567 21416 53576
rect 21364 53533 21373 53567
rect 21373 53533 21407 53567
rect 21407 53533 21416 53567
rect 21364 53524 21416 53533
rect 27160 53524 27212 53576
rect 54024 53592 54076 53601
rect 60648 53592 60700 53644
rect 63040 53592 63092 53644
rect 62856 53524 62908 53576
rect 76104 53592 76156 53644
rect 79968 53592 80020 53644
rect 25688 53456 25740 53508
rect 54024 53456 54076 53508
rect 21088 53388 21140 53440
rect 21364 53388 21416 53440
rect 21640 53431 21692 53440
rect 21640 53397 21649 53431
rect 21649 53397 21683 53431
rect 21683 53397 21692 53431
rect 21640 53388 21692 53397
rect 54208 53388 54260 53440
rect 54392 53456 54444 53508
rect 81072 53456 81124 53508
rect 61016 53388 61068 53440
rect 4246 53286 4298 53338
rect 4310 53286 4362 53338
rect 4374 53286 4426 53338
rect 4438 53286 4490 53338
rect 34966 53286 35018 53338
rect 35030 53286 35082 53338
rect 35094 53286 35146 53338
rect 35158 53286 35210 53338
rect 65686 53286 65738 53338
rect 65750 53286 65802 53338
rect 65814 53286 65866 53338
rect 65878 53286 65930 53338
rect 96406 53286 96458 53338
rect 96470 53286 96522 53338
rect 96534 53286 96586 53338
rect 96598 53286 96650 53338
rect 7840 53184 7892 53236
rect 4436 53116 4488 53168
rect 6184 53116 6236 53168
rect 23020 53116 23072 53168
rect 28264 53116 28316 53168
rect 54024 53116 54076 53168
rect 58256 53116 58308 53168
rect 60464 53159 60516 53168
rect 60464 53125 60473 53159
rect 60473 53125 60507 53159
rect 60507 53125 60516 53159
rect 60464 53116 60516 53125
rect 5816 52912 5868 52964
rect 7564 52912 7616 52964
rect 3976 52844 4028 52896
rect 4988 52844 5040 52896
rect 11428 52844 11480 52896
rect 38292 53048 38344 53100
rect 61384 53116 61436 53168
rect 18696 52980 18748 53032
rect 46296 52980 46348 53032
rect 46848 52980 46900 53032
rect 57520 52980 57572 53032
rect 57704 53023 57756 53032
rect 57704 52989 57713 53023
rect 57713 52989 57747 53023
rect 57747 52989 57756 53023
rect 57704 52980 57756 52989
rect 57980 53023 58032 53032
rect 19892 52912 19944 52964
rect 46756 52912 46808 52964
rect 57980 52989 57989 53023
rect 57989 52989 58023 53023
rect 58023 52989 58032 53023
rect 57980 52980 58032 52989
rect 60648 53023 60700 53032
rect 60648 52989 60657 53023
rect 60657 52989 60691 53023
rect 60691 52989 60700 53023
rect 60648 52980 60700 52989
rect 60924 53023 60976 53032
rect 60924 52989 60933 53023
rect 60933 52989 60967 53023
rect 60967 52989 60976 53023
rect 60924 52980 60976 52989
rect 61016 52980 61068 53032
rect 64604 53116 64656 53168
rect 66904 53116 66956 53168
rect 71136 53116 71188 53168
rect 85764 53116 85816 53168
rect 66076 52980 66128 53032
rect 71688 53048 71740 53100
rect 81072 53091 81124 53100
rect 81072 53057 81081 53091
rect 81081 53057 81115 53091
rect 81115 53057 81124 53091
rect 81072 53048 81124 53057
rect 66996 52980 67048 53032
rect 62028 52912 62080 52964
rect 63684 52912 63736 52964
rect 67364 52887 67416 52896
rect 67364 52853 67373 52887
rect 67373 52853 67407 52887
rect 67407 52853 67416 52887
rect 67364 52844 67416 52853
rect 71780 52887 71832 52896
rect 71780 52853 71789 52887
rect 71789 52853 71823 52887
rect 71823 52853 71832 52887
rect 80704 52980 80756 53032
rect 95792 52980 95844 53032
rect 71780 52844 71832 52853
rect 19606 52742 19658 52794
rect 19670 52742 19722 52794
rect 19734 52742 19786 52794
rect 19798 52742 19850 52794
rect 50326 52742 50378 52794
rect 50390 52742 50442 52794
rect 50454 52742 50506 52794
rect 50518 52742 50570 52794
rect 81046 52742 81098 52794
rect 81110 52742 81162 52794
rect 81174 52742 81226 52794
rect 81238 52742 81290 52794
rect 3976 52683 4028 52692
rect 3976 52649 3985 52683
rect 3985 52649 4019 52683
rect 4019 52649 4028 52683
rect 3976 52640 4028 52649
rect 5080 52640 5132 52692
rect 5540 52640 5592 52692
rect 6460 52640 6512 52692
rect 7840 52640 7892 52692
rect 17868 52640 17920 52692
rect 4436 52547 4488 52556
rect 4436 52513 4445 52547
rect 4445 52513 4479 52547
rect 4479 52513 4488 52547
rect 4436 52504 4488 52513
rect 5816 52572 5868 52624
rect 7656 52615 7708 52624
rect 7656 52581 7665 52615
rect 7665 52581 7699 52615
rect 7699 52581 7708 52615
rect 7656 52572 7708 52581
rect 4988 52547 5040 52556
rect 4988 52513 4997 52547
rect 4997 52513 5031 52547
rect 5031 52513 5040 52547
rect 4988 52504 5040 52513
rect 7840 52547 7892 52556
rect 5540 52436 5592 52488
rect 6552 52436 6604 52488
rect 7840 52513 7849 52547
rect 7849 52513 7883 52547
rect 7883 52513 7892 52547
rect 7840 52504 7892 52513
rect 8116 52479 8168 52488
rect 8116 52445 8125 52479
rect 8125 52445 8159 52479
rect 8159 52445 8168 52479
rect 8116 52436 8168 52445
rect 45560 52640 45612 52692
rect 53656 52640 53708 52692
rect 57980 52640 58032 52692
rect 67364 52640 67416 52692
rect 42708 52615 42760 52624
rect 36268 52547 36320 52556
rect 36268 52513 36277 52547
rect 36277 52513 36311 52547
rect 36311 52513 36320 52547
rect 36268 52504 36320 52513
rect 36636 52547 36688 52556
rect 36636 52513 36645 52547
rect 36645 52513 36679 52547
rect 36679 52513 36688 52547
rect 36636 52504 36688 52513
rect 37004 52547 37056 52556
rect 37004 52513 37013 52547
rect 37013 52513 37047 52547
rect 37047 52513 37056 52547
rect 37004 52504 37056 52513
rect 38016 52504 38068 52556
rect 42156 52547 42208 52556
rect 42156 52513 42165 52547
rect 42165 52513 42199 52547
rect 42199 52513 42208 52547
rect 42156 52504 42208 52513
rect 42708 52581 42717 52615
rect 42717 52581 42751 52615
rect 42751 52581 42760 52615
rect 42708 52572 42760 52581
rect 57520 52572 57572 52624
rect 46480 52504 46532 52556
rect 54392 52504 54444 52556
rect 71136 52504 71188 52556
rect 74448 52504 74500 52556
rect 80152 52547 80204 52556
rect 80152 52513 80161 52547
rect 80161 52513 80195 52547
rect 80195 52513 80204 52547
rect 80152 52504 80204 52513
rect 80520 52547 80572 52556
rect 80520 52513 80529 52547
rect 80529 52513 80563 52547
rect 80563 52513 80572 52547
rect 80888 52547 80940 52556
rect 80520 52504 80572 52513
rect 80888 52513 80897 52547
rect 80897 52513 80931 52547
rect 80931 52513 80940 52547
rect 80888 52504 80940 52513
rect 33784 52436 33836 52488
rect 33968 52436 34020 52488
rect 36452 52479 36504 52488
rect 36452 52445 36461 52479
rect 36461 52445 36495 52479
rect 36495 52445 36504 52479
rect 36452 52436 36504 52445
rect 30196 52368 30248 52420
rect 37372 52479 37424 52488
rect 37372 52445 37381 52479
rect 37381 52445 37415 52479
rect 37415 52445 37424 52479
rect 37372 52436 37424 52445
rect 51724 52436 51776 52488
rect 52276 52436 52328 52488
rect 80980 52436 81032 52488
rect 82912 52436 82964 52488
rect 37832 52368 37884 52420
rect 83280 52368 83332 52420
rect 39304 52300 39356 52352
rect 64420 52300 64472 52352
rect 67364 52300 67416 52352
rect 71044 52300 71096 52352
rect 4246 52198 4298 52250
rect 4310 52198 4362 52250
rect 4374 52198 4426 52250
rect 4438 52198 4490 52250
rect 34966 52198 35018 52250
rect 35030 52198 35082 52250
rect 35094 52198 35146 52250
rect 35158 52198 35210 52250
rect 65686 52198 65738 52250
rect 65750 52198 65802 52250
rect 65814 52198 65866 52250
rect 65878 52198 65930 52250
rect 96406 52198 96458 52250
rect 96470 52198 96522 52250
rect 96534 52198 96586 52250
rect 96598 52198 96650 52250
rect 54576 52096 54628 52148
rect 10600 52028 10652 52080
rect 52644 52028 52696 52080
rect 58808 52028 58860 52080
rect 21364 51960 21416 52012
rect 29552 51960 29604 52012
rect 9864 51892 9916 51944
rect 24216 51892 24268 51944
rect 37004 51892 37056 51944
rect 41880 51892 41932 51944
rect 54576 51935 54628 51944
rect 54576 51901 54585 51935
rect 54585 51901 54619 51935
rect 54619 51901 54628 51935
rect 54576 51892 54628 51901
rect 59268 51935 59320 51944
rect 59268 51901 59277 51935
rect 59277 51901 59311 51935
rect 59311 51901 59320 51935
rect 59268 51892 59320 51901
rect 66352 51892 66404 51944
rect 10600 51824 10652 51876
rect 36636 51824 36688 51876
rect 42156 51824 42208 51876
rect 55128 51867 55180 51876
rect 55128 51833 55137 51867
rect 55137 51833 55171 51867
rect 55171 51833 55180 51867
rect 55128 51824 55180 51833
rect 80520 51824 80572 51876
rect 80980 51824 81032 51876
rect 12164 51756 12216 51808
rect 21640 51756 21692 51808
rect 23112 51756 23164 51808
rect 37832 51756 37884 51808
rect 43076 51756 43128 51808
rect 62028 51756 62080 51808
rect 19606 51654 19658 51706
rect 19670 51654 19722 51706
rect 19734 51654 19786 51706
rect 19798 51654 19850 51706
rect 50326 51654 50378 51706
rect 50390 51654 50442 51706
rect 50454 51654 50506 51706
rect 50518 51654 50570 51706
rect 81046 51654 81098 51706
rect 81110 51654 81162 51706
rect 81174 51654 81226 51706
rect 81238 51654 81290 51706
rect 83280 51552 83332 51604
rect 83740 51552 83792 51604
rect 29920 51348 29972 51400
rect 39672 51212 39724 51264
rect 41696 51255 41748 51264
rect 41696 51221 41705 51255
rect 41705 51221 41739 51255
rect 41739 51221 41748 51255
rect 41696 51212 41748 51221
rect 61384 51212 61436 51264
rect 4246 51110 4298 51162
rect 4310 51110 4362 51162
rect 4374 51110 4426 51162
rect 4438 51110 4490 51162
rect 34966 51110 35018 51162
rect 35030 51110 35082 51162
rect 35094 51110 35146 51162
rect 35158 51110 35210 51162
rect 65686 51110 65738 51162
rect 65750 51110 65802 51162
rect 65814 51110 65866 51162
rect 65878 51110 65930 51162
rect 96406 51110 96458 51162
rect 96470 51110 96522 51162
rect 96534 51110 96586 51162
rect 96598 51110 96650 51162
rect 14924 51008 14976 51060
rect 18972 51008 19024 51060
rect 49516 51008 49568 51060
rect 22468 50940 22520 50992
rect 56048 50940 56100 50992
rect 1124 50872 1176 50924
rect 48044 50872 48096 50924
rect 47584 50847 47636 50856
rect 47584 50813 47593 50847
rect 47593 50813 47627 50847
rect 47627 50813 47636 50847
rect 47584 50804 47636 50813
rect 13452 50736 13504 50788
rect 85212 50736 85264 50788
rect 8668 50668 8720 50720
rect 23296 50668 23348 50720
rect 28356 50668 28408 50720
rect 32956 50668 33008 50720
rect 33600 50668 33652 50720
rect 34428 50668 34480 50720
rect 42340 50668 42392 50720
rect 47584 50668 47636 50720
rect 19606 50566 19658 50618
rect 19670 50566 19722 50618
rect 19734 50566 19786 50618
rect 19798 50566 19850 50618
rect 50326 50566 50378 50618
rect 50390 50566 50442 50618
rect 50454 50566 50506 50618
rect 50518 50566 50570 50618
rect 81046 50566 81098 50618
rect 81110 50566 81162 50618
rect 81174 50566 81226 50618
rect 81238 50566 81290 50618
rect 60096 50464 60148 50516
rect 32956 50396 33008 50448
rect 48044 50439 48096 50448
rect 18788 50328 18840 50380
rect 19892 50328 19944 50380
rect 24492 50328 24544 50380
rect 27804 50328 27856 50380
rect 28356 50328 28408 50380
rect 22468 50303 22520 50312
rect 22468 50269 22477 50303
rect 22477 50269 22511 50303
rect 22511 50269 22520 50303
rect 22468 50260 22520 50269
rect 30380 50260 30432 50312
rect 33600 50328 33652 50380
rect 48044 50405 48053 50439
rect 48053 50405 48087 50439
rect 48087 50405 48096 50439
rect 48044 50396 48096 50405
rect 53380 50396 53432 50448
rect 53748 50396 53800 50448
rect 63776 50396 63828 50448
rect 64696 50396 64748 50448
rect 75368 50396 75420 50448
rect 32220 50303 32272 50312
rect 32220 50269 32229 50303
rect 32229 50269 32263 50303
rect 32263 50269 32272 50303
rect 32220 50260 32272 50269
rect 8300 50192 8352 50244
rect 19524 50192 19576 50244
rect 2044 50124 2096 50176
rect 22652 50192 22704 50244
rect 90456 50371 90508 50380
rect 90456 50337 90465 50371
rect 90465 50337 90499 50371
rect 90499 50337 90508 50371
rect 90456 50328 90508 50337
rect 65064 50260 65116 50312
rect 75184 50260 75236 50312
rect 22284 50167 22336 50176
rect 22284 50133 22293 50167
rect 22293 50133 22327 50167
rect 22327 50133 22336 50167
rect 22284 50124 22336 50133
rect 23848 50124 23900 50176
rect 33416 50124 33468 50176
rect 36820 50124 36872 50176
rect 71596 50192 71648 50244
rect 84568 50124 84620 50176
rect 4246 50022 4298 50074
rect 4310 50022 4362 50074
rect 4374 50022 4426 50074
rect 4438 50022 4490 50074
rect 34966 50022 35018 50074
rect 35030 50022 35082 50074
rect 35094 50022 35146 50074
rect 35158 50022 35210 50074
rect 65686 50022 65738 50074
rect 65750 50022 65802 50074
rect 65814 50022 65866 50074
rect 65878 50022 65930 50074
rect 96406 50022 96458 50074
rect 96470 50022 96522 50074
rect 96534 50022 96586 50074
rect 96598 50022 96650 50074
rect 13452 49963 13504 49972
rect 13452 49929 13461 49963
rect 13461 49929 13495 49963
rect 13495 49929 13504 49963
rect 13452 49920 13504 49929
rect 17868 49920 17920 49972
rect 22928 49920 22980 49972
rect 23020 49920 23072 49972
rect 84844 49920 84896 49972
rect 1400 49759 1452 49768
rect 1400 49725 1409 49759
rect 1409 49725 1443 49759
rect 1443 49725 1452 49759
rect 1400 49716 1452 49725
rect 12256 49759 12308 49768
rect 12256 49725 12265 49759
rect 12265 49725 12299 49759
rect 12299 49725 12308 49759
rect 12256 49716 12308 49725
rect 15108 49852 15160 49904
rect 24032 49895 24084 49904
rect 24032 49861 24041 49895
rect 24041 49861 24075 49895
rect 24075 49861 24084 49895
rect 24032 49852 24084 49861
rect 49516 49852 49568 49904
rect 63776 49852 63828 49904
rect 67640 49852 67692 49904
rect 82268 49784 82320 49836
rect 12992 49759 13044 49768
rect 12992 49725 13001 49759
rect 13001 49725 13035 49759
rect 13035 49725 13044 49759
rect 12992 49716 13044 49725
rect 17408 49716 17460 49768
rect 19524 49716 19576 49768
rect 22652 49716 22704 49768
rect 22928 49759 22980 49768
rect 22928 49725 22937 49759
rect 22937 49725 22971 49759
rect 22971 49725 22980 49759
rect 22928 49716 22980 49725
rect 23020 49716 23072 49768
rect 23296 49759 23348 49768
rect 23296 49725 23305 49759
rect 23305 49725 23339 49759
rect 23339 49725 23348 49759
rect 23848 49759 23900 49768
rect 23296 49716 23348 49725
rect 23848 49725 23857 49759
rect 23857 49725 23891 49759
rect 23891 49725 23900 49759
rect 23848 49716 23900 49725
rect 30380 49716 30432 49768
rect 30564 49759 30616 49768
rect 30564 49725 30573 49759
rect 30573 49725 30607 49759
rect 30607 49725 30616 49759
rect 30564 49716 30616 49725
rect 31760 49716 31812 49768
rect 48412 49716 48464 49768
rect 49516 49716 49568 49768
rect 55956 49759 56008 49768
rect 55956 49725 55965 49759
rect 55965 49725 55999 49759
rect 55999 49725 56008 49759
rect 55956 49716 56008 49725
rect 22376 49623 22428 49632
rect 22376 49589 22385 49623
rect 22385 49589 22419 49623
rect 22419 49589 22428 49623
rect 22376 49580 22428 49589
rect 23020 49580 23072 49632
rect 43352 49648 43404 49700
rect 48228 49648 48280 49700
rect 31576 49580 31628 49632
rect 71688 49759 71740 49768
rect 71688 49725 71697 49759
rect 71697 49725 71731 49759
rect 71731 49725 71740 49759
rect 71688 49716 71740 49725
rect 19606 49478 19658 49530
rect 19670 49478 19722 49530
rect 19734 49478 19786 49530
rect 19798 49478 19850 49530
rect 50326 49478 50378 49530
rect 50390 49478 50442 49530
rect 50454 49478 50506 49530
rect 50518 49478 50570 49530
rect 81046 49478 81098 49530
rect 81110 49478 81162 49530
rect 81174 49478 81226 49530
rect 81238 49478 81290 49530
rect 24032 49376 24084 49428
rect 69664 49376 69716 49428
rect 70124 49376 70176 49428
rect 82728 49376 82780 49428
rect 28448 49308 28500 49360
rect 31576 49308 31628 49360
rect 81992 49308 82044 49360
rect 15016 49240 15068 49292
rect 76196 49240 76248 49292
rect 92848 49240 92900 49292
rect 36728 49172 36780 49224
rect 38200 49172 38252 49224
rect 42340 49215 42392 49224
rect 42340 49181 42349 49215
rect 42349 49181 42383 49215
rect 42383 49181 42392 49215
rect 42340 49172 42392 49181
rect 46204 49172 46256 49224
rect 58808 49172 58860 49224
rect 78036 49172 78088 49224
rect 84200 49215 84252 49224
rect 84200 49181 84209 49215
rect 84209 49181 84243 49215
rect 84243 49181 84252 49215
rect 84200 49172 84252 49181
rect 85948 49215 86000 49224
rect 85948 49181 85957 49215
rect 85957 49181 85991 49215
rect 85991 49181 86000 49215
rect 85948 49172 86000 49181
rect 3700 49104 3752 49156
rect 12992 49104 13044 49156
rect 19248 49104 19300 49156
rect 25872 49104 25924 49156
rect 36084 49104 36136 49156
rect 43352 49104 43404 49156
rect 47032 49104 47084 49156
rect 48228 49104 48280 49156
rect 53748 49104 53800 49156
rect 55404 49104 55456 49156
rect 16120 49036 16172 49088
rect 22652 49079 22704 49088
rect 22652 49045 22661 49079
rect 22661 49045 22695 49079
rect 22695 49045 22704 49079
rect 22652 49036 22704 49045
rect 24308 49079 24360 49088
rect 24308 49045 24317 49079
rect 24317 49045 24351 49079
rect 24351 49045 24360 49079
rect 24308 49036 24360 49045
rect 43720 49079 43772 49088
rect 43720 49045 43729 49079
rect 43729 49045 43763 49079
rect 43763 49045 43772 49079
rect 43720 49036 43772 49045
rect 4246 48934 4298 48986
rect 4310 48934 4362 48986
rect 4374 48934 4426 48986
rect 4438 48934 4490 48986
rect 34966 48934 35018 48986
rect 35030 48934 35082 48986
rect 35094 48934 35146 48986
rect 35158 48934 35210 48986
rect 65686 48934 65738 48986
rect 65750 48934 65802 48986
rect 65814 48934 65866 48986
rect 65878 48934 65930 48986
rect 96406 48934 96458 48986
rect 96470 48934 96522 48986
rect 96534 48934 96586 48986
rect 96598 48934 96650 48986
rect 24308 48832 24360 48884
rect 30104 48832 30156 48884
rect 48964 48832 49016 48884
rect 84200 48832 84252 48884
rect 18604 48764 18656 48816
rect 15384 48696 15436 48748
rect 22652 48764 22704 48816
rect 87512 48764 87564 48816
rect 18972 48671 19024 48680
rect 18972 48637 18981 48671
rect 18981 48637 19015 48671
rect 19015 48637 19024 48671
rect 18972 48628 19024 48637
rect 19248 48671 19300 48680
rect 19248 48637 19257 48671
rect 19257 48637 19291 48671
rect 19291 48637 19300 48671
rect 19248 48628 19300 48637
rect 67548 48696 67600 48748
rect 22836 48560 22888 48612
rect 23940 48560 23992 48612
rect 24216 48560 24268 48612
rect 65064 48628 65116 48680
rect 67732 48671 67784 48680
rect 67732 48637 67741 48671
rect 67741 48637 67775 48671
rect 67775 48637 67784 48671
rect 67732 48628 67784 48637
rect 52460 48560 52512 48612
rect 20536 48492 20588 48544
rect 19606 48390 19658 48442
rect 19670 48390 19722 48442
rect 19734 48390 19786 48442
rect 19798 48390 19850 48442
rect 50326 48390 50378 48442
rect 50390 48390 50442 48442
rect 50454 48390 50506 48442
rect 50518 48390 50570 48442
rect 81046 48390 81098 48442
rect 81110 48390 81162 48442
rect 81174 48390 81226 48442
rect 81238 48390 81290 48442
rect 4896 48195 4948 48204
rect 4896 48161 4905 48195
rect 4905 48161 4939 48195
rect 4939 48161 4948 48195
rect 4896 48152 4948 48161
rect 34060 48220 34112 48272
rect 42340 48152 42392 48204
rect 36636 48084 36688 48136
rect 45284 48288 45336 48340
rect 52460 48152 52512 48204
rect 53196 48152 53248 48204
rect 58256 48220 58308 48272
rect 63592 48220 63644 48272
rect 64512 48220 64564 48272
rect 91744 48220 91796 48272
rect 57888 48195 57940 48204
rect 57888 48161 57897 48195
rect 57897 48161 57931 48195
rect 57931 48161 57940 48195
rect 57888 48152 57940 48161
rect 52000 48084 52052 48136
rect 58072 48152 58124 48204
rect 83648 48152 83700 48204
rect 8300 48016 8352 48068
rect 8392 48016 8444 48068
rect 11796 47948 11848 48000
rect 37832 47991 37884 48000
rect 37832 47957 37841 47991
rect 37841 47957 37875 47991
rect 37875 47957 37884 47991
rect 37832 47948 37884 47957
rect 46020 47991 46072 48000
rect 46020 47957 46029 47991
rect 46029 47957 46063 47991
rect 46063 47957 46072 47991
rect 46020 47948 46072 47957
rect 57428 47948 57480 48000
rect 58256 47991 58308 48000
rect 58256 47957 58265 47991
rect 58265 47957 58299 47991
rect 58299 47957 58308 47991
rect 58256 47948 58308 47957
rect 71688 47948 71740 48000
rect 83096 47948 83148 48000
rect 92480 47948 92532 48000
rect 4246 47846 4298 47898
rect 4310 47846 4362 47898
rect 4374 47846 4426 47898
rect 4438 47846 4490 47898
rect 34966 47846 35018 47898
rect 35030 47846 35082 47898
rect 35094 47846 35146 47898
rect 35158 47846 35210 47898
rect 65686 47846 65738 47898
rect 65750 47846 65802 47898
rect 65814 47846 65866 47898
rect 65878 47846 65930 47898
rect 96406 47846 96458 47898
rect 96470 47846 96522 47898
rect 96534 47846 96586 47898
rect 96598 47846 96650 47898
rect 5724 47744 5776 47796
rect 8392 47744 8444 47796
rect 28448 47787 28500 47796
rect 28448 47753 28457 47787
rect 28457 47753 28491 47787
rect 28491 47753 28500 47787
rect 28448 47744 28500 47753
rect 28816 47744 28868 47796
rect 57428 47744 57480 47796
rect 73988 47744 74040 47796
rect 86960 47744 87012 47796
rect 91744 47744 91796 47796
rect 7104 47676 7156 47728
rect 57888 47676 57940 47728
rect 71228 47676 71280 47728
rect 27528 47608 27580 47660
rect 28172 47651 28224 47660
rect 7472 47540 7524 47592
rect 21824 47540 21876 47592
rect 28172 47617 28181 47651
rect 28181 47617 28215 47651
rect 28215 47617 28224 47651
rect 28172 47608 28224 47617
rect 27528 47404 27580 47456
rect 27988 47583 28040 47592
rect 27988 47549 27996 47583
rect 27996 47549 28030 47583
rect 28030 47549 28040 47583
rect 27988 47540 28040 47549
rect 54760 47608 54812 47660
rect 63408 47608 63460 47660
rect 73896 47540 73948 47592
rect 76656 47540 76708 47592
rect 77300 47540 77352 47592
rect 86684 47608 86736 47660
rect 92480 47651 92532 47660
rect 92480 47617 92489 47651
rect 92489 47617 92523 47651
rect 92523 47617 92532 47651
rect 92480 47608 92532 47617
rect 86868 47540 86920 47592
rect 86960 47583 87012 47592
rect 86960 47549 86969 47583
rect 86969 47549 87003 47583
rect 87003 47549 87012 47583
rect 86960 47540 87012 47549
rect 87328 47583 87380 47592
rect 36728 47472 36780 47524
rect 36912 47472 36964 47524
rect 62396 47472 62448 47524
rect 86684 47472 86736 47524
rect 87328 47549 87337 47583
rect 87337 47549 87371 47583
rect 87371 47549 87380 47583
rect 87328 47540 87380 47549
rect 87420 47540 87472 47592
rect 87604 47472 87656 47524
rect 87972 47540 88024 47592
rect 91744 47540 91796 47592
rect 86868 47404 86920 47456
rect 92848 47583 92900 47592
rect 92848 47549 92857 47583
rect 92857 47549 92891 47583
rect 92891 47549 92900 47583
rect 92848 47540 92900 47549
rect 88156 47447 88208 47456
rect 88156 47413 88165 47447
rect 88165 47413 88199 47447
rect 88199 47413 88208 47447
rect 88156 47404 88208 47413
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 50326 47302 50378 47354
rect 50390 47302 50442 47354
rect 50454 47302 50506 47354
rect 50518 47302 50570 47354
rect 81046 47302 81098 47354
rect 81110 47302 81162 47354
rect 81174 47302 81226 47354
rect 81238 47302 81290 47354
rect 8208 47200 8260 47252
rect 31484 47200 31536 47252
rect 88156 47200 88208 47252
rect 38016 47132 38068 47184
rect 74080 47132 74132 47184
rect 77300 47132 77352 47184
rect 87420 47132 87472 47184
rect 14740 47064 14792 47116
rect 37096 47064 37148 47116
rect 64696 47107 64748 47116
rect 50804 46996 50856 47048
rect 64696 47073 64705 47107
rect 64705 47073 64739 47107
rect 64739 47073 64748 47107
rect 64696 47064 64748 47073
rect 65064 47107 65116 47116
rect 65064 47073 65078 47107
rect 65078 47073 65112 47107
rect 65112 47073 65116 47107
rect 65064 47064 65116 47073
rect 76012 47064 76064 47116
rect 76288 47064 76340 47116
rect 77116 47064 77168 47116
rect 87328 47064 87380 47116
rect 68928 46996 68980 47048
rect 9956 46860 10008 46912
rect 27068 46928 27120 46980
rect 27528 46928 27580 46980
rect 58900 46928 58952 46980
rect 65248 46971 65300 46980
rect 34336 46860 34388 46912
rect 45376 46860 45428 46912
rect 65248 46937 65257 46971
rect 65257 46937 65291 46971
rect 65291 46937 65300 46971
rect 65248 46928 65300 46937
rect 73252 46860 73304 46912
rect 79508 46860 79560 46912
rect 81532 46860 81584 46912
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 65686 46758 65738 46810
rect 65750 46758 65802 46810
rect 65814 46758 65866 46810
rect 65878 46758 65930 46810
rect 96406 46758 96458 46810
rect 96470 46758 96522 46810
rect 96534 46758 96586 46810
rect 96598 46758 96650 46810
rect 11888 46656 11940 46708
rect 14832 46656 14884 46708
rect 25688 46656 25740 46708
rect 75828 46656 75880 46708
rect 76012 46656 76064 46708
rect 18420 46588 18472 46640
rect 96896 46588 96948 46640
rect 19248 46563 19300 46572
rect 19248 46529 19257 46563
rect 19257 46529 19291 46563
rect 19291 46529 19300 46563
rect 19248 46520 19300 46529
rect 43260 46520 43312 46572
rect 71780 46520 71832 46572
rect 74264 46520 74316 46572
rect 13636 46359 13688 46368
rect 13636 46325 13645 46359
rect 13645 46325 13679 46359
rect 13679 46325 13688 46359
rect 13636 46316 13688 46325
rect 14740 46452 14792 46504
rect 14832 46495 14884 46504
rect 14832 46461 14841 46495
rect 14841 46461 14875 46495
rect 14875 46461 14884 46495
rect 18696 46495 18748 46504
rect 14832 46452 14884 46461
rect 18696 46461 18705 46495
rect 18705 46461 18739 46495
rect 18739 46461 18748 46495
rect 18696 46452 18748 46461
rect 66168 46384 66220 46436
rect 81532 46384 81584 46436
rect 87788 46495 87840 46504
rect 16488 46316 16540 46368
rect 71228 46316 71280 46368
rect 74264 46316 74316 46368
rect 84844 46316 84896 46368
rect 87788 46461 87797 46495
rect 87797 46461 87831 46495
rect 87831 46461 87840 46495
rect 87788 46452 87840 46461
rect 88156 46520 88208 46572
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 50326 46214 50378 46266
rect 50390 46214 50442 46266
rect 50454 46214 50506 46266
rect 50518 46214 50570 46266
rect 81046 46214 81098 46266
rect 81110 46214 81162 46266
rect 81174 46214 81226 46266
rect 81238 46214 81290 46266
rect 11244 46112 11296 46164
rect 11612 46112 11664 46164
rect 14740 46112 14792 46164
rect 16948 46112 17000 46164
rect 53564 46112 53616 46164
rect 60372 46112 60424 46164
rect 9680 46044 9732 46096
rect 18696 46044 18748 46096
rect 34336 46044 34388 46096
rect 87788 46044 87840 46096
rect 13636 45976 13688 46028
rect 90548 45976 90600 46028
rect 77668 45772 77720 45824
rect 85948 45772 86000 45824
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 65686 45670 65738 45722
rect 65750 45670 65802 45722
rect 65814 45670 65866 45722
rect 65878 45670 65930 45722
rect 96406 45670 96458 45722
rect 96470 45670 96522 45722
rect 96534 45670 96586 45722
rect 96598 45670 96650 45722
rect 3056 45500 3108 45552
rect 10324 45432 10376 45484
rect 77852 45568 77904 45620
rect 17316 45432 17368 45484
rect 41880 45432 41932 45484
rect 77668 45500 77720 45552
rect 90456 45500 90508 45552
rect 6644 45364 6696 45416
rect 26884 45364 26936 45416
rect 47584 45364 47636 45416
rect 77852 45432 77904 45484
rect 7656 45296 7708 45348
rect 18144 45296 18196 45348
rect 40316 45296 40368 45348
rect 63132 45296 63184 45348
rect 74264 45296 74316 45348
rect 82268 45296 82320 45348
rect 15108 45228 15160 45280
rect 21364 45228 21416 45280
rect 23296 45228 23348 45280
rect 44272 45228 44324 45280
rect 57888 45228 57940 45280
rect 82452 45228 82504 45280
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 50326 45126 50378 45178
rect 50390 45126 50442 45178
rect 50454 45126 50506 45178
rect 50518 45126 50570 45178
rect 81046 45126 81098 45178
rect 81110 45126 81162 45178
rect 81174 45126 81226 45178
rect 81238 45126 81290 45178
rect 8116 45024 8168 45076
rect 58900 45024 58952 45076
rect 70676 45024 70728 45076
rect 4804 44956 4856 45008
rect 7656 44888 7708 44940
rect 17316 44956 17368 45008
rect 21364 44956 21416 45008
rect 72516 44956 72568 45008
rect 17960 44931 18012 44940
rect 17960 44897 17969 44931
rect 17969 44897 18003 44931
rect 18003 44897 18012 44931
rect 18236 44931 18288 44940
rect 17960 44888 18012 44897
rect 18236 44897 18245 44931
rect 18245 44897 18279 44931
rect 18279 44897 18288 44931
rect 18236 44888 18288 44897
rect 19248 44888 19300 44940
rect 57980 44888 58032 44940
rect 74264 44999 74316 45008
rect 74264 44965 74273 44999
rect 74273 44965 74307 44999
rect 74307 44965 74316 44999
rect 74264 44956 74316 44965
rect 73160 44888 73212 44940
rect 4620 44752 4672 44804
rect 1676 44727 1728 44736
rect 1676 44693 1685 44727
rect 1685 44693 1719 44727
rect 1719 44693 1728 44727
rect 1676 44684 1728 44693
rect 6644 44727 6696 44736
rect 6644 44693 6653 44727
rect 6653 44693 6687 44727
rect 6687 44693 6696 44727
rect 6644 44684 6696 44693
rect 18604 44820 18656 44872
rect 32404 44820 32456 44872
rect 54760 44820 54812 44872
rect 64788 44820 64840 44872
rect 74448 44931 74500 44940
rect 74448 44897 74462 44931
rect 74462 44897 74496 44931
rect 74496 44897 74500 44931
rect 74448 44888 74500 44897
rect 17960 44752 18012 44804
rect 18236 44684 18288 44736
rect 45928 44684 45980 44736
rect 74632 44727 74684 44736
rect 74632 44693 74641 44727
rect 74641 44693 74675 44727
rect 74675 44693 74684 44727
rect 74632 44684 74684 44693
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 65686 44582 65738 44634
rect 65750 44582 65802 44634
rect 65814 44582 65866 44634
rect 65878 44582 65930 44634
rect 96406 44582 96458 44634
rect 96470 44582 96522 44634
rect 96534 44582 96586 44634
rect 96598 44582 96650 44634
rect 40316 44412 40368 44464
rect 41880 44412 41932 44464
rect 17684 44276 17736 44328
rect 23572 44319 23624 44328
rect 23572 44285 23581 44319
rect 23581 44285 23615 44319
rect 23615 44285 23624 44319
rect 23572 44276 23624 44285
rect 62856 44276 62908 44328
rect 44272 44208 44324 44260
rect 45100 44208 45152 44260
rect 70492 44344 70544 44396
rect 71688 44344 71740 44396
rect 24860 44183 24912 44192
rect 24860 44149 24869 44183
rect 24869 44149 24903 44183
rect 24903 44149 24912 44183
rect 24860 44140 24912 44149
rect 46848 44140 46900 44192
rect 53748 44140 53800 44192
rect 69572 44183 69624 44192
rect 69572 44149 69581 44183
rect 69581 44149 69615 44183
rect 69615 44149 69624 44183
rect 69572 44140 69624 44149
rect 84936 44140 84988 44192
rect 86500 44140 86552 44192
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 50326 44038 50378 44090
rect 50390 44038 50442 44090
rect 50454 44038 50506 44090
rect 50518 44038 50570 44090
rect 81046 44038 81098 44090
rect 81110 44038 81162 44090
rect 81174 44038 81226 44090
rect 81238 44038 81290 44090
rect 10416 43936 10468 43988
rect 39764 43936 39816 43988
rect 72424 43936 72476 43988
rect 72976 43936 73028 43988
rect 74080 43936 74132 43988
rect 78128 43936 78180 43988
rect 64328 43868 64380 43920
rect 66720 43868 66772 43920
rect 24584 43800 24636 43852
rect 24492 43732 24544 43784
rect 31024 43732 31076 43784
rect 37556 43775 37608 43784
rect 37556 43741 37565 43775
rect 37565 43741 37599 43775
rect 37599 43741 37608 43775
rect 37556 43732 37608 43741
rect 59544 43732 59596 43784
rect 38844 43707 38896 43716
rect 38844 43673 38853 43707
rect 38853 43673 38887 43707
rect 38887 43673 38896 43707
rect 38844 43664 38896 43673
rect 40040 43664 40092 43716
rect 69204 43664 69256 43716
rect 63132 43596 63184 43648
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 65686 43494 65738 43546
rect 65750 43494 65802 43546
rect 65814 43494 65866 43546
rect 65878 43494 65930 43546
rect 96406 43494 96458 43546
rect 96470 43494 96522 43546
rect 96534 43494 96586 43546
rect 96598 43494 96650 43546
rect 7656 43392 7708 43444
rect 35256 43392 35308 43444
rect 38844 43392 38896 43444
rect 50804 43392 50856 43444
rect 52184 43392 52236 43444
rect 82360 43392 82412 43444
rect 16488 43324 16540 43376
rect 38660 43324 38712 43376
rect 29828 43256 29880 43308
rect 40040 43367 40092 43376
rect 40040 43333 40049 43367
rect 40049 43333 40083 43367
rect 40083 43333 40092 43367
rect 40040 43324 40092 43333
rect 45100 43299 45152 43308
rect 45100 43265 45109 43299
rect 45109 43265 45143 43299
rect 45143 43265 45152 43299
rect 45100 43256 45152 43265
rect 82544 43256 82596 43308
rect 40224 43231 40276 43240
rect 40224 43197 40233 43231
rect 40233 43197 40267 43231
rect 40267 43197 40276 43231
rect 40224 43188 40276 43197
rect 44732 43231 44784 43240
rect 40500 43163 40552 43172
rect 40500 43129 40509 43163
rect 40509 43129 40543 43163
rect 40543 43129 40552 43163
rect 40500 43120 40552 43129
rect 44732 43197 44741 43231
rect 44741 43197 44775 43231
rect 44775 43197 44784 43231
rect 44732 43188 44784 43197
rect 59544 43231 59596 43240
rect 59544 43197 59553 43231
rect 59553 43197 59587 43231
rect 59587 43197 59596 43231
rect 94044 43256 94096 43308
rect 59544 43188 59596 43197
rect 53656 43120 53708 43172
rect 56048 43120 56100 43172
rect 55128 43052 55180 43104
rect 58348 43052 58400 43104
rect 58624 43052 58676 43104
rect 71136 43052 71188 43104
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 50326 42950 50378 43002
rect 50390 42950 50442 43002
rect 50454 42950 50506 43002
rect 50518 42950 50570 43002
rect 81046 42950 81098 43002
rect 81110 42950 81162 43002
rect 81174 42950 81226 43002
rect 81238 42950 81290 43002
rect 38660 42848 38712 42900
rect 42892 42848 42944 42900
rect 72424 42848 72476 42900
rect 17408 42780 17460 42832
rect 80888 42780 80940 42832
rect 85580 42780 85632 42832
rect 12072 42712 12124 42764
rect 12256 42712 12308 42764
rect 46112 42712 46164 42764
rect 49424 42712 49476 42764
rect 60740 42712 60792 42764
rect 73528 42755 73580 42764
rect 73528 42721 73537 42755
rect 73537 42721 73571 42755
rect 73571 42721 73580 42755
rect 73528 42712 73580 42721
rect 74448 42712 74500 42764
rect 78680 42712 78732 42764
rect 79968 42712 80020 42764
rect 86224 42712 86276 42764
rect 21548 42644 21600 42696
rect 72516 42687 72568 42696
rect 72516 42653 72525 42687
rect 72525 42653 72559 42687
rect 72559 42653 72568 42687
rect 72516 42644 72568 42653
rect 73068 42687 73120 42696
rect 73068 42653 73077 42687
rect 73077 42653 73111 42687
rect 73111 42653 73120 42687
rect 73068 42644 73120 42653
rect 55956 42576 56008 42628
rect 62212 42508 62264 42560
rect 73528 42508 73580 42560
rect 80704 42619 80756 42628
rect 80704 42585 80713 42619
rect 80713 42585 80747 42619
rect 80747 42585 80756 42619
rect 80704 42576 80756 42585
rect 91928 42576 91980 42628
rect 86592 42508 86644 42560
rect 86868 42508 86920 42560
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 65686 42406 65738 42458
rect 65750 42406 65802 42458
rect 65814 42406 65866 42458
rect 65878 42406 65930 42458
rect 96406 42406 96458 42458
rect 96470 42406 96522 42458
rect 96534 42406 96586 42458
rect 96598 42406 96650 42458
rect 72516 42304 72568 42356
rect 72884 42304 72936 42356
rect 95700 42236 95752 42288
rect 96528 42236 96580 42288
rect 39764 42168 39816 42220
rect 92848 42211 92900 42220
rect 16948 42100 17000 42152
rect 42800 42100 42852 42152
rect 16212 42032 16264 42084
rect 21548 42032 21600 42084
rect 44364 42007 44416 42016
rect 44364 41973 44373 42007
rect 44373 41973 44407 42007
rect 44407 41973 44416 42007
rect 92848 42177 92857 42211
rect 92857 42177 92891 42211
rect 92891 42177 92900 42211
rect 92848 42168 92900 42177
rect 92572 42143 92624 42152
rect 92572 42109 92581 42143
rect 92581 42109 92615 42143
rect 92615 42109 92624 42143
rect 92572 42100 92624 42109
rect 78680 42032 78732 42084
rect 44364 41964 44416 41973
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 50326 41862 50378 41914
rect 50390 41862 50442 41914
rect 50454 41862 50506 41914
rect 50518 41862 50570 41914
rect 81046 41862 81098 41914
rect 81110 41862 81162 41914
rect 81174 41862 81226 41914
rect 81238 41862 81290 41914
rect 80060 41760 80112 41812
rect 80428 41760 80480 41812
rect 42800 41692 42852 41744
rect 42984 41692 43036 41744
rect 72516 41692 72568 41744
rect 86868 41692 86920 41744
rect 29276 41624 29328 41676
rect 95516 41624 95568 41676
rect 31300 41599 31352 41608
rect 31300 41565 31309 41599
rect 31309 41565 31343 41599
rect 31343 41565 31352 41599
rect 31300 41556 31352 41565
rect 49424 41599 49476 41608
rect 49424 41565 49433 41599
rect 49433 41565 49467 41599
rect 49467 41565 49476 41599
rect 49424 41556 49476 41565
rect 96160 41599 96212 41608
rect 96160 41565 96169 41599
rect 96169 41565 96203 41599
rect 96203 41565 96212 41599
rect 96160 41556 96212 41565
rect 96528 41599 96580 41608
rect 96528 41565 96537 41599
rect 96537 41565 96571 41599
rect 96571 41565 96580 41599
rect 96528 41556 96580 41565
rect 18144 41488 18196 41540
rect 18788 41420 18840 41472
rect 80060 41420 80112 41472
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 65686 41318 65738 41370
rect 65750 41318 65802 41370
rect 65814 41318 65866 41370
rect 65878 41318 65930 41370
rect 96406 41318 96458 41370
rect 96470 41318 96522 41370
rect 96534 41318 96586 41370
rect 96598 41318 96650 41370
rect 12348 41216 12400 41268
rect 24860 41216 24912 41268
rect 44272 41216 44324 41268
rect 66904 41216 66956 41268
rect 25596 41148 25648 41200
rect 34428 41148 34480 41200
rect 44640 41148 44692 41200
rect 48136 41148 48188 41200
rect 14372 41080 14424 41132
rect 26976 41080 27028 41132
rect 8300 41012 8352 41064
rect 36544 41012 36596 41064
rect 14832 40944 14884 40996
rect 42524 40944 42576 40996
rect 86868 40944 86920 40996
rect 92112 40944 92164 40996
rect 11888 40876 11940 40928
rect 12348 40876 12400 40928
rect 24860 40876 24912 40928
rect 53748 40876 53800 40928
rect 66904 40876 66956 40928
rect 88432 40876 88484 40928
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 50326 40774 50378 40826
rect 50390 40774 50442 40826
rect 50454 40774 50506 40826
rect 50518 40774 50570 40826
rect 81046 40774 81098 40826
rect 81110 40774 81162 40826
rect 81174 40774 81226 40826
rect 81238 40774 81290 40826
rect 19984 40672 20036 40724
rect 68560 40672 68612 40724
rect 31760 40536 31812 40588
rect 32404 40536 32456 40588
rect 86408 40672 86460 40724
rect 86868 40672 86920 40724
rect 90548 40715 90600 40724
rect 90548 40681 90557 40715
rect 90557 40681 90591 40715
rect 90591 40681 90600 40715
rect 90548 40672 90600 40681
rect 95516 40715 95568 40724
rect 95516 40681 95525 40715
rect 95525 40681 95559 40715
rect 95559 40681 95568 40715
rect 95516 40672 95568 40681
rect 36360 40468 36412 40520
rect 36544 40468 36596 40520
rect 67732 40468 67784 40520
rect 68560 40468 68612 40520
rect 68928 40468 68980 40520
rect 34428 40400 34480 40452
rect 74080 40468 74132 40520
rect 92020 40468 92072 40520
rect 92388 40511 92440 40520
rect 92388 40477 92397 40511
rect 92397 40477 92431 40511
rect 92431 40477 92440 40511
rect 92388 40468 92440 40477
rect 66168 40332 66220 40384
rect 77668 40375 77720 40384
rect 77668 40341 77677 40375
rect 77677 40341 77711 40375
rect 77711 40341 77720 40375
rect 77668 40332 77720 40341
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 65686 40230 65738 40282
rect 65750 40230 65802 40282
rect 65814 40230 65866 40282
rect 65878 40230 65930 40282
rect 96406 40230 96458 40282
rect 96470 40230 96522 40282
rect 96534 40230 96586 40282
rect 96598 40230 96650 40282
rect 53656 40128 53708 40180
rect 77668 40128 77720 40180
rect 34244 40060 34296 40112
rect 35808 40060 35860 40112
rect 39764 40060 39816 40112
rect 43812 40060 43864 40112
rect 44824 40060 44876 40112
rect 47032 40060 47084 40112
rect 48964 40060 49016 40112
rect 67732 40060 67784 40112
rect 68652 40060 68704 40112
rect 12992 39992 13044 40044
rect 14648 39992 14700 40044
rect 10876 39924 10928 39976
rect 7748 39856 7800 39908
rect 10048 39856 10100 39908
rect 18972 39924 19024 39976
rect 28264 39788 28316 39840
rect 28724 39924 28776 39976
rect 34428 39967 34480 39976
rect 34428 39933 34437 39967
rect 34437 39933 34471 39967
rect 34471 39933 34480 39967
rect 34428 39924 34480 39933
rect 34612 39967 34664 39976
rect 34612 39933 34621 39967
rect 34621 39933 34655 39967
rect 34655 39933 34664 39967
rect 34612 39924 34664 39933
rect 35256 39924 35308 39976
rect 40776 39967 40828 39976
rect 40776 39933 40785 39967
rect 40785 39933 40819 39967
rect 40819 39933 40828 39967
rect 40776 39924 40828 39933
rect 31024 39856 31076 39908
rect 34704 39899 34756 39908
rect 34704 39865 34713 39899
rect 34713 39865 34747 39899
rect 34747 39865 34756 39899
rect 34704 39856 34756 39865
rect 49700 39992 49752 40044
rect 50068 40035 50120 40044
rect 50068 40001 50077 40035
rect 50077 40001 50111 40035
rect 50111 40001 50120 40035
rect 50068 39992 50120 40001
rect 60924 40035 60976 40044
rect 41604 39967 41656 39976
rect 41052 39856 41104 39908
rect 29736 39831 29788 39840
rect 29736 39797 29745 39831
rect 29745 39797 29779 39831
rect 29779 39797 29788 39831
rect 29736 39788 29788 39797
rect 32864 39788 32916 39840
rect 34060 39788 34112 39840
rect 34796 39788 34848 39840
rect 40592 39831 40644 39840
rect 40592 39797 40601 39831
rect 40601 39797 40635 39831
rect 40635 39797 40644 39831
rect 40592 39788 40644 39797
rect 41604 39933 41613 39967
rect 41613 39933 41647 39967
rect 41647 39933 41656 39967
rect 41604 39924 41656 39933
rect 44824 39924 44876 39976
rect 45192 39924 45244 39976
rect 57336 39924 57388 39976
rect 60924 40001 60933 40035
rect 60933 40001 60967 40035
rect 60967 40001 60976 40035
rect 60924 39992 60976 40001
rect 73620 39992 73672 40044
rect 61568 39924 61620 39976
rect 71504 39924 71556 39976
rect 72056 39967 72108 39976
rect 72056 39933 72065 39967
rect 72065 39933 72099 39967
rect 72099 39933 72108 39967
rect 72056 39924 72108 39933
rect 41236 39856 41288 39908
rect 44824 39788 44876 39840
rect 64052 39788 64104 39840
rect 73344 39856 73396 39908
rect 73160 39831 73212 39840
rect 73160 39797 73169 39831
rect 73169 39797 73203 39831
rect 73203 39797 73212 39831
rect 73160 39788 73212 39797
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 50326 39686 50378 39738
rect 50390 39686 50442 39738
rect 50454 39686 50506 39738
rect 50518 39686 50570 39738
rect 81046 39686 81098 39738
rect 81110 39686 81162 39738
rect 81174 39686 81226 39738
rect 81238 39686 81290 39738
rect 6184 39627 6236 39636
rect 6184 39593 6193 39627
rect 6193 39593 6227 39627
rect 6227 39593 6236 39627
rect 6184 39584 6236 39593
rect 28264 39584 28316 39636
rect 31116 39584 31168 39636
rect 33692 39584 33744 39636
rect 34152 39627 34204 39636
rect 34152 39593 34161 39627
rect 34161 39593 34195 39627
rect 34195 39593 34204 39627
rect 34152 39584 34204 39593
rect 40776 39584 40828 39636
rect 42064 39584 42116 39636
rect 49700 39584 49752 39636
rect 50988 39584 51040 39636
rect 70032 39584 70084 39636
rect 76840 39584 76892 39636
rect 5080 39491 5132 39500
rect 5080 39457 5089 39491
rect 5089 39457 5123 39491
rect 5123 39457 5132 39491
rect 5080 39448 5132 39457
rect 29552 39448 29604 39500
rect 31576 39448 31628 39500
rect 32956 39491 33008 39500
rect 6092 39380 6144 39432
rect 32496 39423 32548 39432
rect 32496 39389 32505 39423
rect 32505 39389 32539 39423
rect 32539 39389 32548 39423
rect 32496 39380 32548 39389
rect 32956 39457 32965 39491
rect 32965 39457 32999 39491
rect 32999 39457 33008 39491
rect 32956 39448 33008 39457
rect 33600 39491 33652 39500
rect 33600 39457 33609 39491
rect 33609 39457 33643 39491
rect 33643 39457 33652 39491
rect 33600 39448 33652 39457
rect 32864 39355 32916 39364
rect 32864 39321 32873 39355
rect 32873 39321 32907 39355
rect 32907 39321 32916 39355
rect 32864 39312 32916 39321
rect 24216 39244 24268 39296
rect 33508 39380 33560 39432
rect 33692 39423 33744 39432
rect 33692 39389 33701 39423
rect 33701 39389 33735 39423
rect 33735 39389 33744 39423
rect 33692 39380 33744 39389
rect 34060 39516 34112 39568
rect 44272 39516 44324 39568
rect 53748 39516 53800 39568
rect 78312 39516 78364 39568
rect 33968 39491 34020 39500
rect 33968 39457 33977 39491
rect 33977 39457 34011 39491
rect 34011 39457 34020 39491
rect 33968 39448 34020 39457
rect 34704 39448 34756 39500
rect 44916 39448 44968 39500
rect 55496 39448 55548 39500
rect 69020 39491 69072 39500
rect 69020 39457 69029 39491
rect 69029 39457 69063 39491
rect 69063 39457 69072 39491
rect 69020 39448 69072 39457
rect 63408 39380 63460 39432
rect 97448 39380 97500 39432
rect 35716 39244 35768 39296
rect 41236 39244 41288 39296
rect 69204 39312 69256 39364
rect 78404 39312 78456 39364
rect 66996 39244 67048 39296
rect 68928 39287 68980 39296
rect 68928 39253 68937 39287
rect 68937 39253 68971 39287
rect 68971 39253 68980 39287
rect 68928 39244 68980 39253
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 65686 39142 65738 39194
rect 65750 39142 65802 39194
rect 65814 39142 65866 39194
rect 65878 39142 65930 39194
rect 96406 39142 96458 39194
rect 96470 39142 96522 39194
rect 96534 39142 96586 39194
rect 96598 39142 96650 39194
rect 33508 39040 33560 39092
rect 34520 39040 34572 39092
rect 35532 39040 35584 39092
rect 40040 39040 40092 39092
rect 41144 39040 41196 39092
rect 68928 39040 68980 39092
rect 7564 38972 7616 39024
rect 40592 38972 40644 39024
rect 60372 38972 60424 39024
rect 73160 38972 73212 39024
rect 18236 38904 18288 38956
rect 18972 38904 19024 38956
rect 33600 38904 33652 38956
rect 33048 38811 33100 38820
rect 33048 38777 33057 38811
rect 33057 38777 33091 38811
rect 33091 38777 33100 38811
rect 33048 38768 33100 38777
rect 43536 38768 43588 38820
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 50326 38598 50378 38650
rect 50390 38598 50442 38650
rect 50454 38598 50506 38650
rect 50518 38598 50570 38650
rect 81046 38598 81098 38650
rect 81110 38598 81162 38650
rect 81174 38598 81226 38650
rect 81238 38598 81290 38650
rect 33048 38496 33100 38548
rect 43260 38496 43312 38548
rect 43352 38496 43404 38548
rect 94228 38496 94280 38548
rect 10508 38292 10560 38344
rect 10968 38360 11020 38412
rect 11336 38428 11388 38480
rect 16028 38360 16080 38412
rect 38108 38360 38160 38412
rect 42524 38403 42576 38412
rect 42524 38369 42533 38403
rect 42533 38369 42567 38403
rect 42567 38369 42576 38403
rect 42524 38360 42576 38369
rect 42892 38403 42944 38412
rect 20168 38292 20220 38344
rect 31024 38335 31076 38344
rect 31024 38301 31033 38335
rect 31033 38301 31067 38335
rect 31067 38301 31076 38335
rect 31024 38292 31076 38301
rect 31484 38292 31536 38344
rect 41328 38292 41380 38344
rect 42892 38369 42901 38403
rect 42901 38369 42935 38403
rect 42935 38369 42944 38403
rect 42892 38360 42944 38369
rect 43076 38403 43128 38412
rect 43076 38369 43085 38403
rect 43085 38369 43119 38403
rect 43119 38369 43128 38403
rect 43076 38360 43128 38369
rect 42984 38292 43036 38344
rect 11244 38224 11296 38276
rect 42524 38224 42576 38276
rect 46756 38360 46808 38412
rect 48136 38403 48188 38412
rect 48136 38369 48145 38403
rect 48145 38369 48179 38403
rect 48179 38369 48188 38403
rect 48136 38360 48188 38369
rect 48504 38360 48556 38412
rect 49608 38360 49660 38412
rect 73344 38428 73396 38480
rect 87604 38428 87656 38480
rect 72240 38292 72292 38344
rect 73068 38292 73120 38344
rect 48412 38224 48464 38276
rect 10876 38156 10928 38208
rect 24400 38156 24452 38208
rect 26240 38156 26292 38208
rect 34060 38199 34112 38208
rect 34060 38165 34069 38199
rect 34069 38165 34103 38199
rect 34103 38165 34112 38199
rect 34060 38156 34112 38165
rect 73528 38292 73580 38344
rect 74724 38335 74776 38344
rect 74724 38301 74733 38335
rect 74733 38301 74767 38335
rect 74767 38301 74776 38335
rect 74724 38292 74776 38301
rect 74448 38224 74500 38276
rect 91836 38224 91888 38276
rect 73620 38156 73672 38208
rect 77576 38156 77628 38208
rect 81164 38156 81216 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 65686 38054 65738 38106
rect 65750 38054 65802 38106
rect 65814 38054 65866 38106
rect 65878 38054 65930 38106
rect 96406 38054 96458 38106
rect 96470 38054 96522 38106
rect 96534 38054 96586 38106
rect 96598 38054 96650 38106
rect 11244 37952 11296 38004
rect 17684 37952 17736 38004
rect 17500 37884 17552 37936
rect 17868 37884 17920 37936
rect 26240 37952 26292 38004
rect 78404 37995 78456 38004
rect 42892 37884 42944 37936
rect 43352 37884 43404 37936
rect 47032 37927 47084 37936
rect 6092 37748 6144 37800
rect 6736 37748 6788 37800
rect 10968 37816 11020 37868
rect 46664 37859 46716 37868
rect 9404 37791 9456 37800
rect 9404 37757 9413 37791
rect 9413 37757 9447 37791
rect 9447 37757 9456 37791
rect 9404 37748 9456 37757
rect 12440 37748 12492 37800
rect 17040 37748 17092 37800
rect 17868 37748 17920 37800
rect 19892 37791 19944 37800
rect 19892 37757 19901 37791
rect 19901 37757 19935 37791
rect 19935 37757 19944 37791
rect 19892 37748 19944 37757
rect 26332 37791 26384 37800
rect 26332 37757 26341 37791
rect 26341 37757 26375 37791
rect 26375 37757 26384 37791
rect 26332 37748 26384 37757
rect 5448 37612 5500 37664
rect 46296 37791 46348 37800
rect 46296 37757 46305 37791
rect 46305 37757 46339 37791
rect 46339 37757 46348 37791
rect 46296 37748 46348 37757
rect 46664 37825 46673 37859
rect 46673 37825 46707 37859
rect 46707 37825 46716 37859
rect 46664 37816 46716 37825
rect 47032 37893 47041 37927
rect 47041 37893 47075 37927
rect 47075 37893 47084 37927
rect 47032 37884 47084 37893
rect 48412 37816 48464 37868
rect 46572 37791 46624 37800
rect 46572 37757 46581 37791
rect 46581 37757 46615 37791
rect 46615 37757 46624 37791
rect 46848 37791 46900 37800
rect 46572 37748 46624 37757
rect 43812 37680 43864 37732
rect 46848 37757 46857 37791
rect 46857 37757 46891 37791
rect 46891 37757 46900 37791
rect 46848 37748 46900 37757
rect 78404 37961 78413 37995
rect 78413 37961 78447 37995
rect 78447 37961 78456 37995
rect 78404 37952 78456 37961
rect 81164 37952 81216 38004
rect 89812 37952 89864 38004
rect 92388 37884 92440 37936
rect 78956 37859 79008 37868
rect 49516 37748 49568 37800
rect 50896 37791 50948 37800
rect 50896 37757 50905 37791
rect 50905 37757 50939 37791
rect 50939 37757 50948 37791
rect 50896 37748 50948 37757
rect 78588 37791 78640 37800
rect 57336 37680 57388 37732
rect 57704 37680 57756 37732
rect 18512 37612 18564 37664
rect 50160 37612 50212 37664
rect 50804 37655 50856 37664
rect 50804 37621 50813 37655
rect 50813 37621 50847 37655
rect 50847 37621 50856 37655
rect 50804 37612 50856 37621
rect 73528 37655 73580 37664
rect 73528 37621 73537 37655
rect 73537 37621 73571 37655
rect 73571 37621 73580 37655
rect 78588 37757 78597 37791
rect 78597 37757 78631 37791
rect 78631 37757 78640 37791
rect 78588 37748 78640 37757
rect 78956 37825 78965 37859
rect 78965 37825 78999 37859
rect 78999 37825 79008 37859
rect 78956 37816 79008 37825
rect 81164 37859 81216 37868
rect 81164 37825 81173 37859
rect 81173 37825 81207 37859
rect 81207 37825 81216 37859
rect 81164 37816 81216 37825
rect 87696 37859 87748 37868
rect 87696 37825 87705 37859
rect 87705 37825 87739 37859
rect 87739 37825 87748 37859
rect 87696 37816 87748 37825
rect 87788 37816 87840 37868
rect 78864 37791 78916 37800
rect 78864 37757 78873 37791
rect 78873 37757 78907 37791
rect 78907 37757 78916 37791
rect 79140 37791 79192 37800
rect 78864 37748 78916 37757
rect 79140 37757 79156 37791
rect 79156 37757 79192 37791
rect 79140 37748 79192 37757
rect 93860 37748 93912 37800
rect 87512 37723 87564 37732
rect 87512 37689 87521 37723
rect 87521 37689 87555 37723
rect 87555 37689 87564 37723
rect 87512 37680 87564 37689
rect 79232 37655 79284 37664
rect 73528 37612 73580 37621
rect 79232 37621 79241 37655
rect 79241 37621 79275 37655
rect 79275 37621 79284 37655
rect 79232 37612 79284 37621
rect 82544 37655 82596 37664
rect 82544 37621 82553 37655
rect 82553 37621 82587 37655
rect 82587 37621 82596 37655
rect 89628 37680 89680 37732
rect 82544 37612 82596 37621
rect 92664 37612 92716 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 50326 37510 50378 37562
rect 50390 37510 50442 37562
rect 50454 37510 50506 37562
rect 50518 37510 50570 37562
rect 81046 37510 81098 37562
rect 81110 37510 81162 37562
rect 81174 37510 81226 37562
rect 81238 37510 81290 37562
rect 17960 37408 18012 37460
rect 12992 37340 13044 37392
rect 11244 37315 11296 37324
rect 11244 37281 11253 37315
rect 11253 37281 11287 37315
rect 11287 37281 11296 37315
rect 11244 37272 11296 37281
rect 11520 37315 11572 37324
rect 11520 37281 11529 37315
rect 11529 37281 11563 37315
rect 11563 37281 11572 37315
rect 11520 37272 11572 37281
rect 17776 37315 17828 37324
rect 17776 37281 17785 37315
rect 17785 37281 17819 37315
rect 17819 37281 17828 37315
rect 17776 37272 17828 37281
rect 20720 37408 20772 37460
rect 20996 37408 21048 37460
rect 52368 37408 52420 37460
rect 18512 37340 18564 37392
rect 18604 37315 18656 37324
rect 18604 37281 18613 37315
rect 18613 37281 18647 37315
rect 18647 37281 18656 37315
rect 18604 37272 18656 37281
rect 36176 37340 36228 37392
rect 19984 37272 20036 37324
rect 73252 37340 73304 37392
rect 74080 37272 74132 37324
rect 74540 37315 74592 37324
rect 18512 37204 18564 37256
rect 74540 37281 74549 37315
rect 74549 37281 74583 37315
rect 74583 37281 74592 37315
rect 74540 37272 74592 37281
rect 74448 37247 74500 37256
rect 74448 37213 74457 37247
rect 74457 37213 74491 37247
rect 74491 37213 74500 37247
rect 74448 37204 74500 37213
rect 76380 37272 76432 37324
rect 79692 37272 79744 37324
rect 87512 37408 87564 37460
rect 87972 37408 88024 37460
rect 94228 37315 94280 37324
rect 94228 37281 94237 37315
rect 94237 37281 94271 37315
rect 94271 37281 94280 37315
rect 94228 37272 94280 37281
rect 78036 37204 78088 37256
rect 93032 37136 93084 37188
rect 83648 37068 83700 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 65686 36966 65738 37018
rect 65750 36966 65802 37018
rect 65814 36966 65866 37018
rect 65878 36966 65930 37018
rect 96406 36966 96458 37018
rect 96470 36966 96522 37018
rect 96534 36966 96586 37018
rect 96598 36966 96650 37018
rect 3332 36907 3384 36916
rect 3332 36873 3341 36907
rect 3341 36873 3375 36907
rect 3375 36873 3384 36907
rect 3332 36864 3384 36873
rect 49608 36864 49660 36916
rect 76196 36907 76248 36916
rect 33692 36796 33744 36848
rect 63316 36796 63368 36848
rect 76196 36873 76205 36907
rect 76205 36873 76239 36907
rect 76239 36873 76248 36907
rect 76196 36864 76248 36873
rect 6000 36728 6052 36780
rect 9956 36728 10008 36780
rect 52368 36728 52420 36780
rect 57336 36728 57388 36780
rect 89260 36728 89312 36780
rect 8208 36660 8260 36712
rect 16028 36660 16080 36712
rect 49608 36660 49660 36712
rect 75000 36703 75052 36712
rect 75000 36669 75009 36703
rect 75009 36669 75043 36703
rect 75043 36669 75052 36703
rect 75000 36660 75052 36669
rect 75184 36703 75236 36712
rect 75184 36669 75193 36703
rect 75193 36669 75227 36703
rect 75227 36669 75236 36703
rect 75184 36660 75236 36669
rect 75368 36703 75420 36712
rect 75368 36669 75377 36703
rect 75377 36669 75411 36703
rect 75411 36669 75420 36703
rect 75368 36660 75420 36669
rect 75736 36703 75788 36712
rect 75736 36669 75745 36703
rect 75745 36669 75779 36703
rect 75779 36669 75788 36703
rect 75736 36660 75788 36669
rect 75828 36660 75880 36712
rect 6460 36592 6512 36644
rect 19432 36592 19484 36644
rect 20628 36592 20680 36644
rect 48412 36592 48464 36644
rect 88432 36703 88484 36712
rect 88432 36669 88441 36703
rect 88441 36669 88475 36703
rect 88475 36669 88484 36703
rect 88432 36660 88484 36669
rect 8576 36524 8628 36576
rect 59268 36524 59320 36576
rect 88432 36567 88484 36576
rect 88432 36533 88441 36567
rect 88441 36533 88475 36567
rect 88475 36533 88484 36567
rect 88432 36524 88484 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 50326 36422 50378 36474
rect 50390 36422 50442 36474
rect 50454 36422 50506 36474
rect 50518 36422 50570 36474
rect 81046 36422 81098 36474
rect 81110 36422 81162 36474
rect 81174 36422 81226 36474
rect 81238 36422 81290 36474
rect 20628 36320 20680 36372
rect 51356 36320 51408 36372
rect 51448 36320 51500 36372
rect 66812 36320 66864 36372
rect 40868 36252 40920 36304
rect 41328 36252 41380 36304
rect 35808 36227 35860 36236
rect 35808 36193 35817 36227
rect 35817 36193 35851 36227
rect 35851 36193 35860 36227
rect 35808 36184 35860 36193
rect 42064 36184 42116 36236
rect 51448 36227 51500 36236
rect 51448 36193 51457 36227
rect 51457 36193 51491 36227
rect 51491 36193 51500 36227
rect 51448 36184 51500 36193
rect 51632 36227 51684 36236
rect 51632 36193 51640 36227
rect 51640 36193 51674 36227
rect 51674 36193 51684 36227
rect 51816 36227 51868 36236
rect 51632 36184 51684 36193
rect 51816 36193 51825 36227
rect 51825 36193 51859 36227
rect 51859 36193 51868 36227
rect 51816 36184 51868 36193
rect 52184 36227 52236 36236
rect 52184 36193 52193 36227
rect 52193 36193 52227 36227
rect 52227 36193 52236 36227
rect 52184 36184 52236 36193
rect 63040 36227 63092 36236
rect 63040 36193 63049 36227
rect 63049 36193 63083 36227
rect 63083 36193 63092 36227
rect 63040 36184 63092 36193
rect 63592 36227 63644 36236
rect 63592 36193 63601 36227
rect 63601 36193 63635 36227
rect 63635 36193 63644 36227
rect 63592 36184 63644 36193
rect 64696 36184 64748 36236
rect 75736 36320 75788 36372
rect 76012 36320 76064 36372
rect 76932 36320 76984 36372
rect 75368 36252 75420 36304
rect 75920 36252 75972 36304
rect 76748 36252 76800 36304
rect 20720 36116 20772 36168
rect 39764 36116 39816 36168
rect 51724 36159 51776 36168
rect 51724 36125 51733 36159
rect 51733 36125 51767 36159
rect 51767 36125 51776 36159
rect 51724 36116 51776 36125
rect 51908 36116 51960 36168
rect 63316 36159 63368 36168
rect 63316 36125 63325 36159
rect 63325 36125 63359 36159
rect 63359 36125 63368 36159
rect 63316 36116 63368 36125
rect 63408 36159 63460 36168
rect 63408 36125 63417 36159
rect 63417 36125 63451 36159
rect 63451 36125 63460 36159
rect 63408 36116 63460 36125
rect 74264 36116 74316 36168
rect 77944 36159 77996 36168
rect 77944 36125 77953 36159
rect 77953 36125 77987 36159
rect 77987 36125 77996 36159
rect 77944 36116 77996 36125
rect 23572 36048 23624 36100
rect 78312 36227 78364 36236
rect 78312 36193 78321 36227
rect 78321 36193 78355 36227
rect 78355 36193 78364 36227
rect 78312 36184 78364 36193
rect 63684 36023 63736 36032
rect 63684 35989 63693 36023
rect 63693 35989 63727 36023
rect 63727 35989 63736 36023
rect 63684 35980 63736 35989
rect 70308 35980 70360 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 65686 35878 65738 35930
rect 65750 35878 65802 35930
rect 65814 35878 65866 35930
rect 65878 35878 65930 35930
rect 96406 35878 96458 35930
rect 96470 35878 96522 35930
rect 96534 35878 96586 35930
rect 96598 35878 96650 35930
rect 57336 35776 57388 35828
rect 57612 35776 57664 35828
rect 73436 35776 73488 35828
rect 73988 35776 74040 35828
rect 11796 35572 11848 35624
rect 73804 35572 73856 35624
rect 23940 35504 23992 35556
rect 36268 35504 36320 35556
rect 9036 35436 9088 35488
rect 31484 35436 31536 35488
rect 73896 35436 73948 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 50326 35334 50378 35386
rect 50390 35334 50442 35386
rect 50454 35334 50506 35386
rect 50518 35334 50570 35386
rect 81046 35334 81098 35386
rect 81110 35334 81162 35386
rect 81174 35334 81226 35386
rect 81238 35334 81290 35386
rect 10048 35232 10100 35284
rect 40040 35232 40092 35284
rect 42800 35164 42852 35216
rect 51724 35164 51776 35216
rect 39856 35096 39908 35148
rect 63408 35096 63460 35148
rect 31024 35028 31076 35080
rect 31392 35028 31444 35080
rect 66260 34960 66312 35012
rect 66904 34960 66956 35012
rect 73804 34960 73856 35012
rect 29000 34935 29052 34944
rect 29000 34901 29009 34935
rect 29009 34901 29043 34935
rect 29043 34901 29052 34935
rect 29000 34892 29052 34901
rect 65432 34892 65484 34944
rect 66444 34892 66496 34944
rect 72332 34892 72384 34944
rect 84384 34892 84436 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 65686 34790 65738 34842
rect 65750 34790 65802 34842
rect 65814 34790 65866 34842
rect 65878 34790 65930 34842
rect 96406 34790 96458 34842
rect 96470 34790 96522 34842
rect 96534 34790 96586 34842
rect 96598 34790 96650 34842
rect 29000 34688 29052 34740
rect 53564 34688 53616 34740
rect 54668 34688 54720 34740
rect 57336 34688 57388 34740
rect 51816 34620 51868 34672
rect 65432 34620 65484 34672
rect 66444 34688 66496 34740
rect 70308 34688 70360 34740
rect 66628 34620 66680 34672
rect 66904 34663 66956 34672
rect 66904 34629 66913 34663
rect 66913 34629 66947 34663
rect 66947 34629 66956 34663
rect 66904 34620 66956 34629
rect 43536 34552 43588 34604
rect 48044 34552 48096 34604
rect 51724 34552 51776 34604
rect 74264 34552 74316 34604
rect 19892 34484 19944 34536
rect 25688 34484 25740 34536
rect 33324 34484 33376 34536
rect 66260 34527 66312 34536
rect 66260 34493 66269 34527
rect 66269 34493 66303 34527
rect 66303 34493 66312 34527
rect 66260 34484 66312 34493
rect 66444 34527 66496 34536
rect 66444 34493 66453 34527
rect 66453 34493 66487 34527
rect 66487 34493 66496 34527
rect 66444 34484 66496 34493
rect 66628 34527 66680 34536
rect 66628 34493 66638 34527
rect 66638 34493 66672 34527
rect 66672 34493 66680 34527
rect 66628 34484 66680 34493
rect 66904 34484 66956 34536
rect 67824 34527 67876 34536
rect 67824 34493 67833 34527
rect 67833 34493 67867 34527
rect 67867 34493 67876 34527
rect 67824 34484 67876 34493
rect 73436 34484 73488 34536
rect 26516 34416 26568 34468
rect 30380 34416 30432 34468
rect 41604 34416 41656 34468
rect 65432 34416 65484 34468
rect 35256 34348 35308 34400
rect 65616 34348 65668 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 50326 34246 50378 34298
rect 50390 34246 50442 34298
rect 50454 34246 50506 34298
rect 50518 34246 50570 34298
rect 81046 34246 81098 34298
rect 81110 34246 81162 34298
rect 81174 34246 81226 34298
rect 81238 34246 81290 34298
rect 3516 34144 3568 34196
rect 44180 34144 44232 34196
rect 56600 34187 56652 34196
rect 56600 34153 56609 34187
rect 56609 34153 56643 34187
rect 56643 34153 56652 34187
rect 56600 34144 56652 34153
rect 65432 34144 65484 34196
rect 73252 34144 73304 34196
rect 21732 34076 21784 34128
rect 17684 34008 17736 34060
rect 39948 34076 40000 34128
rect 64144 34076 64196 34128
rect 90732 34076 90784 34128
rect 31116 33872 31168 33924
rect 44548 33940 44600 33992
rect 57060 34051 57112 34060
rect 57060 34017 57069 34051
rect 57069 34017 57103 34051
rect 57103 34017 57112 34051
rect 57060 34008 57112 34017
rect 62948 34008 63000 34060
rect 63408 34008 63460 34060
rect 65616 34008 65668 34060
rect 74448 34008 74500 34060
rect 56968 33983 57020 33992
rect 56968 33949 56977 33983
rect 56977 33949 57011 33983
rect 57011 33949 57020 33983
rect 56968 33940 57020 33949
rect 57796 33940 57848 33992
rect 92940 33940 92992 33992
rect 33048 33804 33100 33856
rect 34520 33804 34572 33856
rect 67824 33872 67876 33924
rect 40960 33804 41012 33856
rect 57428 33847 57480 33856
rect 57428 33813 57437 33847
rect 57437 33813 57471 33847
rect 57471 33813 57480 33847
rect 57428 33804 57480 33813
rect 95792 33804 95844 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 65686 33702 65738 33754
rect 65750 33702 65802 33754
rect 65814 33702 65866 33754
rect 65878 33702 65930 33754
rect 96406 33702 96458 33754
rect 96470 33702 96522 33754
rect 96534 33702 96586 33754
rect 96598 33702 96650 33754
rect 10876 33600 10928 33652
rect 90824 33600 90876 33652
rect 65432 33532 65484 33584
rect 66168 33532 66220 33584
rect 9588 33464 9640 33516
rect 56968 33464 57020 33516
rect 31024 33396 31076 33448
rect 33048 33439 33100 33448
rect 33048 33405 33057 33439
rect 33057 33405 33091 33439
rect 33091 33405 33100 33439
rect 33048 33396 33100 33405
rect 33324 33439 33376 33448
rect 33324 33405 33333 33439
rect 33333 33405 33367 33439
rect 33367 33405 33376 33439
rect 33324 33396 33376 33405
rect 97540 33396 97592 33448
rect 31208 33260 31260 33312
rect 66260 33260 66312 33312
rect 66904 33260 66956 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 50326 33158 50378 33210
rect 50390 33158 50442 33210
rect 50454 33158 50506 33210
rect 50518 33158 50570 33210
rect 81046 33158 81098 33210
rect 81110 33158 81162 33210
rect 81174 33158 81226 33210
rect 81238 33158 81290 33210
rect 31944 33056 31996 33108
rect 40776 33056 40828 33108
rect 70952 33056 71004 33108
rect 71320 33056 71372 33108
rect 58900 33031 58952 33040
rect 58900 32997 58909 33031
rect 58909 32997 58943 33031
rect 58943 32997 58952 33031
rect 58900 32988 58952 32997
rect 58072 32963 58124 32972
rect 58072 32929 58081 32963
rect 58081 32929 58115 32963
rect 58115 32929 58124 32963
rect 58072 32920 58124 32929
rect 14004 32784 14056 32836
rect 34152 32784 34204 32836
rect 56048 32716 56100 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 65686 32614 65738 32666
rect 65750 32614 65802 32666
rect 65814 32614 65866 32666
rect 65878 32614 65930 32666
rect 96406 32614 96458 32666
rect 96470 32614 96522 32666
rect 96534 32614 96586 32666
rect 96598 32614 96650 32666
rect 9036 32512 9088 32564
rect 16212 32512 16264 32564
rect 30288 32512 30340 32564
rect 24124 32444 24176 32496
rect 92388 32487 92440 32496
rect 92388 32453 92397 32487
rect 92397 32453 92431 32487
rect 92431 32453 92440 32487
rect 92388 32444 92440 32453
rect 3056 32351 3108 32360
rect 3056 32317 3065 32351
rect 3065 32317 3099 32351
rect 3099 32317 3108 32351
rect 3056 32308 3108 32317
rect 6368 32376 6420 32428
rect 43536 32376 43588 32428
rect 47308 32376 47360 32428
rect 67088 32376 67140 32428
rect 92480 32419 92532 32428
rect 92480 32385 92489 32419
rect 92489 32385 92523 32419
rect 92523 32385 92532 32419
rect 92480 32376 92532 32385
rect 6736 32308 6788 32360
rect 12164 32308 12216 32360
rect 30748 32308 30800 32360
rect 95056 32308 95108 32360
rect 83740 32240 83792 32292
rect 4344 32215 4396 32224
rect 4344 32181 4353 32215
rect 4353 32181 4387 32215
rect 4387 32181 4396 32215
rect 4344 32172 4396 32181
rect 41788 32172 41840 32224
rect 45008 32172 45060 32224
rect 73068 32172 73120 32224
rect 88984 32172 89036 32224
rect 92756 32215 92808 32224
rect 92756 32181 92765 32215
rect 92765 32181 92799 32215
rect 92799 32181 92808 32215
rect 92756 32172 92808 32181
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 50326 32070 50378 32122
rect 50390 32070 50442 32122
rect 50454 32070 50506 32122
rect 50518 32070 50570 32122
rect 81046 32070 81098 32122
rect 81110 32070 81162 32122
rect 81174 32070 81226 32122
rect 81238 32070 81290 32122
rect 4344 31968 4396 32020
rect 12348 31968 12400 32020
rect 85028 31968 85080 32020
rect 95056 32011 95108 32020
rect 69848 31900 69900 31952
rect 70216 31900 70268 31952
rect 40776 31832 40828 31884
rect 88984 31832 89036 31884
rect 94044 31900 94096 31952
rect 95056 31977 95065 32011
rect 95065 31977 95099 32011
rect 95099 31977 95108 32011
rect 95056 31968 95108 31977
rect 39948 31764 40000 31816
rect 43076 31807 43128 31816
rect 43076 31773 43085 31807
rect 43085 31773 43119 31807
rect 43119 31773 43128 31807
rect 43076 31764 43128 31773
rect 43352 31807 43404 31816
rect 43352 31773 43361 31807
rect 43361 31773 43395 31807
rect 43395 31773 43404 31807
rect 43352 31764 43404 31773
rect 71320 31764 71372 31816
rect 92664 31764 92716 31816
rect 63960 31628 64012 31680
rect 69480 31628 69532 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 65686 31526 65738 31578
rect 65750 31526 65802 31578
rect 65814 31526 65866 31578
rect 65878 31526 65930 31578
rect 96406 31526 96458 31578
rect 96470 31526 96522 31578
rect 96534 31526 96586 31578
rect 96598 31526 96650 31578
rect 64604 31467 64656 31476
rect 64604 31433 64613 31467
rect 64613 31433 64647 31467
rect 64647 31433 64656 31467
rect 64604 31424 64656 31433
rect 67824 31424 67876 31476
rect 64144 31356 64196 31408
rect 70032 31356 70084 31408
rect 53840 31288 53892 31340
rect 64328 31288 64380 31340
rect 68652 31288 68704 31340
rect 77852 31288 77904 31340
rect 48136 31220 48188 31272
rect 34796 31152 34848 31204
rect 64144 31152 64196 31204
rect 71596 31263 71648 31272
rect 71596 31229 71605 31263
rect 71605 31229 71639 31263
rect 71639 31229 71648 31263
rect 71596 31220 71648 31229
rect 81532 31220 81584 31272
rect 24216 31084 24268 31136
rect 33416 31084 33468 31136
rect 63960 31084 64012 31136
rect 64052 31084 64104 31136
rect 64604 31084 64656 31136
rect 67088 31084 67140 31136
rect 68744 31084 68796 31136
rect 71412 31127 71464 31136
rect 71412 31093 71421 31127
rect 71421 31093 71455 31127
rect 71455 31093 71464 31127
rect 71412 31084 71464 31093
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 50326 30982 50378 31034
rect 50390 30982 50442 31034
rect 50454 30982 50506 31034
rect 50518 30982 50570 31034
rect 81046 30982 81098 31034
rect 81110 30982 81162 31034
rect 81174 30982 81226 31034
rect 81238 30982 81290 31034
rect 26516 30880 26568 30932
rect 30012 30880 30064 30932
rect 31116 30880 31168 30932
rect 31300 30880 31352 30932
rect 9956 30787 10008 30796
rect 9956 30753 9965 30787
rect 9965 30753 9999 30787
rect 9999 30753 10008 30787
rect 9956 30744 10008 30753
rect 11888 30812 11940 30864
rect 32220 30812 32272 30864
rect 67916 30812 67968 30864
rect 10600 30744 10652 30796
rect 15200 30744 15252 30796
rect 64328 30744 64380 30796
rect 67824 30787 67876 30796
rect 67824 30753 67833 30787
rect 67833 30753 67867 30787
rect 67867 30753 67876 30787
rect 84844 30880 84896 30932
rect 69480 30855 69532 30864
rect 69480 30821 69489 30855
rect 69489 30821 69523 30855
rect 69523 30821 69532 30855
rect 69480 30812 69532 30821
rect 67824 30744 67876 30753
rect 68652 30744 68704 30796
rect 69664 30787 69716 30796
rect 69664 30753 69673 30787
rect 69673 30753 69707 30787
rect 69707 30753 69716 30787
rect 69664 30744 69716 30753
rect 70032 30787 70084 30796
rect 70032 30753 70041 30787
rect 70041 30753 70075 30787
rect 70075 30753 70084 30787
rect 70032 30744 70084 30753
rect 21364 30676 21416 30728
rect 22284 30676 22336 30728
rect 2872 30608 2924 30660
rect 9772 30651 9824 30660
rect 9772 30617 9781 30651
rect 9781 30617 9815 30651
rect 9815 30617 9824 30651
rect 9772 30608 9824 30617
rect 68744 30676 68796 30728
rect 70492 30744 70544 30796
rect 92388 30676 92440 30728
rect 67088 30583 67140 30592
rect 67088 30549 67097 30583
rect 67097 30549 67131 30583
rect 67131 30549 67140 30583
rect 67088 30540 67140 30549
rect 70032 30540 70084 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 65686 30438 65738 30490
rect 65750 30438 65802 30490
rect 65814 30438 65866 30490
rect 65878 30438 65930 30490
rect 96406 30438 96458 30490
rect 96470 30438 96522 30490
rect 96534 30438 96586 30490
rect 96598 30438 96650 30490
rect 20076 30336 20128 30388
rect 67824 30336 67876 30388
rect 67916 30336 67968 30388
rect 70032 30336 70084 30388
rect 81532 30336 81584 30388
rect 82360 30336 82412 30388
rect 84568 30336 84620 30388
rect 84844 30336 84896 30388
rect 34520 30268 34572 30320
rect 43076 30268 43128 30320
rect 43720 30268 43772 30320
rect 25780 30200 25832 30252
rect 77760 30200 77812 30252
rect 78496 30243 78548 30252
rect 78496 30209 78505 30243
rect 78505 30209 78539 30243
rect 78539 30209 78548 30243
rect 78496 30200 78548 30209
rect 26056 30132 26108 30184
rect 41236 30175 41288 30184
rect 41236 30141 41245 30175
rect 41245 30141 41279 30175
rect 41279 30141 41288 30175
rect 41236 30132 41288 30141
rect 58164 30132 58216 30184
rect 26700 29996 26752 30048
rect 36544 29996 36596 30048
rect 41052 29996 41104 30048
rect 69756 30064 69808 30116
rect 86224 30132 86276 30184
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 50326 29894 50378 29946
rect 50390 29894 50442 29946
rect 50454 29894 50506 29946
rect 50518 29894 50570 29946
rect 81046 29894 81098 29946
rect 81110 29894 81162 29946
rect 81174 29894 81226 29946
rect 81238 29894 81290 29946
rect 40040 29792 40092 29844
rect 40500 29792 40552 29844
rect 46296 29792 46348 29844
rect 87512 29792 87564 29844
rect 88064 29792 88116 29844
rect 21272 29767 21324 29776
rect 21272 29733 21281 29767
rect 21281 29733 21315 29767
rect 21315 29733 21324 29767
rect 21272 29724 21324 29733
rect 26148 29724 26200 29776
rect 48320 29724 48372 29776
rect 84936 29724 84988 29776
rect 16212 29656 16264 29708
rect 21916 29699 21968 29708
rect 21916 29665 21925 29699
rect 21925 29665 21959 29699
rect 21959 29665 21968 29699
rect 21916 29656 21968 29665
rect 26792 29699 26844 29708
rect 26792 29665 26801 29699
rect 26801 29665 26835 29699
rect 26835 29665 26844 29699
rect 26792 29656 26844 29665
rect 27804 29656 27856 29708
rect 27988 29656 28040 29708
rect 34704 29588 34756 29640
rect 34796 29588 34848 29640
rect 46664 29588 46716 29640
rect 26424 29520 26476 29572
rect 22192 29495 22244 29504
rect 22192 29461 22201 29495
rect 22201 29461 22235 29495
rect 22235 29461 22244 29495
rect 22192 29452 22244 29461
rect 22284 29452 22336 29504
rect 45008 29520 45060 29572
rect 46296 29520 46348 29572
rect 88064 29588 88116 29640
rect 89260 29631 89312 29640
rect 89260 29597 89269 29631
rect 89269 29597 89303 29631
rect 89303 29597 89312 29631
rect 89260 29588 89312 29597
rect 96160 29588 96212 29640
rect 46572 29452 46624 29504
rect 84108 29452 84160 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 65686 29350 65738 29402
rect 65750 29350 65802 29402
rect 65814 29350 65866 29402
rect 65878 29350 65930 29402
rect 96406 29350 96458 29402
rect 96470 29350 96522 29402
rect 96534 29350 96586 29402
rect 96598 29350 96650 29402
rect 17684 29248 17736 29300
rect 25780 29248 25832 29300
rect 26240 29248 26292 29300
rect 26424 29248 26476 29300
rect 26792 29248 26844 29300
rect 22192 29180 22244 29232
rect 36544 29248 36596 29300
rect 45008 29248 45060 29300
rect 45100 29248 45152 29300
rect 46848 29248 46900 29300
rect 35348 29112 35400 29164
rect 40132 29180 40184 29232
rect 41236 29112 41288 29164
rect 78772 29248 78824 29300
rect 89260 29248 89312 29300
rect 90640 29248 90692 29300
rect 66996 29180 67048 29232
rect 22284 29044 22336 29096
rect 16212 28976 16264 29028
rect 16488 28976 16540 29028
rect 25688 28976 25740 29028
rect 26056 29087 26108 29096
rect 26056 29053 26065 29087
rect 26065 29053 26099 29087
rect 26099 29053 26108 29087
rect 26056 29044 26108 29053
rect 26240 29044 26292 29096
rect 26516 29087 26568 29096
rect 26516 29053 26525 29087
rect 26525 29053 26559 29087
rect 26559 29053 26568 29087
rect 26516 29044 26568 29053
rect 26700 29087 26752 29096
rect 26700 29053 26709 29087
rect 26709 29053 26743 29087
rect 26743 29053 26752 29087
rect 26700 29044 26752 29053
rect 43720 29044 43772 29096
rect 46848 29044 46900 29096
rect 78220 29112 78272 29164
rect 75092 29087 75144 29096
rect 75092 29053 75101 29087
rect 75101 29053 75135 29087
rect 75135 29053 75144 29087
rect 75092 29044 75144 29053
rect 34796 28976 34848 29028
rect 26056 28908 26108 28960
rect 40040 28908 40092 28960
rect 63960 28908 64012 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 50326 28806 50378 28858
rect 50390 28806 50442 28858
rect 50454 28806 50506 28858
rect 50518 28806 50570 28858
rect 81046 28806 81098 28858
rect 81110 28806 81162 28858
rect 81174 28806 81226 28858
rect 81238 28806 81290 28858
rect 53472 28704 53524 28756
rect 23204 28636 23256 28688
rect 40132 28636 40184 28688
rect 63500 28679 63552 28688
rect 15476 28568 15528 28620
rect 15660 28611 15712 28620
rect 15660 28577 15669 28611
rect 15669 28577 15703 28611
rect 15703 28577 15712 28611
rect 15660 28568 15712 28577
rect 60740 28568 60792 28620
rect 61292 28568 61344 28620
rect 63500 28645 63509 28679
rect 63509 28645 63543 28679
rect 63543 28645 63552 28679
rect 63500 28636 63552 28645
rect 63960 28679 64012 28688
rect 63960 28645 63969 28679
rect 63969 28645 64003 28679
rect 64003 28645 64012 28679
rect 63960 28636 64012 28645
rect 91928 28636 91980 28688
rect 77668 28611 77720 28620
rect 60648 28543 60700 28552
rect 60648 28509 60657 28543
rect 60657 28509 60691 28543
rect 60691 28509 60700 28543
rect 60648 28500 60700 28509
rect 77668 28577 77677 28611
rect 77677 28577 77711 28611
rect 77711 28577 77720 28611
rect 77668 28568 77720 28577
rect 77944 28543 77996 28552
rect 77944 28509 77953 28543
rect 77953 28509 77987 28543
rect 77987 28509 77996 28543
rect 77944 28500 77996 28509
rect 17868 28364 17920 28416
rect 21364 28364 21416 28416
rect 44640 28364 44692 28416
rect 84936 28432 84988 28484
rect 77668 28364 77720 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 65686 28262 65738 28314
rect 65750 28262 65802 28314
rect 65814 28262 65866 28314
rect 65878 28262 65930 28314
rect 96406 28262 96458 28314
rect 96470 28262 96522 28314
rect 96534 28262 96586 28314
rect 96598 28262 96650 28314
rect 8208 27956 8260 28008
rect 44180 28160 44232 28212
rect 9404 27888 9456 27940
rect 43720 27956 43772 28008
rect 43996 27999 44048 28008
rect 43996 27965 44005 27999
rect 44005 27965 44039 27999
rect 44039 27965 44048 27999
rect 43996 27956 44048 27965
rect 44180 27999 44232 28008
rect 44180 27965 44189 27999
rect 44189 27965 44223 27999
rect 44223 27965 44232 27999
rect 44180 27956 44232 27965
rect 44548 27999 44600 28008
rect 44272 27888 44324 27940
rect 44548 27965 44557 27999
rect 44557 27965 44591 27999
rect 44591 27965 44600 27999
rect 44548 27956 44600 27965
rect 77944 28160 77996 28212
rect 91652 28160 91704 28212
rect 95976 28160 96028 28212
rect 83188 28092 83240 28144
rect 55956 28067 56008 28076
rect 55956 28033 55965 28067
rect 55965 28033 55999 28067
rect 55999 28033 56008 28067
rect 55956 28024 56008 28033
rect 49424 27956 49476 28008
rect 55772 27999 55824 28008
rect 55772 27965 55780 27999
rect 55780 27965 55814 27999
rect 55814 27965 55824 27999
rect 55772 27956 55824 27965
rect 74632 28024 74684 28076
rect 56232 27956 56284 28008
rect 83464 27956 83516 28008
rect 8116 27820 8168 27872
rect 44548 27820 44600 27872
rect 60648 27888 60700 27940
rect 56232 27863 56284 27872
rect 56232 27829 56241 27863
rect 56241 27829 56275 27863
rect 56275 27829 56284 27863
rect 56232 27820 56284 27829
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 50326 27718 50378 27770
rect 50390 27718 50442 27770
rect 50454 27718 50506 27770
rect 50518 27718 50570 27770
rect 81046 27718 81098 27770
rect 81110 27718 81162 27770
rect 81174 27718 81226 27770
rect 81238 27718 81290 27770
rect 2412 27616 2464 27668
rect 7472 27616 7524 27668
rect 8208 27616 8260 27668
rect 28632 27616 28684 27668
rect 28908 27616 28960 27668
rect 43720 27616 43772 27668
rect 56232 27616 56284 27668
rect 88800 27616 88852 27668
rect 16028 27548 16080 27600
rect 90180 27548 90232 27600
rect 12808 27523 12860 27532
rect 12808 27489 12817 27523
rect 12817 27489 12851 27523
rect 12851 27489 12860 27523
rect 12808 27480 12860 27489
rect 15476 27480 15528 27532
rect 17132 27480 17184 27532
rect 21732 27480 21784 27532
rect 42064 27480 42116 27532
rect 42800 27523 42852 27532
rect 42800 27489 42809 27523
rect 42809 27489 42843 27523
rect 42843 27489 42852 27523
rect 42800 27480 42852 27489
rect 42892 27480 42944 27532
rect 51908 27480 51960 27532
rect 73344 27480 73396 27532
rect 74448 27480 74500 27532
rect 89628 27480 89680 27532
rect 14924 27455 14976 27464
rect 14924 27421 14933 27455
rect 14933 27421 14967 27455
rect 14967 27421 14976 27455
rect 14924 27412 14976 27421
rect 25412 27455 25464 27464
rect 25412 27421 25421 27455
rect 25421 27421 25455 27455
rect 25455 27421 25464 27455
rect 25412 27412 25464 27421
rect 42708 27455 42760 27464
rect 42708 27421 42717 27455
rect 42717 27421 42751 27455
rect 42751 27421 42760 27455
rect 42708 27412 42760 27421
rect 42984 27412 43036 27464
rect 43536 27455 43588 27464
rect 43536 27421 43545 27455
rect 43545 27421 43579 27455
rect 43579 27421 43588 27455
rect 43536 27412 43588 27421
rect 46112 27412 46164 27464
rect 60188 27412 60240 27464
rect 60280 27344 60332 27396
rect 64696 27344 64748 27396
rect 42616 27276 42668 27328
rect 56600 27319 56652 27328
rect 56600 27285 56609 27319
rect 56609 27285 56643 27319
rect 56643 27285 56652 27319
rect 56600 27276 56652 27285
rect 70400 27276 70452 27328
rect 71412 27276 71464 27328
rect 77576 27344 77628 27396
rect 78220 27344 78272 27396
rect 84844 27276 84896 27328
rect 95240 27276 95292 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 65686 27174 65738 27226
rect 65750 27174 65802 27226
rect 65814 27174 65866 27226
rect 65878 27174 65930 27226
rect 96406 27174 96458 27226
rect 96470 27174 96522 27226
rect 96534 27174 96586 27226
rect 96598 27174 96650 27226
rect 16028 27072 16080 27124
rect 11704 27004 11756 27056
rect 12624 27004 12676 27056
rect 84844 27072 84896 27124
rect 28908 27004 28960 27056
rect 42616 27004 42668 27056
rect 46112 27004 46164 27056
rect 7472 26911 7524 26920
rect 7472 26877 7481 26911
rect 7481 26877 7515 26911
rect 7515 26877 7524 26911
rect 7472 26868 7524 26877
rect 17868 26936 17920 26988
rect 8116 26868 8168 26920
rect 20536 26911 20588 26920
rect 12624 26800 12676 26852
rect 20536 26877 20545 26911
rect 20545 26877 20579 26911
rect 20579 26877 20588 26911
rect 20536 26868 20588 26877
rect 21088 26911 21140 26920
rect 21088 26877 21097 26911
rect 21097 26877 21131 26911
rect 21131 26877 21140 26911
rect 21088 26868 21140 26877
rect 41420 26936 41472 26988
rect 46296 26936 46348 26988
rect 87052 26936 87104 26988
rect 45008 26868 45060 26920
rect 57060 26868 57112 26920
rect 70400 26868 70452 26920
rect 21364 26800 21416 26852
rect 23020 26800 23072 26852
rect 35348 26800 35400 26852
rect 41696 26732 41748 26784
rect 46296 26732 46348 26784
rect 61568 26732 61620 26784
rect 62028 26732 62080 26784
rect 69020 26732 69072 26784
rect 69756 26732 69808 26784
rect 87052 26732 87104 26784
rect 87420 26732 87472 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 50326 26630 50378 26682
rect 50390 26630 50442 26682
rect 50454 26630 50506 26682
rect 50518 26630 50570 26682
rect 81046 26630 81098 26682
rect 81110 26630 81162 26682
rect 81174 26630 81226 26682
rect 81238 26630 81290 26682
rect 21732 26528 21784 26580
rect 32956 26528 33008 26580
rect 40040 26528 40092 26580
rect 87420 26528 87472 26580
rect 17224 26392 17276 26444
rect 34704 26435 34756 26444
rect 34704 26401 34713 26435
rect 34713 26401 34747 26435
rect 34747 26401 34756 26435
rect 34704 26392 34756 26401
rect 17684 26256 17736 26308
rect 19432 26256 19484 26308
rect 21088 26324 21140 26376
rect 34520 26231 34572 26240
rect 34520 26197 34529 26231
rect 34529 26197 34563 26231
rect 34563 26197 34572 26231
rect 42800 26256 42852 26308
rect 43260 26256 43312 26308
rect 84384 26256 84436 26308
rect 95976 26256 96028 26308
rect 34520 26188 34572 26197
rect 72332 26188 72384 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 65686 26086 65738 26138
rect 65750 26086 65802 26138
rect 65814 26086 65866 26138
rect 65878 26086 65930 26138
rect 96406 26086 96458 26138
rect 96470 26086 96522 26138
rect 96534 26086 96586 26138
rect 96598 26086 96650 26138
rect 10600 25984 10652 26036
rect 21088 25984 21140 26036
rect 22652 25984 22704 26036
rect 43812 25984 43864 26036
rect 44088 25984 44140 26036
rect 44456 25984 44508 26036
rect 69480 25984 69532 26036
rect 13268 25916 13320 25968
rect 44272 25916 44324 25968
rect 7748 25848 7800 25900
rect 57336 25916 57388 25968
rect 72792 25848 72844 25900
rect 80152 25848 80204 25900
rect 42248 25780 42300 25832
rect 5908 25712 5960 25764
rect 45100 25712 45152 25764
rect 49608 25780 49660 25832
rect 75000 25823 75052 25832
rect 75000 25789 75009 25823
rect 75009 25789 75043 25823
rect 75043 25789 75052 25823
rect 75000 25780 75052 25789
rect 49700 25712 49752 25764
rect 56784 25712 56836 25764
rect 73896 25712 73948 25764
rect 75920 25712 75972 25764
rect 10508 25644 10560 25696
rect 66076 25644 66128 25696
rect 66260 25644 66312 25696
rect 67088 25644 67140 25696
rect 92480 25644 92532 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 50326 25542 50378 25594
rect 50390 25542 50442 25594
rect 50454 25542 50506 25594
rect 50518 25542 50570 25594
rect 81046 25542 81098 25594
rect 81110 25542 81162 25594
rect 81174 25542 81226 25594
rect 81238 25542 81290 25594
rect 27804 25440 27856 25492
rect 39396 25440 39448 25492
rect 44088 25440 44140 25492
rect 66260 25440 66312 25492
rect 71320 25440 71372 25492
rect 35532 25372 35584 25424
rect 80152 25415 80204 25424
rect 80152 25381 80161 25415
rect 80161 25381 80195 25415
rect 80195 25381 80204 25415
rect 80152 25372 80204 25381
rect 65156 25304 65208 25356
rect 44364 25236 44416 25288
rect 78220 25279 78272 25288
rect 78220 25245 78229 25279
rect 78229 25245 78263 25279
rect 78263 25245 78272 25279
rect 78220 25236 78272 25245
rect 78496 25279 78548 25288
rect 78496 25245 78505 25279
rect 78505 25245 78539 25279
rect 78539 25245 78548 25279
rect 78496 25236 78548 25245
rect 80244 25236 80296 25288
rect 72332 25168 72384 25220
rect 72700 25168 72752 25220
rect 46848 25100 46900 25152
rect 73804 25100 73856 25152
rect 75920 25100 75972 25152
rect 76656 25100 76708 25152
rect 79600 25143 79652 25152
rect 79600 25109 79609 25143
rect 79609 25109 79643 25143
rect 79643 25109 79652 25143
rect 79600 25100 79652 25109
rect 80980 25143 81032 25152
rect 80980 25109 80989 25143
rect 80989 25109 81023 25143
rect 81023 25109 81032 25143
rect 80980 25100 81032 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 65686 24998 65738 25050
rect 65750 24998 65802 25050
rect 65814 24998 65866 25050
rect 65878 24998 65930 25050
rect 96406 24998 96458 25050
rect 96470 24998 96522 25050
rect 96534 24998 96586 25050
rect 96598 24998 96650 25050
rect 9956 24871 10008 24880
rect 9956 24837 9965 24871
rect 9965 24837 9999 24871
rect 9999 24837 10008 24871
rect 9956 24828 10008 24837
rect 10048 24803 10100 24812
rect 10048 24769 10057 24803
rect 10057 24769 10091 24803
rect 10091 24769 10100 24803
rect 10048 24760 10100 24769
rect 71412 24896 71464 24948
rect 72792 24896 72844 24948
rect 77024 24896 77076 24948
rect 80244 24896 80296 24948
rect 16028 24828 16080 24880
rect 18788 24828 18840 24880
rect 43352 24828 43404 24880
rect 80980 24828 81032 24880
rect 10508 24760 10560 24812
rect 9128 24599 9180 24608
rect 9128 24565 9137 24599
rect 9137 24565 9171 24599
rect 9171 24565 9180 24599
rect 12716 24692 12768 24744
rect 14924 24692 14976 24744
rect 19156 24692 19208 24744
rect 19432 24692 19484 24744
rect 30564 24760 30616 24812
rect 36084 24760 36136 24812
rect 54208 24760 54260 24812
rect 20076 24692 20128 24744
rect 34520 24692 34572 24744
rect 35808 24692 35860 24744
rect 59360 24692 59412 24744
rect 80796 24692 80848 24744
rect 85580 24692 85632 24744
rect 86224 24735 86276 24744
rect 86224 24701 86233 24735
rect 86233 24701 86267 24735
rect 86267 24701 86276 24735
rect 86224 24692 86276 24701
rect 86408 24735 86460 24744
rect 86408 24701 86417 24735
rect 86417 24701 86451 24735
rect 86451 24701 86460 24735
rect 86408 24692 86460 24701
rect 10600 24599 10652 24608
rect 9128 24556 9180 24565
rect 10600 24565 10609 24599
rect 10609 24565 10643 24599
rect 10643 24565 10652 24599
rect 10600 24556 10652 24565
rect 21272 24599 21324 24608
rect 21272 24565 21281 24599
rect 21281 24565 21315 24599
rect 21315 24565 21324 24599
rect 21272 24556 21324 24565
rect 35440 24599 35492 24608
rect 35440 24565 35449 24599
rect 35449 24565 35483 24599
rect 35483 24565 35492 24599
rect 35440 24556 35492 24565
rect 35716 24599 35768 24608
rect 35716 24565 35725 24599
rect 35725 24565 35759 24599
rect 35759 24565 35768 24599
rect 35716 24556 35768 24565
rect 36084 24556 36136 24608
rect 85212 24556 85264 24608
rect 85396 24556 85448 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 50326 24454 50378 24506
rect 50390 24454 50442 24506
rect 50454 24454 50506 24506
rect 50518 24454 50570 24506
rect 81046 24454 81098 24506
rect 81110 24454 81162 24506
rect 81174 24454 81226 24506
rect 81238 24454 81290 24506
rect 9128 24352 9180 24404
rect 41420 24352 41472 24404
rect 21272 24284 21324 24336
rect 36636 24284 36688 24336
rect 9956 24216 10008 24268
rect 35348 24216 35400 24268
rect 36636 24148 36688 24200
rect 52276 24148 52328 24200
rect 11060 24080 11112 24132
rect 11796 24080 11848 24132
rect 31392 24080 31444 24132
rect 40960 24080 41012 24132
rect 64972 24080 65024 24132
rect 20076 24012 20128 24064
rect 80060 24012 80112 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 65686 23910 65738 23962
rect 65750 23910 65802 23962
rect 65814 23910 65866 23962
rect 65878 23910 65930 23962
rect 96406 23910 96458 23962
rect 96470 23910 96522 23962
rect 96534 23910 96586 23962
rect 96598 23910 96650 23962
rect 9772 23808 9824 23860
rect 85212 23808 85264 23860
rect 10600 23740 10652 23792
rect 41696 23740 41748 23792
rect 42248 23740 42300 23792
rect 49424 23740 49476 23792
rect 5724 23672 5776 23724
rect 12716 23672 12768 23724
rect 40316 23672 40368 23724
rect 66904 23672 66956 23724
rect 31668 23604 31720 23656
rect 40040 23647 40092 23656
rect 40040 23613 40049 23647
rect 40049 23613 40083 23647
rect 40083 23613 40092 23647
rect 40040 23604 40092 23613
rect 11060 23536 11112 23588
rect 49240 23536 49292 23588
rect 48964 23468 49016 23520
rect 49516 23468 49568 23520
rect 72884 23468 72936 23520
rect 77852 23604 77904 23656
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 50326 23366 50378 23418
rect 50390 23366 50442 23418
rect 50454 23366 50506 23418
rect 50518 23366 50570 23418
rect 81046 23366 81098 23418
rect 81110 23366 81162 23418
rect 81174 23366 81226 23418
rect 81238 23366 81290 23418
rect 16120 23264 16172 23316
rect 78772 23264 78824 23316
rect 44548 23196 44600 23248
rect 16396 23128 16448 23180
rect 29552 23060 29604 23112
rect 46020 23060 46072 23112
rect 59728 23128 59780 23180
rect 60372 23171 60424 23180
rect 60372 23137 60381 23171
rect 60381 23137 60415 23171
rect 60415 23137 60424 23171
rect 60372 23128 60424 23137
rect 60740 23171 60792 23180
rect 60740 23137 60749 23171
rect 60749 23137 60783 23171
rect 60783 23137 60792 23171
rect 60740 23128 60792 23137
rect 61568 23128 61620 23180
rect 78220 23128 78272 23180
rect 90180 23128 90232 23180
rect 60096 23103 60148 23112
rect 60096 23069 60105 23103
rect 60105 23069 60139 23103
rect 60139 23069 60148 23103
rect 60096 23060 60148 23069
rect 3424 22992 3476 23044
rect 35440 22992 35492 23044
rect 43720 22992 43772 23044
rect 77944 23103 77996 23112
rect 77944 23069 77953 23103
rect 77953 23069 77987 23103
rect 77987 23069 77996 23103
rect 77944 23060 77996 23069
rect 72056 22992 72108 23044
rect 59728 22967 59780 22976
rect 59728 22933 59737 22967
rect 59737 22933 59771 22967
rect 59771 22933 59780 22967
rect 59728 22924 59780 22933
rect 79416 22924 79468 22976
rect 85120 22924 85172 22976
rect 95884 22924 95936 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 65686 22822 65738 22874
rect 65750 22822 65802 22874
rect 65814 22822 65866 22874
rect 65878 22822 65930 22874
rect 96406 22822 96458 22874
rect 96470 22822 96522 22874
rect 96534 22822 96586 22874
rect 96598 22822 96650 22874
rect 6368 22720 6420 22772
rect 66996 22720 67048 22772
rect 49516 22652 49568 22704
rect 79508 22652 79560 22704
rect 15108 22584 15160 22636
rect 57520 22584 57572 22636
rect 19156 22559 19208 22568
rect 19156 22525 19165 22559
rect 19165 22525 19199 22559
rect 19199 22525 19208 22559
rect 19156 22516 19208 22525
rect 19432 22559 19484 22568
rect 19432 22525 19441 22559
rect 19441 22525 19475 22559
rect 19475 22525 19484 22559
rect 19432 22516 19484 22525
rect 22100 22448 22152 22500
rect 23112 22448 23164 22500
rect 48872 22516 48924 22568
rect 47584 22448 47636 22500
rect 48320 22448 48372 22500
rect 79416 22448 79468 22500
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 50326 22278 50378 22330
rect 50390 22278 50442 22330
rect 50454 22278 50506 22330
rect 50518 22278 50570 22330
rect 81046 22278 81098 22330
rect 81110 22278 81162 22330
rect 81174 22278 81226 22330
rect 81238 22278 81290 22330
rect 19432 22176 19484 22228
rect 61844 22176 61896 22228
rect 36176 22151 36228 22160
rect 36176 22117 36185 22151
rect 36185 22117 36219 22151
rect 36219 22117 36228 22151
rect 36176 22108 36228 22117
rect 65524 22108 65576 22160
rect 72240 22108 72292 22160
rect 76564 22108 76616 22160
rect 36912 22083 36964 22092
rect 36912 22049 36921 22083
rect 36921 22049 36955 22083
rect 36955 22049 36964 22083
rect 36912 22040 36964 22049
rect 36084 21972 36136 22024
rect 43076 21972 43128 22024
rect 47400 21972 47452 22024
rect 47952 22040 48004 22092
rect 71136 22040 71188 22092
rect 88156 21972 88208 22024
rect 33784 21904 33836 21956
rect 34336 21904 34388 21956
rect 26792 21836 26844 21888
rect 35624 21836 35676 21888
rect 50068 21904 50120 21956
rect 64420 21904 64472 21956
rect 63040 21836 63092 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 65686 21734 65738 21786
rect 65750 21734 65802 21786
rect 65814 21734 65866 21786
rect 65878 21734 65930 21786
rect 96406 21734 96458 21786
rect 96470 21734 96522 21786
rect 96534 21734 96586 21786
rect 96598 21734 96650 21786
rect 11980 21632 12032 21684
rect 28816 21632 28868 21684
rect 35348 21632 35400 21684
rect 35716 21632 35768 21684
rect 43720 21632 43772 21684
rect 69572 21632 69624 21684
rect 22376 21564 22428 21616
rect 22836 21564 22888 21616
rect 48872 21564 48924 21616
rect 76564 21564 76616 21616
rect 76932 21564 76984 21616
rect 15384 21496 15436 21548
rect 28264 21496 28316 21548
rect 28356 21496 28408 21548
rect 64512 21496 64564 21548
rect 76748 21496 76800 21548
rect 12716 21428 12768 21480
rect 26792 21428 26844 21480
rect 26976 21428 27028 21480
rect 33876 21428 33928 21480
rect 80612 21471 80664 21480
rect 80612 21437 80621 21471
rect 80621 21437 80655 21471
rect 80655 21437 80664 21471
rect 80612 21428 80664 21437
rect 80796 21471 80848 21480
rect 80796 21437 80805 21471
rect 80805 21437 80839 21471
rect 80839 21437 80848 21471
rect 80796 21428 80848 21437
rect 1676 21360 1728 21412
rect 28632 21360 28684 21412
rect 33968 21360 34020 21412
rect 35624 21292 35676 21344
rect 56140 21360 56192 21412
rect 58992 21360 59044 21412
rect 57152 21292 57204 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 50326 21190 50378 21242
rect 50390 21190 50442 21242
rect 50454 21190 50506 21242
rect 50518 21190 50570 21242
rect 81046 21190 81098 21242
rect 81110 21190 81162 21242
rect 81174 21190 81226 21242
rect 81238 21190 81290 21242
rect 77668 21088 77720 21140
rect 77668 20995 77720 21004
rect 77668 20961 77677 20995
rect 77677 20961 77711 20995
rect 77711 20961 77720 20995
rect 97172 21088 97224 21140
rect 77668 20952 77720 20961
rect 90180 20952 90232 21004
rect 20720 20748 20772 20800
rect 21916 20748 21968 20800
rect 50068 20748 50120 20800
rect 71320 20748 71372 20800
rect 95240 20748 95292 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 65686 20646 65738 20698
rect 65750 20646 65802 20698
rect 65814 20646 65866 20698
rect 65878 20646 65930 20698
rect 96406 20646 96458 20698
rect 96470 20646 96522 20698
rect 96534 20646 96586 20698
rect 96598 20646 96650 20698
rect 21916 20544 21968 20596
rect 24216 20544 24268 20596
rect 64236 20544 64288 20596
rect 66260 20544 66312 20596
rect 10784 20476 10836 20528
rect 4804 20340 4856 20392
rect 5264 20340 5316 20392
rect 15844 20340 15896 20392
rect 19432 20340 19484 20392
rect 23940 20383 23992 20392
rect 23940 20349 23949 20383
rect 23949 20349 23983 20383
rect 23983 20349 23992 20383
rect 23940 20340 23992 20349
rect 24308 20451 24360 20460
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24308 20408 24360 20417
rect 24216 20383 24268 20392
rect 24216 20349 24225 20383
rect 24225 20349 24259 20383
rect 24259 20349 24268 20383
rect 30196 20408 30248 20460
rect 88432 20408 88484 20460
rect 24216 20340 24268 20349
rect 24492 20383 24544 20392
rect 24492 20349 24501 20383
rect 24501 20349 24535 20383
rect 24535 20349 24544 20383
rect 24492 20340 24544 20349
rect 24860 20340 24912 20392
rect 55036 20340 55088 20392
rect 78128 20383 78180 20392
rect 78128 20349 78137 20383
rect 78137 20349 78171 20383
rect 78171 20349 78180 20383
rect 78128 20340 78180 20349
rect 45284 20272 45336 20324
rect 12808 20204 12860 20256
rect 24492 20204 24544 20256
rect 28172 20204 28224 20256
rect 43628 20204 43680 20256
rect 62856 20204 62908 20256
rect 74172 20204 74224 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 50326 20102 50378 20154
rect 50390 20102 50442 20154
rect 50454 20102 50506 20154
rect 50518 20102 50570 20154
rect 81046 20102 81098 20154
rect 81110 20102 81162 20154
rect 81174 20102 81226 20154
rect 81238 20102 81290 20154
rect 16120 20000 16172 20052
rect 24308 20000 24360 20052
rect 65156 20043 65208 20052
rect 65156 20009 65165 20043
rect 65165 20009 65199 20043
rect 65199 20009 65208 20043
rect 65156 20000 65208 20009
rect 71688 20000 71740 20052
rect 95240 20000 95292 20052
rect 19064 19932 19116 19984
rect 24216 19932 24268 19984
rect 24860 19932 24912 19984
rect 25872 19932 25924 19984
rect 62212 19932 62264 19984
rect 64696 19932 64748 19984
rect 83648 19932 83700 19984
rect 88800 19975 88852 19984
rect 88800 19941 88809 19975
rect 88809 19941 88843 19975
rect 88843 19941 88852 19975
rect 88800 19932 88852 19941
rect 28172 19864 28224 19916
rect 61752 19864 61804 19916
rect 64972 19907 65024 19916
rect 64972 19873 64981 19907
rect 64981 19873 65015 19907
rect 65015 19873 65024 19907
rect 64972 19864 65024 19873
rect 68376 19864 68428 19916
rect 72884 19907 72936 19916
rect 72884 19873 72893 19907
rect 72893 19873 72927 19907
rect 72927 19873 72936 19907
rect 72884 19864 72936 19873
rect 73252 19907 73304 19916
rect 45284 19796 45336 19848
rect 50896 19796 50948 19848
rect 73252 19873 73261 19907
rect 73261 19873 73295 19907
rect 73295 19873 73304 19907
rect 73252 19864 73304 19873
rect 82636 19864 82688 19916
rect 85856 19864 85908 19916
rect 90548 19864 90600 19916
rect 90180 19796 90232 19848
rect 90456 19796 90508 19848
rect 56140 19728 56192 19780
rect 43076 19660 43128 19712
rect 46112 19660 46164 19712
rect 89628 19660 89680 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 65686 19558 65738 19610
rect 65750 19558 65802 19610
rect 65814 19558 65866 19610
rect 65878 19558 65930 19610
rect 96406 19558 96458 19610
rect 96470 19558 96522 19610
rect 96534 19558 96586 19610
rect 96598 19558 96650 19610
rect 8944 19320 8996 19372
rect 43076 19456 43128 19508
rect 44548 19388 44600 19440
rect 44456 19320 44508 19372
rect 12256 19252 12308 19304
rect 20996 19252 21048 19304
rect 24124 19252 24176 19304
rect 43168 19252 43220 19304
rect 44640 19295 44692 19304
rect 44640 19261 44649 19295
rect 44649 19261 44683 19295
rect 44683 19261 44692 19295
rect 45100 19320 45152 19372
rect 45376 19320 45428 19372
rect 46112 19320 46164 19372
rect 71688 19320 71740 19372
rect 44640 19252 44692 19261
rect 45008 19295 45060 19304
rect 45008 19261 45017 19295
rect 45017 19261 45051 19295
rect 45051 19261 45060 19295
rect 45008 19252 45060 19261
rect 45192 19295 45244 19304
rect 45192 19261 45201 19295
rect 45201 19261 45235 19295
rect 45235 19261 45244 19295
rect 45192 19252 45244 19261
rect 50620 19295 50672 19304
rect 50620 19261 50629 19295
rect 50629 19261 50663 19295
rect 50663 19261 50672 19295
rect 50620 19252 50672 19261
rect 67640 19252 67692 19304
rect 28540 19116 28592 19168
rect 62120 19184 62172 19236
rect 62764 19184 62816 19236
rect 86868 19184 86920 19236
rect 50160 19116 50212 19168
rect 50620 19116 50672 19168
rect 54116 19116 54168 19168
rect 73436 19116 73488 19168
rect 95240 19184 95292 19236
rect 90640 19116 90692 19168
rect 97264 19116 97316 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 50326 19014 50378 19066
rect 50390 19014 50442 19066
rect 50454 19014 50506 19066
rect 50518 19014 50570 19066
rect 81046 19014 81098 19066
rect 81110 19014 81162 19066
rect 81174 19014 81226 19066
rect 81238 19014 81290 19066
rect 3976 18912 4028 18964
rect 29000 18844 29052 18896
rect 29736 18844 29788 18896
rect 45192 18844 45244 18896
rect 53380 18844 53432 18896
rect 62948 18844 63000 18896
rect 63408 18844 63460 18896
rect 65432 18912 65484 18964
rect 96160 18912 96212 18964
rect 64880 18844 64932 18896
rect 70584 18844 70636 18896
rect 73436 18844 73488 18896
rect 79416 18844 79468 18896
rect 39488 18776 39540 18828
rect 57428 18776 57480 18828
rect 65340 18776 65392 18828
rect 96988 18819 97040 18828
rect 96988 18785 96997 18819
rect 96997 18785 97031 18819
rect 97031 18785 97040 18819
rect 96988 18776 97040 18785
rect 42800 18708 42852 18760
rect 47400 18751 47452 18760
rect 47400 18717 47409 18751
rect 47409 18717 47443 18751
rect 47443 18717 47452 18751
rect 47400 18708 47452 18717
rect 55036 18708 55088 18760
rect 61936 18751 61988 18760
rect 61936 18717 61945 18751
rect 61945 18717 61979 18751
rect 61979 18717 61988 18751
rect 61936 18708 61988 18717
rect 62672 18708 62724 18760
rect 97264 18819 97316 18828
rect 97264 18785 97273 18819
rect 97273 18785 97307 18819
rect 97307 18785 97316 18819
rect 97264 18776 97316 18785
rect 12256 18640 12308 18692
rect 20720 18640 20772 18692
rect 34520 18640 34572 18692
rect 35808 18640 35860 18692
rect 38108 18640 38160 18692
rect 46848 18572 46900 18624
rect 50620 18640 50672 18692
rect 59452 18640 59504 18692
rect 49976 18572 50028 18624
rect 55956 18572 56008 18624
rect 77944 18640 77996 18692
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 65686 18470 65738 18522
rect 65750 18470 65802 18522
rect 65814 18470 65866 18522
rect 65878 18470 65930 18522
rect 96406 18470 96458 18522
rect 96470 18470 96522 18522
rect 96534 18470 96586 18522
rect 96598 18470 96650 18522
rect 62120 18368 62172 18420
rect 73344 18411 73396 18420
rect 58256 18300 58308 18352
rect 67640 18300 67692 18352
rect 19432 18232 19484 18284
rect 19892 18232 19944 18284
rect 28356 18232 28408 18284
rect 34520 18232 34572 18284
rect 19340 18207 19392 18216
rect 19340 18173 19349 18207
rect 19349 18173 19383 18207
rect 19383 18173 19392 18207
rect 19340 18164 19392 18173
rect 30196 18207 30248 18216
rect 30196 18173 30205 18207
rect 30205 18173 30239 18207
rect 30239 18173 30248 18207
rect 30196 18164 30248 18173
rect 31668 18164 31720 18216
rect 55036 18207 55088 18216
rect 18604 18096 18656 18148
rect 55036 18173 55045 18207
rect 55045 18173 55079 18207
rect 55079 18173 55088 18207
rect 55036 18164 55088 18173
rect 55312 18207 55364 18216
rect 55312 18173 55321 18207
rect 55321 18173 55355 18207
rect 55355 18173 55364 18207
rect 55312 18164 55364 18173
rect 55956 18232 56008 18284
rect 67732 18232 67784 18284
rect 71136 18300 71188 18352
rect 71320 18343 71372 18352
rect 71320 18309 71329 18343
rect 71329 18309 71363 18343
rect 71363 18309 71372 18343
rect 71320 18300 71372 18309
rect 70584 18207 70636 18216
rect 70584 18173 70593 18207
rect 70593 18173 70627 18207
rect 70627 18173 70636 18207
rect 70584 18164 70636 18173
rect 71688 18164 71740 18216
rect 73344 18377 73353 18411
rect 73353 18377 73387 18411
rect 73387 18377 73396 18411
rect 73344 18368 73396 18377
rect 59728 18096 59780 18148
rect 70492 18096 70544 18148
rect 71320 18096 71372 18148
rect 96712 18096 96764 18148
rect 96988 18096 97040 18148
rect 38108 18028 38160 18080
rect 42800 18028 42852 18080
rect 51264 18028 51316 18080
rect 53288 18028 53340 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 50326 17926 50378 17978
rect 50390 17926 50442 17978
rect 50454 17926 50506 17978
rect 50518 17926 50570 17978
rect 81046 17926 81098 17978
rect 81110 17926 81162 17978
rect 81174 17926 81226 17978
rect 81238 17926 81290 17978
rect 60280 17824 60332 17876
rect 61108 17824 61160 17876
rect 66996 17824 67048 17876
rect 69848 17824 69900 17876
rect 34060 17620 34112 17672
rect 39856 17620 39908 17672
rect 44456 17620 44508 17672
rect 48320 17620 48372 17672
rect 73712 17620 73764 17672
rect 24768 17552 24820 17604
rect 77668 17552 77720 17604
rect 17132 17527 17184 17536
rect 17132 17493 17141 17527
rect 17141 17493 17175 17527
rect 17175 17493 17184 17527
rect 17132 17484 17184 17493
rect 25964 17484 26016 17536
rect 31116 17484 31168 17536
rect 34244 17484 34296 17536
rect 43812 17484 43864 17536
rect 62396 17484 62448 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 65686 17382 65738 17434
rect 65750 17382 65802 17434
rect 65814 17382 65866 17434
rect 65878 17382 65930 17434
rect 96406 17382 96458 17434
rect 96470 17382 96522 17434
rect 96534 17382 96586 17434
rect 96598 17382 96650 17434
rect 26332 17280 26384 17332
rect 72608 17280 72660 17332
rect 81532 17280 81584 17332
rect 4988 17212 5040 17264
rect 71228 17212 71280 17264
rect 72424 17212 72476 17264
rect 79876 17212 79928 17264
rect 80152 17212 80204 17264
rect 17132 17144 17184 17196
rect 33692 17144 33744 17196
rect 44640 17144 44692 17196
rect 66996 17144 67048 17196
rect 72516 17144 72568 17196
rect 81532 17144 81584 17196
rect 46480 17076 46532 17128
rect 49056 17008 49108 17060
rect 55312 17008 55364 17060
rect 86868 17119 86920 17128
rect 86868 17085 86877 17119
rect 86877 17085 86911 17119
rect 86911 17085 86920 17119
rect 86868 17076 86920 17085
rect 87420 17119 87472 17128
rect 87420 17085 87429 17119
rect 87429 17085 87463 17119
rect 87463 17085 87472 17119
rect 87420 17076 87472 17085
rect 97172 17119 97224 17128
rect 97172 17085 97181 17119
rect 97181 17085 97215 17119
rect 97215 17085 97224 17119
rect 97172 17076 97224 17085
rect 21180 16940 21232 16992
rect 21364 16940 21416 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 50326 16838 50378 16890
rect 50390 16838 50442 16890
rect 50454 16838 50506 16890
rect 50518 16838 50570 16890
rect 81046 16838 81098 16890
rect 81110 16838 81162 16890
rect 81174 16838 81226 16890
rect 81238 16838 81290 16890
rect 44732 16779 44784 16788
rect 6276 16668 6328 16720
rect 8576 16668 8628 16720
rect 44732 16745 44741 16779
rect 44741 16745 44775 16779
rect 44775 16745 44784 16779
rect 44732 16736 44784 16745
rect 47676 16779 47728 16788
rect 47676 16745 47685 16779
rect 47685 16745 47719 16779
rect 47719 16745 47728 16779
rect 47676 16736 47728 16745
rect 24308 16668 24360 16720
rect 24768 16668 24820 16720
rect 8944 16600 8996 16652
rect 20260 16600 20312 16652
rect 44456 16668 44508 16720
rect 44640 16711 44692 16720
rect 44640 16677 44649 16711
rect 44649 16677 44683 16711
rect 44683 16677 44692 16711
rect 44640 16668 44692 16677
rect 48044 16736 48096 16788
rect 48320 16736 48372 16788
rect 48504 16600 48556 16652
rect 58624 16736 58676 16788
rect 68376 16736 68428 16788
rect 97172 16736 97224 16788
rect 49700 16600 49752 16652
rect 50160 16600 50212 16652
rect 14556 16532 14608 16584
rect 79416 16532 79468 16584
rect 46204 16396 46256 16448
rect 67548 16396 67600 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 65686 16294 65738 16346
rect 65750 16294 65802 16346
rect 65814 16294 65866 16346
rect 65878 16294 65930 16346
rect 96406 16294 96458 16346
rect 96470 16294 96522 16346
rect 96534 16294 96586 16346
rect 96598 16294 96650 16346
rect 25964 16192 26016 16244
rect 42432 16192 42484 16244
rect 59268 16192 59320 16244
rect 95976 16192 96028 16244
rect 37832 16124 37884 16176
rect 85948 16124 86000 16176
rect 9864 16056 9916 16108
rect 29000 16056 29052 16108
rect 40040 16056 40092 16108
rect 89076 16056 89128 16108
rect 19248 15988 19300 16040
rect 71412 15988 71464 16040
rect 2504 15920 2556 15972
rect 13636 15920 13688 15972
rect 17776 15920 17828 15972
rect 80336 15920 80388 15972
rect 2412 15852 2464 15904
rect 69756 15852 69808 15904
rect 79416 15852 79468 15904
rect 93860 15852 93912 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 50326 15750 50378 15802
rect 50390 15750 50442 15802
rect 50454 15750 50506 15802
rect 50518 15750 50570 15802
rect 81046 15750 81098 15802
rect 81110 15750 81162 15802
rect 81174 15750 81226 15802
rect 81238 15750 81290 15802
rect 58072 15691 58124 15700
rect 58072 15657 58081 15691
rect 58081 15657 58115 15691
rect 58115 15657 58124 15691
rect 58072 15648 58124 15657
rect 57980 15623 58032 15632
rect 57980 15589 57989 15623
rect 57989 15589 58023 15623
rect 58023 15589 58032 15623
rect 57980 15580 58032 15589
rect 13636 15376 13688 15428
rect 31668 15376 31720 15428
rect 92296 15308 92348 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 65686 15206 65738 15258
rect 65750 15206 65802 15258
rect 65814 15206 65866 15258
rect 65878 15206 65930 15258
rect 96406 15206 96458 15258
rect 96470 15206 96522 15258
rect 96534 15206 96586 15258
rect 96598 15206 96650 15258
rect 14004 15104 14056 15156
rect 14556 15104 14608 15156
rect 15568 15104 15620 15156
rect 18696 15036 18748 15088
rect 55772 15104 55824 15156
rect 84384 15104 84436 15156
rect 59452 15036 59504 15088
rect 61844 15036 61896 15088
rect 97816 15036 97868 15088
rect 13636 14943 13688 14952
rect 13636 14909 13645 14943
rect 13645 14909 13679 14943
rect 13679 14909 13688 14943
rect 13636 14900 13688 14909
rect 15936 14968 15988 15020
rect 63408 14968 63460 15020
rect 14004 14943 14056 14952
rect 14004 14909 14013 14943
rect 14013 14909 14047 14943
rect 14047 14909 14056 14943
rect 14004 14900 14056 14909
rect 35256 14900 35308 14952
rect 44824 14900 44876 14952
rect 13820 14832 13872 14884
rect 17224 14832 17276 14884
rect 33968 14832 34020 14884
rect 55220 14832 55272 14884
rect 97908 14900 97960 14952
rect 66812 14764 66864 14816
rect 96068 14832 96120 14884
rect 87788 14764 87840 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 50326 14662 50378 14714
rect 50390 14662 50442 14714
rect 50454 14662 50506 14714
rect 50518 14662 50570 14714
rect 81046 14662 81098 14714
rect 81110 14662 81162 14714
rect 81174 14662 81226 14714
rect 81238 14662 81290 14714
rect 18512 14560 18564 14612
rect 81624 14560 81676 14612
rect 23020 14492 23072 14544
rect 92112 14492 92164 14544
rect 13544 14424 13596 14476
rect 42984 14424 43036 14476
rect 44364 14467 44416 14476
rect 44364 14433 44373 14467
rect 44373 14433 44407 14467
rect 44407 14433 44416 14467
rect 44364 14424 44416 14433
rect 44732 14467 44784 14476
rect 44732 14433 44741 14467
rect 44741 14433 44775 14467
rect 44775 14433 44784 14467
rect 44732 14424 44784 14433
rect 44824 14424 44876 14476
rect 45008 14424 45060 14476
rect 75000 14424 75052 14476
rect 82912 14467 82964 14476
rect 82912 14433 82921 14467
rect 82921 14433 82955 14467
rect 82955 14433 82964 14467
rect 82912 14424 82964 14433
rect 22100 14288 22152 14340
rect 44548 14288 44600 14340
rect 77024 14356 77076 14408
rect 45376 14288 45428 14340
rect 57244 14288 57296 14340
rect 61660 14288 61712 14340
rect 67180 14288 67232 14340
rect 37740 14263 37792 14272
rect 37740 14229 37749 14263
rect 37749 14229 37783 14263
rect 37783 14229 37792 14263
rect 37740 14220 37792 14229
rect 46664 14220 46716 14272
rect 49700 14220 49752 14272
rect 54484 14220 54536 14272
rect 55220 14220 55272 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 65686 14118 65738 14170
rect 65750 14118 65802 14170
rect 65814 14118 65866 14170
rect 65878 14118 65930 14170
rect 96406 14118 96458 14170
rect 96470 14118 96522 14170
rect 96534 14118 96586 14170
rect 96598 14118 96650 14170
rect 37740 14016 37792 14068
rect 62488 14016 62540 14068
rect 49608 13948 49660 14000
rect 46664 13880 46716 13932
rect 49700 13880 49752 13932
rect 12164 13812 12216 13864
rect 16304 13812 16356 13864
rect 23204 13812 23256 13864
rect 39764 13855 39816 13864
rect 39764 13821 39773 13855
rect 39773 13821 39807 13855
rect 39807 13821 39816 13855
rect 39764 13812 39816 13821
rect 29368 13744 29420 13796
rect 29736 13744 29788 13796
rect 92204 13744 92256 13796
rect 94044 13744 94096 13796
rect 44732 13676 44784 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 50326 13574 50378 13626
rect 50390 13574 50442 13626
rect 50454 13574 50506 13626
rect 50518 13574 50570 13626
rect 81046 13574 81098 13626
rect 81110 13574 81162 13626
rect 81174 13574 81226 13626
rect 81238 13574 81290 13626
rect 10968 13472 11020 13524
rect 36452 13472 36504 13524
rect 37188 13472 37240 13524
rect 11428 13336 11480 13388
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 12532 13404 12584 13456
rect 19984 13404 20036 13456
rect 9312 13268 9364 13320
rect 31024 13336 31076 13388
rect 67364 13379 67416 13388
rect 67364 13345 67373 13379
rect 67373 13345 67407 13379
rect 67407 13345 67416 13379
rect 67364 13336 67416 13345
rect 12532 13268 12584 13320
rect 43260 13268 43312 13320
rect 61568 13268 61620 13320
rect 69756 13268 69808 13320
rect 39580 13200 39632 13252
rect 41420 13200 41472 13252
rect 61476 13200 61528 13252
rect 66628 13200 66680 13252
rect 88248 13200 88300 13252
rect 16948 13175 17000 13184
rect 16948 13141 16957 13175
rect 16957 13141 16991 13175
rect 16991 13141 17000 13175
rect 16948 13132 17000 13141
rect 28908 13132 28960 13184
rect 63776 13132 63828 13184
rect 66352 13132 66404 13184
rect 92204 13132 92256 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 65686 13030 65738 13082
rect 65750 13030 65802 13082
rect 65814 13030 65866 13082
rect 65878 13030 65930 13082
rect 96406 13030 96458 13082
rect 96470 13030 96522 13082
rect 96534 13030 96586 13082
rect 96598 13030 96650 13082
rect 37188 12928 37240 12980
rect 55956 12928 56008 12980
rect 60096 12928 60148 12980
rect 6092 12860 6144 12912
rect 6828 12860 6880 12912
rect 41052 12903 41104 12912
rect 41052 12869 41061 12903
rect 41061 12869 41095 12903
rect 41095 12869 41104 12903
rect 41052 12860 41104 12869
rect 32496 12792 32548 12844
rect 41144 12835 41196 12844
rect 41144 12801 41153 12835
rect 41153 12801 41187 12835
rect 41187 12801 41196 12835
rect 41144 12792 41196 12801
rect 41604 12860 41656 12912
rect 19064 12767 19116 12776
rect 19064 12733 19073 12767
rect 19073 12733 19107 12767
rect 19107 12733 19116 12767
rect 19064 12724 19116 12733
rect 23112 12724 23164 12776
rect 41604 12724 41656 12776
rect 56140 12860 56192 12912
rect 69756 12928 69808 12980
rect 55956 12792 56008 12844
rect 40776 12699 40828 12708
rect 40776 12665 40785 12699
rect 40785 12665 40819 12699
rect 40819 12665 40828 12699
rect 40776 12656 40828 12665
rect 56140 12724 56192 12776
rect 66352 12724 66404 12776
rect 66628 12767 66680 12776
rect 66628 12733 66637 12767
rect 66637 12733 66671 12767
rect 66671 12733 66680 12767
rect 66628 12724 66680 12733
rect 66812 12724 66864 12776
rect 66996 12767 67048 12776
rect 66996 12733 67005 12767
rect 67005 12733 67039 12767
rect 67039 12733 67048 12767
rect 66996 12724 67048 12733
rect 67088 12724 67140 12776
rect 67548 12767 67600 12776
rect 67548 12733 67557 12767
rect 67557 12733 67591 12767
rect 67591 12733 67600 12767
rect 67548 12724 67600 12733
rect 96712 12767 96764 12776
rect 29736 12588 29788 12640
rect 41052 12588 41104 12640
rect 82544 12656 82596 12708
rect 96712 12733 96721 12767
rect 96721 12733 96755 12767
rect 96755 12733 96764 12767
rect 96712 12724 96764 12733
rect 97816 12903 97868 12912
rect 97816 12869 97825 12903
rect 97825 12869 97859 12903
rect 97859 12869 97868 12903
rect 97816 12860 97868 12869
rect 84476 12588 84528 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 50326 12486 50378 12538
rect 50390 12486 50442 12538
rect 50454 12486 50506 12538
rect 50518 12486 50570 12538
rect 81046 12486 81098 12538
rect 81110 12486 81162 12538
rect 81174 12486 81226 12538
rect 81238 12486 81290 12538
rect 27712 12384 27764 12436
rect 27988 12384 28040 12436
rect 38108 12291 38160 12300
rect 38108 12257 38117 12291
rect 38117 12257 38151 12291
rect 38151 12257 38160 12291
rect 38108 12248 38160 12257
rect 63684 12384 63736 12436
rect 67640 12384 67692 12436
rect 67732 12316 67784 12368
rect 85672 12248 85724 12300
rect 85856 12248 85908 12300
rect 86500 12291 86552 12300
rect 82176 12180 82228 12232
rect 86500 12257 86509 12291
rect 86509 12257 86543 12291
rect 86543 12257 86552 12291
rect 86500 12248 86552 12257
rect 86408 12223 86460 12232
rect 86408 12189 86417 12223
rect 86417 12189 86451 12223
rect 86451 12189 86460 12223
rect 86408 12180 86460 12189
rect 3056 12112 3108 12164
rect 95240 12248 95292 12300
rect 96804 12223 96856 12232
rect 96804 12189 96813 12223
rect 96813 12189 96847 12223
rect 96847 12189 96856 12223
rect 96804 12180 96856 12189
rect 96988 12223 97040 12232
rect 96988 12189 96997 12223
rect 96997 12189 97031 12223
rect 97031 12189 97040 12223
rect 96988 12180 97040 12189
rect 63592 12044 63644 12096
rect 77116 12044 77168 12096
rect 80704 12044 80756 12096
rect 97540 12087 97592 12096
rect 97540 12053 97549 12087
rect 97549 12053 97583 12087
rect 97583 12053 97592 12087
rect 97540 12044 97592 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 65686 11942 65738 11994
rect 65750 11942 65802 11994
rect 65814 11942 65866 11994
rect 65878 11942 65930 11994
rect 96406 11942 96458 11994
rect 96470 11942 96522 11994
rect 96534 11942 96586 11994
rect 96598 11942 96650 11994
rect 3424 11883 3476 11892
rect 3424 11849 3433 11883
rect 3433 11849 3467 11883
rect 3467 11849 3476 11883
rect 3424 11840 3476 11849
rect 30196 11840 30248 11892
rect 97540 11840 97592 11892
rect 20628 11772 20680 11824
rect 48228 11772 48280 11824
rect 80520 11815 80572 11824
rect 80520 11781 80529 11815
rect 80529 11781 80563 11815
rect 80563 11781 80572 11815
rect 80520 11772 80572 11781
rect 80704 11772 80756 11824
rect 85304 11772 85356 11824
rect 3700 11747 3752 11756
rect 3700 11713 3709 11747
rect 3709 11713 3743 11747
rect 3743 11713 3752 11747
rect 3700 11704 3752 11713
rect 3976 11636 4028 11688
rect 12072 11636 12124 11688
rect 17960 11704 18012 11756
rect 35348 11704 35400 11756
rect 41236 11704 41288 11756
rect 53840 11704 53892 11756
rect 77116 11636 77168 11688
rect 17960 11568 18012 11620
rect 27712 11568 27764 11620
rect 33784 11568 33836 11620
rect 37556 11568 37608 11620
rect 44180 11568 44232 11620
rect 51080 11568 51132 11620
rect 52000 11568 52052 11620
rect 80888 11704 80940 11756
rect 31668 11500 31720 11552
rect 80888 11543 80940 11552
rect 80888 11509 80897 11543
rect 80897 11509 80931 11543
rect 80931 11509 80940 11543
rect 80888 11500 80940 11509
rect 96988 11500 97040 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 50326 11398 50378 11450
rect 50390 11398 50442 11450
rect 50454 11398 50506 11450
rect 50518 11398 50570 11450
rect 81046 11398 81098 11450
rect 81110 11398 81162 11450
rect 81174 11398 81226 11450
rect 81238 11398 81290 11450
rect 89352 11296 89404 11348
rect 8760 11228 8812 11280
rect 27160 11203 27212 11212
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 27160 11169 27169 11203
rect 27169 11169 27203 11203
rect 27203 11169 27212 11203
rect 27160 11160 27212 11169
rect 27712 11203 27764 11212
rect 27712 11169 27721 11203
rect 27721 11169 27755 11203
rect 27755 11169 27764 11203
rect 27712 11160 27764 11169
rect 27988 11228 28040 11280
rect 44456 11228 44508 11280
rect 47216 11228 47268 11280
rect 48228 11228 48280 11280
rect 50804 11228 50856 11280
rect 37372 11160 37424 11212
rect 42800 11160 42852 11212
rect 44088 11160 44140 11212
rect 44180 11160 44232 11212
rect 47492 11092 47544 11144
rect 38016 11024 38068 11076
rect 19156 10956 19208 11008
rect 44456 11067 44508 11076
rect 44456 11033 44465 11067
rect 44465 11033 44499 11067
rect 44499 11033 44508 11067
rect 53196 11067 53248 11076
rect 44456 11024 44508 11033
rect 53196 11033 53205 11067
rect 53205 11033 53239 11067
rect 53239 11033 53248 11067
rect 53840 11203 53892 11212
rect 53840 11169 53849 11203
rect 53849 11169 53883 11203
rect 53883 11169 53892 11203
rect 53840 11160 53892 11169
rect 80796 11228 80848 11280
rect 54300 11160 54352 11212
rect 55036 11092 55088 11144
rect 53196 11024 53248 11033
rect 55220 11024 55272 11076
rect 51080 10956 51132 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 65686 10854 65738 10906
rect 65750 10854 65802 10906
rect 65814 10854 65866 10906
rect 65878 10854 65930 10906
rect 96406 10854 96458 10906
rect 96470 10854 96522 10906
rect 96534 10854 96586 10906
rect 96598 10854 96650 10906
rect 5724 10752 5776 10804
rect 16948 10752 17000 10804
rect 55220 10752 55272 10804
rect 3884 10659 3936 10668
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 14464 10684 14516 10736
rect 78864 10684 78916 10736
rect 6184 10616 6236 10668
rect 8576 10616 8628 10668
rect 12900 10659 12952 10668
rect 6644 10548 6696 10600
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 24032 10591 24084 10600
rect 11336 10480 11388 10532
rect 24032 10557 24041 10591
rect 24041 10557 24075 10591
rect 24075 10557 24084 10591
rect 24032 10548 24084 10557
rect 24308 10548 24360 10600
rect 36360 10591 36412 10600
rect 36360 10557 36369 10591
rect 36369 10557 36403 10591
rect 36403 10557 36412 10591
rect 36360 10548 36412 10557
rect 36636 10591 36688 10600
rect 36636 10557 36645 10591
rect 36645 10557 36679 10591
rect 36679 10557 36688 10591
rect 36636 10548 36688 10557
rect 36728 10591 36780 10600
rect 36728 10557 36742 10591
rect 36742 10557 36776 10591
rect 36776 10557 36780 10591
rect 93216 10616 93268 10668
rect 36728 10548 36780 10557
rect 40684 10480 40736 10532
rect 54300 10548 54352 10600
rect 55036 10591 55088 10600
rect 55036 10557 55045 10591
rect 55045 10557 55079 10591
rect 55079 10557 55088 10591
rect 55036 10548 55088 10557
rect 55312 10548 55364 10600
rect 55588 10591 55640 10600
rect 55588 10557 55597 10591
rect 55597 10557 55631 10591
rect 55631 10557 55640 10591
rect 55588 10548 55640 10557
rect 75184 10480 75236 10532
rect 13176 10412 13228 10464
rect 30104 10412 30156 10464
rect 38200 10412 38252 10464
rect 93584 10412 93636 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 50326 10310 50378 10362
rect 50390 10310 50442 10362
rect 50454 10310 50506 10362
rect 50518 10310 50570 10362
rect 81046 10310 81098 10362
rect 81110 10310 81162 10362
rect 81174 10310 81226 10362
rect 81238 10310 81290 10362
rect 4804 10140 4856 10192
rect 20628 10208 20680 10260
rect 40224 10208 40276 10260
rect 61752 10251 61804 10260
rect 61752 10217 61761 10251
rect 61761 10217 61795 10251
rect 61795 10217 61804 10251
rect 61752 10208 61804 10217
rect 62212 10251 62264 10260
rect 62212 10217 62221 10251
rect 62221 10217 62255 10251
rect 62255 10217 62264 10251
rect 62212 10208 62264 10217
rect 35532 10140 35584 10192
rect 39948 10140 40000 10192
rect 17684 10004 17736 10056
rect 62948 10004 63000 10056
rect 63684 10140 63736 10192
rect 63408 10004 63460 10056
rect 80888 10072 80940 10124
rect 93400 10072 93452 10124
rect 63868 10004 63920 10056
rect 92756 10004 92808 10056
rect 17224 9936 17276 9988
rect 17684 9868 17736 9920
rect 17868 9911 17920 9920
rect 17868 9877 17877 9911
rect 17877 9877 17911 9911
rect 17911 9877 17920 9911
rect 17868 9868 17920 9877
rect 24032 9868 24084 9920
rect 24400 9868 24452 9920
rect 63592 9936 63644 9988
rect 94136 9936 94188 9988
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 65686 9766 65738 9818
rect 65750 9766 65802 9818
rect 65814 9766 65866 9818
rect 65878 9766 65930 9818
rect 96406 9766 96458 9818
rect 96470 9766 96522 9818
rect 96534 9766 96586 9818
rect 96598 9766 96650 9818
rect 1952 9664 2004 9716
rect 91008 9664 91060 9716
rect 13176 9528 13228 9580
rect 27068 9528 27120 9580
rect 23204 9460 23256 9512
rect 44364 9460 44416 9512
rect 48964 9596 49016 9648
rect 92572 9596 92624 9648
rect 45284 9503 45336 9512
rect 45284 9469 45293 9503
rect 45293 9469 45327 9503
rect 45327 9469 45336 9503
rect 45284 9460 45336 9469
rect 45652 9460 45704 9512
rect 53104 9528 53156 9580
rect 58072 9528 58124 9580
rect 60188 9528 60240 9580
rect 86408 9528 86460 9580
rect 55588 9460 55640 9512
rect 63408 9460 63460 9512
rect 68284 9460 68336 9512
rect 92848 9460 92900 9512
rect 20536 9392 20588 9444
rect 44456 9392 44508 9444
rect 70768 9392 70820 9444
rect 73804 9392 73856 9444
rect 82820 9392 82872 9444
rect 94044 9435 94096 9444
rect 94044 9401 94053 9435
rect 94053 9401 94087 9435
rect 94087 9401 94096 9435
rect 94044 9392 94096 9401
rect 94412 9392 94464 9444
rect 16672 9324 16724 9376
rect 40868 9324 40920 9376
rect 47584 9324 47636 9376
rect 79508 9324 79560 9376
rect 83464 9324 83516 9376
rect 91284 9324 91336 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 50326 9222 50378 9274
rect 50390 9222 50442 9274
rect 50454 9222 50506 9274
rect 50518 9222 50570 9274
rect 81046 9222 81098 9274
rect 81110 9222 81162 9274
rect 81174 9222 81226 9274
rect 81238 9222 81290 9274
rect 3240 9120 3292 9172
rect 39672 9120 39724 9172
rect 49056 9120 49108 9172
rect 91468 9120 91520 9172
rect 9772 9052 9824 9104
rect 53196 9052 53248 9104
rect 56048 9052 56100 9104
rect 97448 9052 97500 9104
rect 3976 8984 4028 9036
rect 40776 8984 40828 9036
rect 49608 8984 49660 9036
rect 96896 8984 96948 9036
rect 25412 8916 25464 8968
rect 96068 8916 96120 8968
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 65686 8678 65738 8730
rect 65750 8678 65802 8730
rect 65814 8678 65866 8730
rect 65878 8678 65930 8730
rect 96406 8678 96458 8730
rect 96470 8678 96522 8730
rect 96534 8678 96586 8730
rect 96598 8678 96650 8730
rect 4804 8619 4856 8628
rect 4804 8585 4813 8619
rect 4813 8585 4847 8619
rect 4847 8585 4856 8619
rect 4804 8576 4856 8585
rect 11704 8576 11756 8628
rect 12348 8576 12400 8628
rect 60188 8508 60240 8560
rect 32864 8440 32916 8492
rect 4068 8304 4120 8356
rect 75092 8372 75144 8424
rect 50712 8304 50764 8356
rect 63776 8304 63828 8356
rect 67088 8304 67140 8356
rect 20628 8236 20680 8288
rect 22928 8236 22980 8288
rect 23848 8236 23900 8288
rect 25504 8236 25556 8288
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 50326 8134 50378 8186
rect 50390 8134 50442 8186
rect 50454 8134 50506 8186
rect 50518 8134 50570 8186
rect 81046 8134 81098 8186
rect 81110 8134 81162 8186
rect 81174 8134 81226 8186
rect 81238 8134 81290 8186
rect 18880 8032 18932 8084
rect 22836 8032 22888 8084
rect 28908 8032 28960 8084
rect 74816 8032 74868 8084
rect 21456 7964 21508 8016
rect 22100 7964 22152 8016
rect 64420 8007 64472 8016
rect 64420 7973 64429 8007
rect 64429 7973 64463 8007
rect 64463 7973 64472 8007
rect 64420 7964 64472 7973
rect 79140 7964 79192 8016
rect 96804 8032 96856 8084
rect 93860 7939 93912 7948
rect 93860 7905 93869 7939
rect 93869 7905 93903 7939
rect 93903 7905 93912 7939
rect 93860 7896 93912 7905
rect 50988 7828 51040 7880
rect 61384 7828 61436 7880
rect 62764 7871 62816 7880
rect 62764 7837 62773 7871
rect 62773 7837 62807 7871
rect 62807 7837 62816 7871
rect 62764 7828 62816 7837
rect 79232 7828 79284 7880
rect 79692 7828 79744 7880
rect 94412 7939 94464 7948
rect 94412 7905 94421 7939
rect 94421 7905 94455 7939
rect 94455 7905 94464 7939
rect 94412 7896 94464 7905
rect 2964 7760 3016 7812
rect 8760 7692 8812 7744
rect 9128 7692 9180 7744
rect 24492 7760 24544 7812
rect 31116 7760 31168 7812
rect 45100 7760 45152 7812
rect 59360 7760 59412 7812
rect 29920 7692 29972 7744
rect 39764 7692 39816 7744
rect 78496 7760 78548 7812
rect 94412 7692 94464 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 65686 7590 65738 7642
rect 65750 7590 65802 7642
rect 65814 7590 65866 7642
rect 65878 7590 65930 7642
rect 96406 7590 96458 7642
rect 96470 7590 96522 7642
rect 96534 7590 96586 7642
rect 96598 7590 96650 7642
rect 16212 7488 16264 7540
rect 64420 7488 64472 7540
rect 41052 7420 41104 7472
rect 17868 7352 17920 7404
rect 43352 7216 43404 7268
rect 13360 7148 13412 7200
rect 16396 7148 16448 7200
rect 29644 7148 29696 7200
rect 44088 7148 44140 7200
rect 84752 7284 84804 7336
rect 85580 7284 85632 7336
rect 87972 7148 88024 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 50326 7046 50378 7098
rect 50390 7046 50442 7098
rect 50454 7046 50506 7098
rect 50518 7046 50570 7098
rect 81046 7046 81098 7098
rect 81110 7046 81162 7098
rect 81174 7046 81226 7098
rect 81238 7046 81290 7098
rect 2596 6944 2648 6996
rect 94412 6944 94464 6996
rect 13912 6876 13964 6928
rect 16120 6876 16172 6928
rect 45192 6740 45244 6792
rect 38752 6672 38804 6724
rect 48688 6647 48740 6656
rect 48688 6613 48697 6647
rect 48697 6613 48731 6647
rect 48731 6613 48740 6647
rect 59728 6808 59780 6860
rect 62764 6808 62816 6860
rect 98276 6808 98328 6860
rect 53564 6672 53616 6724
rect 60188 6715 60240 6724
rect 60188 6681 60197 6715
rect 60197 6681 60231 6715
rect 60231 6681 60240 6715
rect 60188 6672 60240 6681
rect 56968 6647 57020 6656
rect 48688 6604 48740 6613
rect 56968 6613 56977 6647
rect 56977 6613 57011 6647
rect 57011 6613 57020 6647
rect 56968 6604 57020 6613
rect 59728 6647 59780 6656
rect 59728 6613 59737 6647
rect 59737 6613 59771 6647
rect 59771 6613 59780 6647
rect 59728 6604 59780 6613
rect 84660 6672 84712 6724
rect 78036 6604 78088 6656
rect 97540 6604 97592 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 65686 6502 65738 6554
rect 65750 6502 65802 6554
rect 65814 6502 65866 6554
rect 65878 6502 65930 6554
rect 96406 6502 96458 6554
rect 96470 6502 96522 6554
rect 96534 6502 96586 6554
rect 96598 6502 96650 6554
rect 14188 6400 14240 6452
rect 48688 6400 48740 6452
rect 53840 6400 53892 6452
rect 78036 6400 78088 6452
rect 92112 6443 92164 6452
rect 92112 6409 92121 6443
rect 92121 6409 92155 6443
rect 92155 6409 92164 6443
rect 92112 6400 92164 6409
rect 14004 6264 14056 6316
rect 38752 6264 38804 6316
rect 52460 6196 52512 6248
rect 61936 6196 61988 6248
rect 71044 6196 71096 6248
rect 90456 6196 90508 6248
rect 97632 6239 97684 6248
rect 8392 6128 8444 6180
rect 53564 6128 53616 6180
rect 59636 6128 59688 6180
rect 73528 6128 73580 6180
rect 20720 6060 20772 6112
rect 21732 6060 21784 6112
rect 59728 6060 59780 6112
rect 72700 6060 72752 6112
rect 97632 6205 97641 6239
rect 97641 6205 97675 6239
rect 97675 6205 97684 6239
rect 97632 6196 97684 6205
rect 98828 6128 98880 6180
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 50326 5958 50378 6010
rect 50390 5958 50442 6010
rect 50454 5958 50506 6010
rect 50518 5958 50570 6010
rect 81046 5958 81098 6010
rect 81110 5958 81162 6010
rect 81174 5958 81226 6010
rect 81238 5958 81290 6010
rect 50160 5856 50212 5908
rect 82452 5856 82504 5908
rect 84936 5856 84988 5908
rect 85212 5899 85264 5908
rect 85212 5865 85221 5899
rect 85221 5865 85255 5899
rect 85255 5865 85264 5899
rect 85212 5856 85264 5865
rect 50068 5788 50120 5840
rect 88984 5788 89036 5840
rect 2688 5763 2740 5772
rect 2688 5729 2697 5763
rect 2697 5729 2731 5763
rect 2731 5729 2740 5763
rect 2688 5720 2740 5729
rect 69664 5720 69716 5772
rect 84108 5763 84160 5772
rect 80244 5652 80296 5704
rect 84108 5729 84117 5763
rect 84117 5729 84151 5763
rect 84151 5729 84160 5763
rect 84108 5720 84160 5729
rect 91652 5763 91704 5772
rect 91652 5729 91661 5763
rect 91661 5729 91695 5763
rect 91695 5729 91704 5763
rect 91652 5720 91704 5729
rect 91928 5720 91980 5772
rect 96988 5720 97040 5772
rect 99012 5720 99064 5772
rect 13728 5516 13780 5568
rect 14280 5516 14332 5568
rect 99472 5652 99524 5704
rect 90456 5516 90508 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 65686 5414 65738 5466
rect 65750 5414 65802 5466
rect 65814 5414 65866 5466
rect 65878 5414 65930 5466
rect 96406 5414 96458 5466
rect 96470 5414 96522 5466
rect 96534 5414 96586 5466
rect 96598 5414 96650 5466
rect 6644 5312 6696 5364
rect 68468 5312 68520 5364
rect 82268 5312 82320 5364
rect 85028 5312 85080 5364
rect 16304 5244 16356 5296
rect 46296 5244 46348 5296
rect 67364 5244 67416 5296
rect 80612 5244 80664 5296
rect 3516 5176 3568 5228
rect 1860 5108 1912 5160
rect 7472 5176 7524 5228
rect 16948 5176 17000 5228
rect 17132 5176 17184 5228
rect 35440 5176 35492 5228
rect 3332 5083 3384 5092
rect 3332 5049 3341 5083
rect 3341 5049 3375 5083
rect 3375 5049 3384 5083
rect 3332 5040 3384 5049
rect 480 4972 532 5024
rect 3608 5040 3660 5092
rect 4804 5108 4856 5160
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 10600 5151 10652 5160
rect 10600 5117 10609 5151
rect 10609 5117 10643 5151
rect 10643 5117 10652 5151
rect 10600 5108 10652 5117
rect 11888 5108 11940 5160
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 14280 5151 14332 5160
rect 14280 5117 14289 5151
rect 14289 5117 14323 5151
rect 14323 5117 14332 5151
rect 14280 5108 14332 5117
rect 15476 5151 15528 5160
rect 15476 5117 15485 5151
rect 15485 5117 15519 5151
rect 15519 5117 15528 5151
rect 15476 5108 15528 5117
rect 16856 5108 16908 5160
rect 18604 5151 18656 5160
rect 18604 5117 18613 5151
rect 18613 5117 18647 5151
rect 18647 5117 18656 5151
rect 18604 5108 18656 5117
rect 24400 5151 24452 5160
rect 24400 5117 24409 5151
rect 24409 5117 24443 5151
rect 24443 5117 24452 5151
rect 24400 5108 24452 5117
rect 80520 5151 80572 5160
rect 80520 5117 80529 5151
rect 80529 5117 80563 5151
rect 80563 5117 80572 5151
rect 80520 5108 80572 5117
rect 96252 5108 96304 5160
rect 97816 5151 97868 5160
rect 43444 5040 43496 5092
rect 56968 5040 57020 5092
rect 73712 5040 73764 5092
rect 97816 5117 97825 5151
rect 97825 5117 97859 5151
rect 97859 5117 97868 5151
rect 97816 5108 97868 5117
rect 98460 5040 98512 5092
rect 5172 4972 5224 5024
rect 17224 4972 17276 5024
rect 24584 5015 24636 5024
rect 24584 4981 24593 5015
rect 24593 4981 24627 5015
rect 24627 4981 24636 5015
rect 24584 4972 24636 4981
rect 52460 4972 52512 5024
rect 86960 4972 87012 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 50326 4870 50378 4922
rect 50390 4870 50442 4922
rect 50454 4870 50506 4922
rect 50518 4870 50570 4922
rect 81046 4870 81098 4922
rect 81110 4870 81162 4922
rect 81174 4870 81226 4922
rect 81238 4870 81290 4922
rect 15200 4811 15252 4820
rect 1768 4700 1820 4752
rect 5172 4743 5224 4752
rect 5172 4709 5181 4743
rect 5181 4709 5215 4743
rect 5215 4709 5224 4743
rect 5172 4700 5224 4709
rect 5908 4743 5960 4752
rect 5908 4709 5917 4743
rect 5917 4709 5951 4743
rect 5951 4709 5960 4743
rect 5908 4700 5960 4709
rect 6644 4743 6696 4752
rect 6644 4709 6653 4743
rect 6653 4709 6687 4743
rect 6687 4709 6696 4743
rect 6644 4700 6696 4709
rect 7472 4743 7524 4752
rect 7472 4709 7481 4743
rect 7481 4709 7515 4743
rect 7515 4709 7524 4743
rect 7472 4700 7524 4709
rect 11152 4743 11204 4752
rect 11152 4709 11161 4743
rect 11161 4709 11195 4743
rect 11195 4709 11204 4743
rect 11152 4700 11204 4709
rect 11336 4743 11388 4752
rect 11336 4709 11345 4743
rect 11345 4709 11379 4743
rect 11379 4709 11388 4743
rect 11336 4700 11388 4709
rect 11796 4700 11848 4752
rect 15200 4777 15209 4811
rect 15209 4777 15243 4811
rect 15243 4777 15252 4811
rect 15200 4768 15252 4777
rect 17224 4768 17276 4820
rect 32404 4768 32456 4820
rect 43352 4768 43404 4820
rect 41144 4700 41196 4752
rect 79324 4768 79376 4820
rect 81532 4768 81584 4820
rect 82084 4768 82136 4820
rect 84568 4768 84620 4820
rect 80152 4700 80204 4752
rect 848 4632 900 4684
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 7564 4632 7616 4684
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 12532 4675 12584 4684
rect 12532 4641 12541 4675
rect 12541 4641 12575 4675
rect 12575 4641 12584 4675
rect 12532 4632 12584 4641
rect 15752 4675 15804 4684
rect 5540 4564 5592 4616
rect 6184 4564 6236 4616
rect 12440 4564 12492 4616
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 16120 4632 16172 4684
rect 17132 4632 17184 4684
rect 17316 4632 17368 4684
rect 17960 4632 18012 4684
rect 19432 4632 19484 4684
rect 20352 4632 20404 4684
rect 21088 4632 21140 4684
rect 25044 4632 25096 4684
rect 25688 4632 25740 4684
rect 26424 4632 26476 4684
rect 26884 4632 26936 4684
rect 37280 4675 37332 4684
rect 37280 4641 37289 4675
rect 37289 4641 37323 4675
rect 37323 4641 37332 4675
rect 37280 4632 37332 4641
rect 39120 4675 39172 4684
rect 39120 4641 39129 4675
rect 39129 4641 39163 4675
rect 39163 4641 39172 4675
rect 39120 4632 39172 4641
rect 39672 4632 39724 4684
rect 44088 4632 44140 4684
rect 44548 4675 44600 4684
rect 44548 4641 44557 4675
rect 44557 4641 44591 4675
rect 44591 4641 44600 4675
rect 44548 4632 44600 4641
rect 45836 4632 45888 4684
rect 47032 4675 47084 4684
rect 47032 4641 47041 4675
rect 47041 4641 47075 4675
rect 47075 4641 47084 4675
rect 47032 4632 47084 4641
rect 47584 4632 47636 4684
rect 48228 4632 48280 4684
rect 52552 4675 52604 4684
rect 52552 4641 52561 4675
rect 52561 4641 52595 4675
rect 52595 4641 52604 4675
rect 52552 4632 52604 4641
rect 53104 4632 53156 4684
rect 62856 4675 62908 4684
rect 62856 4641 62865 4675
rect 62865 4641 62899 4675
rect 62899 4641 62908 4675
rect 62856 4632 62908 4641
rect 73804 4675 73856 4684
rect 73804 4641 73813 4675
rect 73813 4641 73847 4675
rect 73847 4641 73856 4675
rect 73804 4632 73856 4641
rect 78772 4675 78824 4684
rect 78772 4641 78781 4675
rect 78781 4641 78815 4675
rect 78815 4641 78824 4675
rect 78772 4632 78824 4641
rect 79324 4632 79376 4684
rect 80060 4675 80112 4684
rect 80060 4641 80069 4675
rect 80069 4641 80103 4675
rect 80103 4641 80112 4675
rect 80060 4632 80112 4641
rect 80796 4675 80848 4684
rect 80796 4641 80805 4675
rect 80805 4641 80839 4675
rect 80839 4641 80848 4675
rect 80796 4632 80848 4641
rect 81440 4675 81492 4684
rect 81440 4641 81449 4675
rect 81449 4641 81483 4675
rect 81483 4641 81492 4675
rect 81440 4632 81492 4641
rect 82912 4675 82964 4684
rect 82912 4641 82921 4675
rect 82921 4641 82955 4675
rect 82955 4641 82964 4675
rect 82912 4632 82964 4641
rect 89720 4632 89772 4684
rect 93400 4675 93452 4684
rect 93400 4641 93409 4675
rect 93409 4641 93443 4675
rect 93443 4641 93452 4675
rect 93400 4632 93452 4641
rect 93952 4632 94004 4684
rect 94596 4632 94648 4684
rect 95240 4632 95292 4684
rect 95792 4632 95844 4684
rect 96712 4632 96764 4684
rect 97264 4675 97316 4684
rect 97264 4641 97273 4675
rect 97273 4641 97307 4675
rect 97307 4641 97316 4675
rect 97264 4632 97316 4641
rect 16304 4564 16356 4616
rect 16948 4564 17000 4616
rect 20720 4564 20772 4616
rect 58532 4564 58584 4616
rect 18512 4496 18564 4548
rect 55864 4496 55916 4548
rect 4620 4428 4672 4480
rect 5080 4471 5132 4480
rect 5080 4437 5089 4471
rect 5089 4437 5123 4471
rect 5123 4437 5132 4471
rect 5080 4428 5132 4437
rect 7472 4428 7524 4480
rect 11612 4428 11664 4480
rect 17132 4428 17184 4480
rect 48504 4428 48556 4480
rect 65156 4471 65208 4480
rect 65156 4437 65165 4471
rect 65165 4437 65199 4471
rect 65199 4437 65208 4471
rect 65156 4428 65208 4437
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 65686 4326 65738 4378
rect 65750 4326 65802 4378
rect 65814 4326 65866 4378
rect 65878 4326 65930 4378
rect 96406 4326 96458 4378
rect 96470 4326 96522 4378
rect 96534 4326 96586 4378
rect 96598 4326 96650 4378
rect 3608 4224 3660 4276
rect 29736 4224 29788 4276
rect 48136 4224 48188 4276
rect 65156 4224 65208 4276
rect 69940 4224 69992 4276
rect 70676 4156 70728 4208
rect 82360 4156 82412 4208
rect 84752 4156 84804 4208
rect 2596 4131 2648 4140
rect 664 4020 716 4072
rect 1492 4020 1544 4072
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 3424 4088 3476 4140
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 2504 3952 2556 4004
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 6368 4020 6420 4072
rect 7656 4063 7708 4072
rect 7656 4029 7665 4063
rect 7665 4029 7699 4063
rect 7699 4029 7708 4063
rect 7656 4020 7708 4029
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 8852 4020 8904 4072
rect 9404 4020 9456 4072
rect 10508 4063 10560 4072
rect 10508 4029 10517 4063
rect 10517 4029 10551 4063
rect 10551 4029 10560 4063
rect 10508 4020 10560 4029
rect 12992 4088 13044 4140
rect 69940 4088 69992 4140
rect 81624 4131 81676 4140
rect 12716 4020 12768 4072
rect 13728 4063 13780 4072
rect 13728 4029 13737 4063
rect 13737 4029 13771 4063
rect 13771 4029 13780 4063
rect 13728 4020 13780 4029
rect 14372 4063 14424 4072
rect 14372 4029 14381 4063
rect 14381 4029 14415 4063
rect 14415 4029 14424 4063
rect 14372 4020 14424 4029
rect 16028 4063 16080 4072
rect 3976 3952 4028 4004
rect 6092 3952 6144 4004
rect 6736 3952 6788 4004
rect 11060 3952 11112 4004
rect 13636 3952 13688 4004
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 17408 4063 17460 4072
rect 17408 4029 17417 4063
rect 17417 4029 17451 4063
rect 17451 4029 17460 4063
rect 17408 4020 17460 4029
rect 18052 4020 18104 4072
rect 18880 4063 18932 4072
rect 18880 4029 18889 4063
rect 18889 4029 18923 4063
rect 18923 4029 18932 4063
rect 18880 4020 18932 4029
rect 19892 4020 19944 4072
rect 20076 4020 20128 4072
rect 22008 4020 22060 4072
rect 22836 4020 22888 4072
rect 23296 4020 23348 4072
rect 23940 4020 23992 4072
rect 24584 4020 24636 4072
rect 25872 4063 25924 4072
rect 25872 4029 25881 4063
rect 25881 4029 25915 4063
rect 25915 4029 25924 4063
rect 25872 4020 25924 4029
rect 26516 4063 26568 4072
rect 26516 4029 26525 4063
rect 26525 4029 26559 4063
rect 26559 4029 26568 4063
rect 26516 4020 26568 4029
rect 27528 4020 27580 4072
rect 28724 4063 28776 4072
rect 28724 4029 28733 4063
rect 28733 4029 28767 4063
rect 28767 4029 28776 4063
rect 28724 4020 28776 4029
rect 29368 4063 29420 4072
rect 29368 4029 29377 4063
rect 29377 4029 29411 4063
rect 29411 4029 29420 4063
rect 29368 4020 29420 4029
rect 30564 4063 30616 4072
rect 30564 4029 30573 4063
rect 30573 4029 30607 4063
rect 30607 4029 30616 4063
rect 30564 4020 30616 4029
rect 31208 4063 31260 4072
rect 31208 4029 31217 4063
rect 31217 4029 31251 4063
rect 31251 4029 31260 4063
rect 31208 4020 31260 4029
rect 31760 4020 31812 4072
rect 33600 4063 33652 4072
rect 33600 4029 33609 4063
rect 33609 4029 33643 4063
rect 33643 4029 33652 4063
rect 33600 4020 33652 4029
rect 34244 4063 34296 4072
rect 34244 4029 34253 4063
rect 34253 4029 34287 4063
rect 34287 4029 34296 4063
rect 34244 4020 34296 4029
rect 34796 4020 34848 4072
rect 35440 4020 35492 4072
rect 36084 4020 36136 4072
rect 36636 4020 36688 4072
rect 37832 4020 37884 4072
rect 38476 4020 38528 4072
rect 39948 4063 40000 4072
rect 39948 4029 39957 4063
rect 39957 4029 39991 4063
rect 39991 4029 40000 4063
rect 39948 4020 40000 4029
rect 40316 4020 40368 4072
rect 40960 4020 41012 4072
rect 41512 4020 41564 4072
rect 42708 4020 42760 4072
rect 46020 4063 46072 4072
rect 20628 3952 20680 4004
rect 43352 3952 43404 4004
rect 1768 3884 1820 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 7196 3884 7248 3936
rect 8024 3884 8076 3936
rect 10508 3884 10560 3936
rect 12348 3884 12400 3936
rect 13452 3884 13504 3936
rect 15936 3884 15988 3936
rect 16396 3884 16448 3936
rect 17776 3884 17828 3936
rect 18328 3884 18380 3936
rect 19064 3884 19116 3936
rect 19984 3884 20036 3936
rect 43996 3884 44048 3936
rect 46020 4029 46029 4063
rect 46029 4029 46063 4063
rect 46063 4029 46072 4063
rect 46020 4020 46072 4029
rect 45192 3952 45244 4004
rect 46388 3884 46440 3936
rect 48412 4020 48464 4072
rect 48872 4020 48924 4072
rect 49608 4020 49660 4072
rect 50160 4020 50212 4072
rect 50804 4020 50856 4072
rect 51448 4020 51500 4072
rect 51908 3952 51960 4004
rect 53748 4020 53800 4072
rect 54300 4020 54352 4072
rect 54944 4020 54996 4072
rect 55588 4020 55640 4072
rect 56140 4020 56192 4072
rect 56784 4020 56836 4072
rect 57428 4020 57480 4072
rect 58624 4020 58676 4072
rect 59176 3952 59228 4004
rect 59820 3952 59872 4004
rect 60464 3884 60516 3936
rect 61016 3952 61068 4004
rect 61752 3952 61804 4004
rect 62304 3884 62356 3936
rect 64144 4020 64196 4072
rect 64788 4020 64840 4072
rect 65984 4020 66036 4072
rect 66536 4063 66588 4072
rect 66536 4029 66545 4063
rect 66545 4029 66579 4063
rect 66579 4029 66588 4063
rect 66536 4020 66588 4029
rect 67180 4063 67232 4072
rect 67180 4029 67189 4063
rect 67189 4029 67223 4063
rect 67223 4029 67232 4063
rect 67180 4020 67232 4029
rect 67732 4020 67784 4072
rect 68468 4063 68520 4072
rect 68468 4029 68477 4063
rect 68477 4029 68511 4063
rect 68511 4029 68520 4063
rect 68468 4020 68520 4029
rect 68928 4020 68980 4072
rect 69572 3952 69624 4004
rect 70768 4020 70820 4072
rect 71412 4020 71464 4072
rect 72056 4020 72108 4072
rect 72608 4020 72660 4072
rect 73252 4020 73304 4072
rect 74448 4020 74500 4072
rect 75092 4020 75144 4072
rect 75736 4020 75788 4072
rect 76380 4020 76432 4072
rect 77024 4020 77076 4072
rect 77668 4020 77720 4072
rect 80244 4063 80296 4072
rect 78128 3952 78180 4004
rect 80244 4029 80253 4063
rect 80253 4029 80287 4063
rect 80287 4029 80296 4063
rect 80244 4020 80296 4029
rect 80336 4020 80388 4072
rect 81624 4097 81633 4131
rect 81633 4097 81667 4131
rect 81667 4097 81676 4131
rect 81624 4088 81676 4097
rect 83556 4088 83608 4140
rect 96896 4131 96948 4140
rect 96896 4097 96905 4131
rect 96905 4097 96939 4131
rect 96939 4097 96948 4131
rect 96896 4088 96948 4097
rect 81992 4020 82044 4072
rect 83648 4063 83700 4072
rect 81808 3952 81860 4004
rect 83648 4029 83657 4063
rect 83657 4029 83691 4063
rect 83691 4029 83700 4063
rect 83648 4020 83700 4029
rect 84200 4020 84252 4072
rect 84844 4020 84896 4072
rect 85396 3952 85448 4004
rect 86684 4020 86736 4072
rect 87236 4020 87288 4072
rect 88524 4063 88576 4072
rect 88524 4029 88533 4063
rect 88533 4029 88567 4063
rect 88567 4029 88576 4063
rect 88524 4020 88576 4029
rect 89076 4020 89128 4072
rect 90272 4020 90324 4072
rect 90916 4020 90968 4072
rect 91560 4020 91612 4072
rect 92112 4020 92164 4072
rect 92756 4020 92808 4072
rect 94136 4063 94188 4072
rect 94136 4029 94145 4063
rect 94145 4029 94179 4063
rect 94179 4029 94188 4063
rect 94136 4020 94188 4029
rect 94780 4063 94832 4072
rect 94780 4029 94789 4063
rect 94789 4029 94823 4063
rect 94823 4029 94832 4063
rect 94780 4020 94832 4029
rect 95976 4063 96028 4072
rect 95976 4029 95985 4063
rect 95985 4029 96019 4063
rect 96019 4029 96028 4063
rect 95976 4020 96028 4029
rect 99288 4020 99340 4072
rect 97448 3952 97500 4004
rect 78220 3884 78272 3936
rect 90180 3884 90232 3936
rect 98000 3927 98052 3936
rect 98000 3893 98009 3927
rect 98009 3893 98043 3927
rect 98043 3893 98052 3927
rect 98000 3884 98052 3893
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 50326 3782 50378 3834
rect 50390 3782 50442 3834
rect 50454 3782 50506 3834
rect 50518 3782 50570 3834
rect 81046 3782 81098 3834
rect 81110 3782 81162 3834
rect 81174 3782 81226 3834
rect 81238 3782 81290 3834
rect 112 3680 164 3732
rect 1124 3680 1176 3732
rect 2964 3723 3016 3732
rect 2964 3689 2973 3723
rect 2973 3689 3007 3723
rect 3007 3689 3016 3723
rect 2964 3680 3016 3689
rect 13360 3680 13412 3732
rect 14924 3680 14976 3732
rect 15752 3680 15804 3732
rect 68652 3680 68704 3732
rect 85028 3723 85080 3732
rect 4068 3612 4120 3664
rect 6276 3612 6328 3664
rect 6460 3655 6512 3664
rect 6460 3621 6469 3655
rect 6469 3621 6503 3655
rect 6503 3621 6512 3655
rect 6460 3612 6512 3621
rect 7380 3612 7432 3664
rect 8576 3612 8628 3664
rect 9772 3655 9824 3664
rect 9772 3621 9781 3655
rect 9781 3621 9815 3655
rect 9815 3621 9824 3655
rect 9772 3612 9824 3621
rect 10784 3612 10836 3664
rect 13268 3655 13320 3664
rect 13268 3621 13277 3655
rect 13277 3621 13311 3655
rect 13311 3621 13320 3655
rect 13268 3612 13320 3621
rect 15384 3655 15436 3664
rect 15384 3621 15393 3655
rect 15393 3621 15427 3655
rect 15427 3621 15436 3655
rect 15384 3612 15436 3621
rect 16488 3655 16540 3664
rect 16488 3621 16497 3655
rect 16497 3621 16531 3655
rect 16531 3621 16540 3655
rect 16488 3612 16540 3621
rect 18236 3612 18288 3664
rect 20168 3612 20220 3664
rect 20996 3655 21048 3664
rect 20996 3621 21005 3655
rect 21005 3621 21039 3655
rect 21039 3621 21048 3655
rect 20996 3612 21048 3621
rect 21916 3612 21968 3664
rect 26976 3612 27028 3664
rect 31576 3612 31628 3664
rect 1124 3544 1176 3596
rect 2228 3544 2280 3596
rect 4712 3544 4764 3596
rect 5448 3544 5500 3596
rect 7196 3587 7248 3596
rect 7196 3553 7205 3587
rect 7205 3553 7239 3587
rect 7239 3553 7248 3587
rect 7196 3544 7248 3553
rect 7748 3544 7800 3596
rect 9128 3544 9180 3596
rect 10232 3544 10284 3596
rect 12072 3544 12124 3596
rect 12624 3544 12676 3596
rect 14464 3544 14516 3596
rect 15016 3544 15068 3596
rect 16304 3544 16356 3596
rect 18144 3544 18196 3596
rect 19984 3587 20036 3596
rect 19984 3553 19993 3587
rect 19993 3553 20027 3587
rect 20027 3553 20036 3587
rect 19984 3544 20036 3553
rect 22192 3544 22244 3596
rect 23480 3544 23532 3596
rect 24676 3544 24728 3596
rect 21364 3476 21416 3528
rect 20812 3408 20864 3460
rect 25228 3408 25280 3460
rect 27068 3544 27120 3596
rect 28080 3587 28132 3596
rect 28080 3553 28089 3587
rect 28089 3553 28123 3587
rect 28123 3553 28132 3587
rect 28080 3544 28132 3553
rect 28908 3587 28960 3596
rect 28908 3553 28917 3587
rect 28917 3553 28951 3587
rect 28951 3553 28960 3587
rect 28908 3544 28960 3553
rect 29920 3544 29972 3596
rect 39764 3612 39816 3664
rect 46756 3655 46808 3664
rect 46756 3621 46765 3655
rect 46765 3621 46799 3655
rect 46799 3621 46808 3655
rect 46756 3612 46808 3621
rect 62396 3612 62448 3664
rect 31944 3544 31996 3596
rect 32496 3544 32548 3596
rect 34428 3587 34480 3596
rect 32956 3476 33008 3528
rect 34428 3553 34437 3587
rect 34437 3553 34471 3587
rect 34471 3553 34480 3587
rect 34428 3544 34480 3553
rect 35624 3544 35676 3596
rect 36820 3587 36872 3596
rect 36820 3553 36829 3587
rect 36829 3553 36863 3587
rect 36863 3553 36872 3587
rect 36820 3544 36872 3553
rect 37464 3587 37516 3596
rect 37464 3553 37473 3587
rect 37473 3553 37507 3587
rect 37507 3553 37516 3587
rect 37464 3544 37516 3553
rect 38108 3587 38160 3596
rect 38108 3553 38117 3587
rect 38117 3553 38151 3587
rect 38151 3553 38160 3587
rect 38108 3544 38160 3553
rect 39304 3587 39356 3596
rect 39304 3553 39313 3587
rect 39313 3553 39347 3587
rect 39347 3553 39356 3587
rect 39304 3544 39356 3553
rect 40500 3544 40552 3596
rect 41696 3587 41748 3596
rect 41696 3553 41705 3587
rect 41705 3553 41739 3587
rect 41739 3553 41748 3587
rect 41696 3544 41748 3553
rect 42340 3587 42392 3596
rect 42340 3553 42349 3587
rect 42349 3553 42383 3587
rect 42383 3553 42392 3587
rect 42340 3544 42392 3553
rect 42984 3587 43036 3596
rect 42984 3553 42993 3587
rect 42993 3553 43027 3587
rect 43027 3553 43036 3587
rect 42984 3544 43036 3553
rect 44824 3587 44876 3596
rect 42156 3476 42208 3528
rect 44824 3553 44833 3587
rect 44833 3553 44867 3587
rect 44867 3553 44876 3587
rect 44824 3544 44876 3553
rect 46296 3587 46348 3596
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 46572 3544 46624 3596
rect 47216 3476 47268 3528
rect 47860 3476 47912 3528
rect 49056 3544 49108 3596
rect 49700 3544 49752 3596
rect 50896 3544 50948 3596
rect 52092 3587 52144 3596
rect 52092 3553 52101 3587
rect 52101 3553 52135 3587
rect 52135 3553 52144 3587
rect 52092 3544 52144 3553
rect 52736 3587 52788 3596
rect 52736 3553 52745 3587
rect 52745 3553 52779 3587
rect 52779 3553 52788 3587
rect 52736 3544 52788 3553
rect 53288 3544 53340 3596
rect 53932 3544 53984 3596
rect 54576 3544 54628 3596
rect 55128 3544 55180 3596
rect 56324 3544 56376 3596
rect 56968 3544 57020 3596
rect 58164 3587 58216 3596
rect 58164 3553 58173 3587
rect 58173 3553 58207 3587
rect 58207 3553 58216 3587
rect 58164 3544 58216 3553
rect 58808 3587 58860 3596
rect 58808 3553 58817 3587
rect 58817 3553 58851 3587
rect 58851 3553 58860 3587
rect 58808 3544 58860 3553
rect 60648 3587 60700 3596
rect 57980 3476 58032 3528
rect 60648 3553 60657 3587
rect 60657 3553 60691 3587
rect 60691 3553 60700 3587
rect 60648 3544 60700 3553
rect 61292 3544 61344 3596
rect 61844 3476 61896 3528
rect 63040 3544 63092 3596
rect 63684 3544 63736 3596
rect 64328 3544 64380 3596
rect 63500 3476 63552 3528
rect 65340 3544 65392 3596
rect 66812 3544 66864 3596
rect 67916 3587 67968 3596
rect 67916 3553 67925 3587
rect 67925 3553 67959 3587
rect 67959 3553 67968 3587
rect 67916 3544 67968 3553
rect 68560 3587 68612 3596
rect 68560 3553 68569 3587
rect 68569 3553 68603 3587
rect 68603 3553 68612 3587
rect 68560 3544 68612 3553
rect 69204 3587 69256 3596
rect 69204 3553 69213 3587
rect 69213 3553 69247 3587
rect 69247 3553 69256 3587
rect 69204 3544 69256 3553
rect 69756 3544 69808 3596
rect 70400 3544 70452 3596
rect 70216 3476 70268 3528
rect 71596 3544 71648 3596
rect 72792 3544 72844 3596
rect 74080 3587 74132 3596
rect 74080 3553 74089 3587
rect 74089 3553 74123 3587
rect 74123 3553 74132 3587
rect 74080 3544 74132 3553
rect 81532 3612 81584 3664
rect 74632 3544 74684 3596
rect 75920 3587 75972 3596
rect 75920 3553 75929 3587
rect 75929 3553 75963 3587
rect 75963 3553 75972 3587
rect 75920 3544 75972 3553
rect 76472 3544 76524 3596
rect 77116 3544 77168 3596
rect 77760 3544 77812 3596
rect 78404 3544 78456 3596
rect 79048 3544 79100 3596
rect 79692 3544 79744 3596
rect 79968 3476 80020 3528
rect 80152 3476 80204 3528
rect 81624 3544 81676 3596
rect 83004 3544 83056 3596
rect 85028 3689 85037 3723
rect 85037 3689 85071 3723
rect 85071 3689 85080 3723
rect 85028 3680 85080 3689
rect 94872 3723 94924 3732
rect 94872 3689 94881 3723
rect 94881 3689 94915 3723
rect 94915 3689 94924 3723
rect 94872 3680 94924 3689
rect 97724 3612 97776 3664
rect 84476 3544 84528 3596
rect 84660 3587 84712 3596
rect 84660 3553 84669 3587
rect 84669 3553 84703 3587
rect 84703 3553 84712 3587
rect 84660 3544 84712 3553
rect 84752 3587 84804 3596
rect 84752 3553 84761 3587
rect 84761 3553 84795 3587
rect 84795 3553 84804 3587
rect 84936 3587 84988 3596
rect 84752 3544 84804 3553
rect 84936 3553 84945 3587
rect 84945 3553 84979 3587
rect 84979 3553 84988 3587
rect 84936 3544 84988 3553
rect 85028 3544 85080 3596
rect 85672 3544 85724 3596
rect 26700 3451 26752 3460
rect 26700 3417 26709 3451
rect 26709 3417 26743 3451
rect 26743 3417 26752 3451
rect 26700 3408 26752 3417
rect 75184 3408 75236 3460
rect 86040 3476 86092 3528
rect 87972 3544 88024 3596
rect 89260 3587 89312 3596
rect 89260 3553 89269 3587
rect 89269 3553 89303 3587
rect 89303 3553 89312 3587
rect 89260 3544 89312 3553
rect 89904 3587 89956 3596
rect 89904 3553 89913 3587
rect 89913 3553 89947 3587
rect 89947 3553 89956 3587
rect 89904 3544 89956 3553
rect 90548 3587 90600 3596
rect 90548 3553 90557 3587
rect 90557 3553 90591 3587
rect 90591 3553 90600 3587
rect 90548 3544 90600 3553
rect 91100 3544 91152 3596
rect 92388 3544 92440 3596
rect 92940 3544 92992 3596
rect 93584 3544 93636 3596
rect 95424 3544 95476 3596
rect 94504 3476 94556 3528
rect 98644 3476 98696 3528
rect 88708 3408 88760 3460
rect 94964 3451 95016 3460
rect 94964 3417 94973 3451
rect 94973 3417 95007 3451
rect 95007 3417 95016 3451
rect 94964 3408 95016 3417
rect 97448 3451 97500 3460
rect 97448 3417 97457 3451
rect 97457 3417 97491 3451
rect 97491 3417 97500 3451
rect 97448 3408 97500 3417
rect 20168 3340 20220 3392
rect 26332 3340 26384 3392
rect 81716 3340 81768 3392
rect 84292 3383 84344 3392
rect 84292 3349 84301 3383
rect 84301 3349 84335 3383
rect 84335 3349 84344 3383
rect 84292 3340 84344 3349
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 65686 3238 65738 3290
rect 65750 3238 65802 3290
rect 65814 3238 65866 3290
rect 65878 3238 65930 3290
rect 96406 3238 96458 3290
rect 96470 3238 96522 3290
rect 96534 3238 96586 3290
rect 96598 3238 96650 3290
rect 9312 3136 9364 3188
rect 13360 3068 13412 3120
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 8760 3000 8812 3052
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 10968 3000 11020 3009
rect 12716 3000 12768 3052
rect 2872 2932 2924 2984
rect 3148 2975 3200 2984
rect 3148 2941 3157 2975
rect 3157 2941 3191 2975
rect 3191 2941 3200 2975
rect 3148 2932 3200 2941
rect 3700 2932 3752 2984
rect 8208 2932 8260 2984
rect 8392 2932 8444 2984
rect 8668 2932 8720 2984
rect 9864 2932 9916 2984
rect 10876 2932 10928 2984
rect 13176 2932 13228 2984
rect 18972 3136 19024 3188
rect 25320 3179 25372 3188
rect 25320 3145 25329 3179
rect 25329 3145 25363 3179
rect 25363 3145 25372 3179
rect 25320 3136 25372 3145
rect 27804 3136 27856 3188
rect 38200 3179 38252 3188
rect 38200 3145 38209 3179
rect 38209 3145 38243 3179
rect 38243 3145 38252 3179
rect 38200 3136 38252 3145
rect 47308 3179 47360 3188
rect 47308 3145 47317 3179
rect 47317 3145 47351 3179
rect 47351 3145 47360 3179
rect 47308 3136 47360 3145
rect 55220 3179 55272 3188
rect 55220 3145 55229 3179
rect 55229 3145 55263 3179
rect 55263 3145 55272 3179
rect 62488 3179 62540 3188
rect 55220 3136 55272 3145
rect 62488 3145 62497 3179
rect 62497 3145 62531 3179
rect 62531 3145 62540 3179
rect 62488 3136 62540 3145
rect 66720 3179 66772 3188
rect 66720 3145 66729 3179
rect 66729 3145 66763 3179
rect 66763 3145 66772 3179
rect 66720 3136 66772 3145
rect 72240 3179 72292 3188
rect 72240 3145 72249 3179
rect 72249 3145 72283 3179
rect 72283 3145 72292 3179
rect 72240 3136 72292 3145
rect 80244 3136 80296 3188
rect 80888 3136 80940 3188
rect 90824 3136 90876 3188
rect 91284 3179 91336 3188
rect 91284 3145 91293 3179
rect 91293 3145 91327 3179
rect 91327 3145 91336 3179
rect 91284 3136 91336 3145
rect 93676 3179 93728 3188
rect 93676 3145 93685 3179
rect 93685 3145 93719 3179
rect 93719 3145 93728 3179
rect 93676 3136 93728 3145
rect 95884 3136 95936 3188
rect 14096 3068 14148 3120
rect 35808 3068 35860 3120
rect 38936 3068 38988 3120
rect 57152 3068 57204 3120
rect 59360 3068 59412 3120
rect 62212 3068 62264 3120
rect 13912 3000 13964 3052
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 17040 3000 17092 3052
rect 19248 3043 19300 3052
rect 19248 3009 19257 3043
rect 19257 3009 19291 3043
rect 19291 3009 19300 3043
rect 19248 3000 19300 3009
rect 20260 3000 20312 3052
rect 20628 3000 20680 3052
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 21456 3000 21508 3009
rect 43536 3000 43588 3052
rect 14004 2975 14056 2984
rect 14004 2941 14013 2975
rect 14013 2941 14047 2975
rect 14047 2941 14056 2975
rect 14004 2932 14056 2941
rect 3976 2907 4028 2916
rect 3976 2873 3985 2907
rect 3985 2873 4019 2907
rect 4019 2873 4028 2907
rect 3976 2864 4028 2873
rect 6000 2864 6052 2916
rect 11428 2864 11480 2916
rect 13912 2864 13964 2916
rect 15752 2932 15804 2984
rect 18788 2932 18840 2984
rect 19340 2932 19392 2984
rect 22652 2975 22704 2984
rect 22652 2941 22661 2975
rect 22661 2941 22695 2975
rect 22695 2941 22704 2975
rect 22652 2932 22704 2941
rect 16212 2864 16264 2916
rect 19248 2864 19300 2916
rect 19432 2864 19484 2916
rect 21640 2864 21692 2916
rect 22928 2864 22980 2916
rect 24032 2932 24084 2984
rect 25320 2932 25372 2984
rect 26332 2975 26384 2984
rect 26332 2941 26341 2975
rect 26341 2941 26375 2975
rect 26375 2941 26384 2975
rect 26332 2932 26384 2941
rect 27804 2932 27856 2984
rect 25504 2907 25556 2916
rect 25504 2873 25513 2907
rect 25513 2873 25547 2907
rect 25547 2873 25556 2907
rect 25504 2864 25556 2873
rect 27712 2864 27764 2916
rect 9220 2796 9272 2848
rect 11244 2796 11296 2848
rect 12532 2796 12584 2848
rect 21364 2796 21416 2848
rect 26056 2796 26108 2848
rect 27344 2796 27396 2848
rect 28356 2796 28408 2848
rect 29552 2932 29604 2984
rect 30104 2932 30156 2984
rect 30748 2932 30800 2984
rect 31392 2932 31444 2984
rect 32588 2932 32640 2984
rect 33232 2932 33284 2984
rect 33784 2932 33836 2984
rect 35532 2932 35584 2984
rect 35256 2907 35308 2916
rect 35256 2873 35265 2907
rect 35265 2873 35299 2907
rect 35299 2873 35308 2907
rect 35256 2864 35308 2873
rect 35348 2864 35400 2916
rect 36268 2932 36320 2984
rect 38200 2932 38252 2984
rect 38660 2932 38712 2984
rect 40224 2975 40276 2984
rect 40224 2941 40233 2975
rect 40233 2941 40267 2975
rect 40267 2941 40276 2975
rect 40224 2932 40276 2941
rect 41604 2932 41656 2984
rect 43720 2975 43772 2984
rect 37648 2864 37700 2916
rect 41328 2907 41380 2916
rect 41328 2873 41337 2907
rect 41337 2873 41371 2907
rect 41371 2873 41380 2907
rect 41328 2864 41380 2873
rect 37096 2796 37148 2848
rect 38752 2796 38804 2848
rect 40132 2796 40184 2848
rect 41144 2796 41196 2848
rect 43720 2941 43729 2975
rect 43729 2941 43763 2975
rect 43763 2941 43772 2975
rect 43720 2932 43772 2941
rect 52368 3000 52420 3052
rect 54852 3000 54904 3052
rect 58348 3000 58400 3052
rect 58440 3000 58492 3052
rect 61568 3000 61620 3052
rect 66168 3000 66220 3052
rect 45744 2975 45796 2984
rect 43168 2864 43220 2916
rect 44180 2864 44232 2916
rect 45744 2941 45753 2975
rect 45753 2941 45787 2975
rect 45787 2941 45796 2975
rect 45744 2932 45796 2941
rect 45560 2907 45612 2916
rect 45560 2873 45569 2907
rect 45569 2873 45603 2907
rect 45603 2873 45612 2907
rect 45560 2864 45612 2873
rect 45376 2796 45428 2848
rect 47308 2932 47360 2984
rect 49516 2932 49568 2984
rect 51264 2975 51316 2984
rect 51264 2941 51273 2975
rect 51273 2941 51307 2975
rect 51307 2941 51316 2975
rect 51264 2932 51316 2941
rect 47400 2907 47452 2916
rect 47400 2873 47409 2907
rect 47409 2873 47443 2907
rect 47443 2873 47452 2907
rect 47400 2864 47452 2873
rect 49240 2907 49292 2916
rect 49240 2873 49249 2907
rect 49249 2873 49283 2907
rect 49283 2873 49292 2907
rect 49240 2864 49292 2873
rect 51080 2907 51132 2916
rect 51080 2873 51089 2907
rect 51089 2873 51123 2907
rect 51123 2873 51132 2907
rect 51080 2864 51132 2873
rect 50160 2796 50212 2848
rect 54116 2975 54168 2984
rect 51448 2864 51500 2916
rect 54116 2941 54125 2975
rect 54125 2941 54159 2975
rect 54159 2941 54168 2975
rect 54116 2932 54168 2941
rect 55220 2932 55272 2984
rect 56876 2932 56928 2984
rect 55312 2907 55364 2916
rect 55312 2873 55321 2907
rect 55321 2873 55355 2907
rect 55355 2873 55364 2907
rect 55312 2864 55364 2873
rect 56600 2907 56652 2916
rect 56600 2873 56609 2907
rect 56609 2873 56643 2907
rect 56643 2873 56652 2907
rect 56600 2864 56652 2873
rect 53564 2796 53616 2848
rect 55864 2796 55916 2848
rect 57612 2932 57664 2984
rect 58992 2864 59044 2916
rect 59544 2932 59596 2984
rect 60096 2932 60148 2984
rect 61660 2975 61712 2984
rect 61660 2941 61669 2975
rect 61669 2941 61703 2975
rect 61703 2941 61712 2975
rect 61660 2932 61712 2941
rect 62488 2932 62540 2984
rect 64696 2975 64748 2984
rect 59636 2864 59688 2916
rect 61476 2907 61528 2916
rect 61476 2873 61485 2907
rect 61485 2873 61519 2907
rect 61519 2873 61528 2907
rect 61476 2864 61528 2873
rect 62672 2907 62724 2916
rect 62672 2873 62681 2907
rect 62681 2873 62715 2907
rect 62715 2873 62724 2907
rect 62672 2864 62724 2873
rect 60188 2796 60240 2848
rect 62120 2796 62172 2848
rect 62488 2796 62540 2848
rect 64696 2941 64705 2975
rect 64705 2941 64739 2975
rect 64739 2941 64748 2975
rect 64696 2932 64748 2941
rect 64880 2932 64932 2984
rect 65524 2932 65576 2984
rect 66720 2932 66772 2984
rect 69940 2975 69992 2984
rect 64512 2907 64564 2916
rect 64512 2873 64521 2907
rect 64521 2873 64555 2907
rect 64555 2873 64564 2907
rect 64512 2864 64564 2873
rect 66904 2907 66956 2916
rect 66904 2873 66913 2907
rect 66913 2873 66947 2907
rect 66947 2873 66956 2907
rect 66904 2864 66956 2873
rect 67364 2864 67416 2916
rect 69940 2941 69949 2975
rect 69949 2941 69983 2975
rect 69983 2941 69992 2975
rect 69940 2932 69992 2941
rect 71044 2932 71096 2984
rect 72240 2932 72292 2984
rect 69388 2864 69440 2916
rect 70584 2907 70636 2916
rect 70584 2873 70593 2907
rect 70593 2873 70627 2907
rect 70627 2873 70636 2907
rect 70584 2864 70636 2873
rect 72424 2907 72476 2916
rect 72424 2873 72433 2907
rect 72433 2873 72467 2907
rect 72467 2873 72476 2907
rect 72424 2864 72476 2873
rect 72240 2796 72292 2848
rect 73436 2932 73488 2984
rect 75184 2975 75236 2984
rect 75184 2941 75193 2975
rect 75193 2941 75227 2975
rect 75227 2941 75236 2975
rect 75184 2932 75236 2941
rect 75276 2932 75328 2984
rect 76840 2975 76892 2984
rect 76840 2941 76849 2975
rect 76849 2941 76883 2975
rect 76883 2941 76892 2975
rect 76840 2932 76892 2941
rect 78220 2932 78272 2984
rect 85120 3068 85172 3120
rect 79968 3000 80020 3052
rect 74908 2864 74960 2916
rect 76656 2907 76708 2916
rect 76656 2873 76665 2907
rect 76665 2873 76699 2907
rect 76699 2873 76708 2907
rect 76656 2864 76708 2873
rect 77944 2907 77996 2916
rect 77944 2873 77953 2907
rect 77953 2873 77987 2907
rect 77987 2873 77996 2907
rect 77944 2864 77996 2873
rect 78036 2864 78088 2916
rect 79784 2864 79836 2916
rect 80428 2907 80480 2916
rect 80428 2873 80437 2907
rect 80437 2873 80471 2907
rect 80471 2873 80480 2907
rect 80428 2864 80480 2873
rect 81348 2932 81400 2984
rect 82360 3000 82412 3052
rect 82912 3000 82964 3052
rect 82636 2932 82688 2984
rect 83280 2932 83332 2984
rect 83924 2932 83976 2984
rect 84384 2864 84436 2916
rect 86224 2932 86276 2984
rect 86868 2932 86920 2984
rect 87512 2932 87564 2984
rect 88156 2932 88208 2984
rect 88800 2932 88852 2984
rect 90824 2932 90876 2984
rect 91284 2932 91336 2984
rect 91744 2932 91796 2984
rect 90088 2864 90140 2916
rect 91008 2864 91060 2916
rect 93676 2932 93728 2984
rect 94412 2932 94464 2984
rect 96068 2975 96120 2984
rect 96068 2941 96077 2975
rect 96077 2941 96111 2975
rect 96111 2941 96120 2975
rect 96068 2932 96120 2941
rect 96804 2932 96856 2984
rect 93124 2907 93176 2916
rect 93124 2873 93133 2907
rect 93133 2873 93167 2907
rect 93167 2873 93176 2907
rect 93124 2864 93176 2873
rect 73620 2796 73672 2848
rect 74724 2796 74776 2848
rect 76104 2796 76156 2848
rect 77300 2796 77352 2848
rect 79232 2839 79284 2848
rect 79232 2805 79241 2839
rect 79241 2805 79275 2839
rect 79275 2805 79284 2839
rect 79232 2796 79284 2805
rect 80336 2796 80388 2848
rect 82176 2796 82228 2848
rect 87052 2796 87104 2848
rect 89628 2796 89680 2848
rect 90364 2796 90416 2848
rect 93768 2864 93820 2916
rect 96252 2864 96304 2916
rect 97540 2907 97592 2916
rect 97540 2873 97549 2907
rect 97549 2873 97583 2907
rect 97583 2873 97592 2907
rect 97540 2864 97592 2873
rect 95608 2796 95660 2848
rect 97724 2796 97776 2848
rect 99840 2796 99892 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 50326 2694 50378 2746
rect 50390 2694 50442 2746
rect 50454 2694 50506 2746
rect 50518 2694 50570 2746
rect 81046 2694 81098 2746
rect 81110 2694 81162 2746
rect 81174 2694 81226 2746
rect 81238 2694 81290 2746
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 22744 2635 22796 2644
rect 22744 2601 22753 2635
rect 22753 2601 22787 2635
rect 22787 2601 22796 2635
rect 22744 2592 22796 2601
rect 2136 2524 2188 2576
rect 3240 2524 3292 2576
rect 4988 2567 5040 2576
rect 4988 2533 4997 2567
rect 4997 2533 5031 2567
rect 5031 2533 5040 2567
rect 4988 2524 5040 2533
rect 7656 2567 7708 2576
rect 7656 2533 7665 2567
rect 7665 2533 7699 2567
rect 7699 2533 7708 2567
rect 7656 2524 7708 2533
rect 10416 2567 10468 2576
rect 10416 2533 10425 2567
rect 10425 2533 10459 2567
rect 10459 2533 10468 2567
rect 10416 2524 10468 2533
rect 11704 2524 11756 2576
rect 12256 2567 12308 2576
rect 12256 2533 12265 2567
rect 12265 2533 12299 2567
rect 12299 2533 12308 2567
rect 12256 2524 12308 2533
rect 13544 2524 13596 2576
rect 13820 2567 13872 2576
rect 13820 2533 13829 2567
rect 13829 2533 13863 2567
rect 13863 2533 13872 2567
rect 13820 2524 13872 2533
rect 15568 2567 15620 2576
rect 15568 2533 15577 2567
rect 15577 2533 15611 2567
rect 15611 2533 15620 2567
rect 15568 2524 15620 2533
rect 16672 2567 16724 2576
rect 16672 2533 16681 2567
rect 16681 2533 16715 2567
rect 16715 2533 16724 2567
rect 16672 2524 16724 2533
rect 18420 2567 18472 2576
rect 18420 2533 18429 2567
rect 18429 2533 18463 2567
rect 18463 2533 18472 2567
rect 18420 2524 18472 2533
rect 19156 2524 19208 2576
rect 20536 2524 20588 2576
rect 21824 2567 21876 2576
rect 21824 2533 21833 2567
rect 21833 2533 21867 2567
rect 21867 2533 21876 2567
rect 21824 2524 21876 2533
rect 26792 2592 26844 2644
rect 23848 2567 23900 2576
rect 23848 2533 23857 2567
rect 23857 2533 23891 2567
rect 23891 2533 23900 2567
rect 23848 2524 23900 2533
rect 24492 2567 24544 2576
rect 24492 2533 24501 2567
rect 24501 2533 24535 2567
rect 24535 2533 24544 2567
rect 24492 2524 24544 2533
rect 25780 2567 25832 2576
rect 25780 2533 25789 2567
rect 25789 2533 25823 2567
rect 25823 2533 25832 2567
rect 25780 2524 25832 2533
rect 28632 2635 28684 2644
rect 28632 2601 28641 2635
rect 28641 2601 28675 2635
rect 28675 2601 28684 2635
rect 28632 2592 28684 2601
rect 28816 2635 28868 2644
rect 28816 2601 28825 2635
rect 28825 2601 28859 2635
rect 28859 2601 28868 2635
rect 29644 2635 29696 2644
rect 28816 2592 28868 2601
rect 29644 2601 29653 2635
rect 29653 2601 29687 2635
rect 29687 2601 29696 2635
rect 29644 2592 29696 2601
rect 30380 2592 30432 2644
rect 31484 2635 31536 2644
rect 31484 2601 31493 2635
rect 31493 2601 31527 2635
rect 31527 2601 31536 2635
rect 31484 2592 31536 2601
rect 34152 2635 34204 2644
rect 34152 2601 34161 2635
rect 34161 2601 34195 2635
rect 34195 2601 34204 2635
rect 34152 2592 34204 2601
rect 32680 2524 32732 2576
rect 33692 2567 33744 2576
rect 33692 2533 33701 2567
rect 33701 2533 33735 2567
rect 33735 2533 33744 2567
rect 33692 2524 33744 2533
rect 35992 2592 36044 2644
rect 36176 2635 36228 2644
rect 36176 2601 36185 2635
rect 36185 2601 36219 2635
rect 36219 2601 36228 2635
rect 36176 2592 36228 2601
rect 36912 2635 36964 2644
rect 36912 2601 36921 2635
rect 36921 2601 36955 2635
rect 36955 2601 36964 2635
rect 36912 2592 36964 2601
rect 39396 2635 39448 2644
rect 37924 2567 37976 2576
rect 37924 2533 37933 2567
rect 37933 2533 37967 2567
rect 37967 2533 37976 2567
rect 37924 2524 37976 2533
rect 38936 2567 38988 2576
rect 38936 2533 38945 2567
rect 38945 2533 38979 2567
rect 38979 2533 38988 2567
rect 38936 2524 38988 2533
rect 39396 2601 39405 2635
rect 39405 2601 39439 2635
rect 39439 2601 39448 2635
rect 39396 2592 39448 2601
rect 40040 2592 40092 2644
rect 41420 2635 41472 2644
rect 39856 2567 39908 2576
rect 39856 2533 39865 2567
rect 39865 2533 39899 2567
rect 39899 2533 39908 2567
rect 39856 2524 39908 2533
rect 41420 2601 41429 2635
rect 41429 2601 41463 2635
rect 41463 2601 41472 2635
rect 41420 2592 41472 2601
rect 45008 2592 45060 2644
rect 49424 2635 49476 2644
rect 49424 2601 49433 2635
rect 49433 2601 49467 2635
rect 49467 2601 49476 2635
rect 49424 2592 49476 2601
rect 296 2456 348 2508
rect 1308 2388 1360 2440
rect 3884 2456 3936 2508
rect 5632 2499 5684 2508
rect 5632 2465 5641 2499
rect 5641 2465 5675 2499
rect 5675 2465 5684 2499
rect 5632 2456 5684 2465
rect 6552 2456 6604 2508
rect 5724 2388 5776 2440
rect 9588 2456 9640 2508
rect 13268 2456 13320 2508
rect 16948 2456 17000 2508
rect 17592 2499 17644 2508
rect 17592 2465 17601 2499
rect 17601 2465 17635 2499
rect 17635 2465 17644 2499
rect 17592 2456 17644 2465
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 24216 2456 24268 2508
rect 14740 2388 14792 2440
rect 23664 2388 23716 2440
rect 27436 2456 27488 2508
rect 33416 2456 33468 2508
rect 38752 2456 38804 2508
rect 42432 2567 42484 2576
rect 42432 2533 42441 2567
rect 42441 2533 42475 2567
rect 42475 2533 42484 2567
rect 42432 2524 42484 2533
rect 43812 2524 43864 2576
rect 44364 2524 44416 2576
rect 45100 2567 45152 2576
rect 45100 2533 45109 2567
rect 45109 2533 45143 2567
rect 45143 2533 45152 2567
rect 45100 2524 45152 2533
rect 45928 2567 45980 2576
rect 45928 2533 45937 2567
rect 45937 2533 45971 2567
rect 45971 2533 45980 2567
rect 45928 2524 45980 2533
rect 48136 2524 48188 2576
rect 48504 2567 48556 2576
rect 48504 2533 48513 2567
rect 48513 2533 48547 2567
rect 48547 2533 48556 2567
rect 48504 2524 48556 2533
rect 50712 2592 50764 2644
rect 54760 2635 54812 2644
rect 50988 2524 51040 2576
rect 54760 2601 54769 2635
rect 54769 2601 54803 2635
rect 54803 2601 54812 2635
rect 54760 2592 54812 2601
rect 52368 2567 52420 2576
rect 52368 2533 52377 2567
rect 52377 2533 52411 2567
rect 52411 2533 52420 2567
rect 52368 2524 52420 2533
rect 53656 2524 53708 2576
rect 53840 2567 53892 2576
rect 53840 2533 53849 2567
rect 53849 2533 53883 2567
rect 53883 2533 53892 2567
rect 53840 2524 53892 2533
rect 58072 2592 58124 2644
rect 55772 2567 55824 2576
rect 55772 2533 55781 2567
rect 55781 2533 55815 2567
rect 55815 2533 55824 2567
rect 55772 2524 55824 2533
rect 56692 2524 56744 2576
rect 57796 2567 57848 2576
rect 57796 2533 57805 2567
rect 57805 2533 57839 2567
rect 57839 2533 57848 2567
rect 57796 2524 57848 2533
rect 58348 2567 58400 2576
rect 58348 2533 58357 2567
rect 58357 2533 58391 2567
rect 58391 2533 58400 2567
rect 58348 2524 58400 2533
rect 60280 2592 60332 2644
rect 59268 2567 59320 2576
rect 59268 2533 59277 2567
rect 59277 2533 59311 2567
rect 59311 2533 59320 2567
rect 59268 2524 59320 2533
rect 62028 2592 62080 2644
rect 66260 2635 66312 2644
rect 66260 2601 66269 2635
rect 66269 2601 66303 2635
rect 66303 2601 66312 2635
rect 68836 2635 68888 2644
rect 66260 2592 66312 2601
rect 61200 2567 61252 2576
rect 61200 2533 61209 2567
rect 61209 2533 61243 2567
rect 61243 2533 61252 2567
rect 61200 2524 61252 2533
rect 61568 2524 61620 2576
rect 61936 2567 61988 2576
rect 61936 2533 61945 2567
rect 61945 2533 61979 2567
rect 61979 2533 61988 2567
rect 61936 2524 61988 2533
rect 63132 2567 63184 2576
rect 63132 2533 63141 2567
rect 63141 2533 63175 2567
rect 63175 2533 63184 2567
rect 63132 2524 63184 2533
rect 64052 2524 64104 2576
rect 66076 2524 66128 2576
rect 68836 2601 68845 2635
rect 68845 2601 68879 2635
rect 68879 2601 68888 2635
rect 68836 2592 68888 2601
rect 67088 2524 67140 2576
rect 68376 2567 68428 2576
rect 68376 2533 68385 2567
rect 68385 2533 68419 2567
rect 68419 2533 68428 2567
rect 68376 2524 68428 2533
rect 69480 2592 69532 2644
rect 70676 2592 70728 2644
rect 71504 2635 71556 2644
rect 71504 2601 71513 2635
rect 71513 2601 71547 2635
rect 71547 2601 71556 2635
rect 74172 2635 74224 2644
rect 71504 2592 71556 2601
rect 74172 2601 74181 2635
rect 74181 2601 74215 2635
rect 74215 2601 74224 2635
rect 74172 2592 74224 2601
rect 72516 2524 72568 2576
rect 74816 2592 74868 2644
rect 77484 2592 77536 2644
rect 78864 2635 78916 2644
rect 30380 2388 30432 2440
rect 32220 2388 32272 2440
rect 34612 2388 34664 2440
rect 38292 2388 38344 2440
rect 46480 2456 46532 2508
rect 49884 2456 49936 2508
rect 54116 2456 54168 2508
rect 59360 2456 59412 2508
rect 62120 2456 62172 2508
rect 8944 2320 8996 2372
rect 9864 2320 9916 2372
rect 15292 2320 15344 2372
rect 21824 2320 21876 2372
rect 23020 2320 23072 2372
rect 24860 2320 24912 2372
rect 27896 2320 27948 2372
rect 28540 2320 28592 2372
rect 29092 2320 29144 2372
rect 29828 2320 29880 2372
rect 31024 2320 31076 2372
rect 32772 2320 32824 2372
rect 8576 2252 8628 2304
rect 22468 2252 22520 2304
rect 31576 2252 31628 2304
rect 33968 2320 34020 2372
rect 38844 2320 38896 2372
rect 36452 2252 36504 2304
rect 40684 2320 40736 2372
rect 42524 2388 42576 2440
rect 43076 2431 43128 2440
rect 43076 2397 43085 2431
rect 43085 2397 43119 2431
rect 43119 2397 43128 2431
rect 43076 2388 43128 2397
rect 43812 2388 43864 2440
rect 48044 2388 48096 2440
rect 51724 2388 51776 2440
rect 55036 2388 55088 2440
rect 59636 2388 59688 2440
rect 63408 2456 63460 2508
rect 66352 2456 66404 2508
rect 69848 2456 69900 2508
rect 63868 2388 63920 2440
rect 67548 2388 67600 2440
rect 71228 2456 71280 2508
rect 76564 2524 76616 2576
rect 77208 2567 77260 2576
rect 77208 2533 77217 2567
rect 77217 2533 77251 2567
rect 77251 2533 77260 2567
rect 77208 2524 77260 2533
rect 77300 2524 77352 2576
rect 78864 2601 78873 2635
rect 78873 2601 78907 2635
rect 78907 2601 78916 2635
rect 79508 2635 79560 2644
rect 78864 2592 78916 2601
rect 79508 2601 79517 2635
rect 79517 2601 79551 2635
rect 79551 2601 79560 2635
rect 79508 2592 79560 2601
rect 73712 2499 73764 2508
rect 73712 2465 73721 2499
rect 73721 2465 73755 2499
rect 73755 2465 73764 2499
rect 73712 2456 73764 2465
rect 74264 2456 74316 2508
rect 80612 2524 80664 2576
rect 82728 2592 82780 2644
rect 84568 2592 84620 2644
rect 88340 2635 88392 2644
rect 88340 2601 88349 2635
rect 88349 2601 88383 2635
rect 88383 2601 88392 2635
rect 89444 2635 89496 2644
rect 88340 2592 88392 2601
rect 82820 2524 82872 2576
rect 85580 2524 85632 2576
rect 85948 2567 86000 2576
rect 85948 2533 85957 2567
rect 85957 2533 85991 2567
rect 85991 2533 86000 2567
rect 85948 2524 86000 2533
rect 86960 2524 87012 2576
rect 87880 2567 87932 2576
rect 87880 2533 87889 2567
rect 87889 2533 87923 2567
rect 87923 2533 87932 2567
rect 87880 2524 87932 2533
rect 89444 2601 89453 2635
rect 89453 2601 89487 2635
rect 89487 2601 89496 2635
rect 89444 2592 89496 2601
rect 89628 2567 89680 2576
rect 89628 2533 89637 2567
rect 89637 2533 89671 2567
rect 89671 2533 89680 2567
rect 89628 2524 89680 2533
rect 90732 2635 90784 2644
rect 90732 2601 90741 2635
rect 90741 2601 90775 2635
rect 90775 2601 90784 2635
rect 90732 2592 90784 2601
rect 91376 2592 91428 2644
rect 92848 2635 92900 2644
rect 91468 2524 91520 2576
rect 92848 2601 92857 2635
rect 92857 2601 92891 2635
rect 92891 2601 92900 2635
rect 92848 2592 92900 2601
rect 94320 2592 94372 2644
rect 95516 2635 95568 2644
rect 93860 2524 93912 2576
rect 95516 2601 95525 2635
rect 95525 2601 95559 2635
rect 95559 2601 95568 2635
rect 95516 2592 95568 2601
rect 96160 2592 96212 2644
rect 97724 2524 97776 2576
rect 95700 2456 95752 2508
rect 73068 2388 73120 2440
rect 77300 2388 77352 2440
rect 81164 2388 81216 2440
rect 81348 2388 81400 2440
rect 84660 2388 84712 2440
rect 86408 2388 86460 2440
rect 46204 2320 46256 2372
rect 41972 2252 42024 2304
rect 46112 2252 46164 2304
rect 47952 2252 48004 2304
rect 50528 2252 50580 2304
rect 51540 2252 51592 2304
rect 52920 2320 52972 2372
rect 57796 2320 57848 2372
rect 55956 2252 56008 2304
rect 60832 2252 60884 2304
rect 63316 2320 63368 2372
rect 66444 2320 66496 2372
rect 69112 2320 69164 2372
rect 71872 2320 71924 2372
rect 75460 2320 75512 2372
rect 65064 2252 65116 2304
rect 70032 2252 70084 2304
rect 74724 2252 74776 2304
rect 78496 2320 78548 2372
rect 84016 2320 84068 2372
rect 85856 2320 85908 2372
rect 87788 2320 87840 2372
rect 82820 2252 82872 2304
rect 83372 2252 83424 2304
rect 85212 2252 85264 2304
rect 88248 2252 88300 2304
rect 91928 2388 91980 2440
rect 91008 2320 91060 2372
rect 93032 2363 93084 2372
rect 93032 2329 93041 2363
rect 93041 2329 93075 2363
rect 93075 2329 93084 2363
rect 93032 2320 93084 2329
rect 90732 2252 90784 2304
rect 94228 2320 94280 2372
rect 99656 2320 99708 2372
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 65686 2150 65738 2202
rect 65750 2150 65802 2202
rect 65814 2150 65866 2202
rect 65878 2150 65930 2202
rect 96406 2150 96458 2202
rect 96470 2150 96522 2202
rect 96534 2150 96586 2202
rect 96598 2150 96650 2202
rect 35992 2048 36044 2100
rect 45652 2048 45704 2100
rect 48688 2048 48740 2100
rect 51540 2048 51592 2100
rect 52276 2048 52328 2100
rect 55036 2048 55088 2100
rect 88892 2048 88944 2100
rect 91008 2048 91060 2100
rect 4344 1844 4396 1896
rect 4804 1844 4856 1896
rect 19800 1844 19852 1896
rect 20076 1844 20128 1896
rect 35072 1504 35124 1556
rect 35348 1504 35400 1556
rect 68744 1436 68796 1488
rect 69848 1436 69900 1488
rect 4528 1368 4580 1420
rect 5632 1368 5684 1420
rect 44364 1368 44416 1420
rect 46112 1368 46164 1420
rect 46848 1368 46900 1420
rect 47952 1368 48004 1420
rect 65708 1368 65760 1420
rect 66444 1368 66496 1420
rect 68192 1368 68244 1420
rect 69112 1368 69164 1420
rect 92572 1368 92624 1420
rect 94228 1368 94280 1420
rect 3976 1300 4028 1352
rect 49792 1300 49844 1352
rect 84292 1300 84344 1352
rect 39488 1164 39540 1216
rect 43076 1164 43128 1216
rect 89536 1164 89588 1216
rect 93032 1164 93084 1216
<< metal2 >>
rect 386 99200 442 100000
rect 1214 99200 1270 100000
rect 2042 99200 2098 100000
rect 2962 99200 3018 100000
rect 3790 99200 3846 100000
rect 4710 99200 4766 100000
rect 5538 99200 5594 100000
rect 6458 99200 6514 100000
rect 7286 99200 7342 100000
rect 8206 99200 8262 100000
rect 9034 99200 9090 100000
rect 9862 99200 9918 100000
rect 10782 99200 10838 100000
rect 11610 99200 11666 100000
rect 12530 99200 12586 100000
rect 13358 99200 13414 100000
rect 14278 99200 14334 100000
rect 15106 99200 15162 100000
rect 16026 99200 16082 100000
rect 16854 99200 16910 100000
rect 17774 99200 17830 100000
rect 18602 99200 18658 100000
rect 19430 99200 19486 100000
rect 20350 99200 20406 100000
rect 21178 99200 21234 100000
rect 22098 99200 22154 100000
rect 22926 99200 22982 100000
rect 23846 99200 23902 100000
rect 24674 99200 24730 100000
rect 25594 99200 25650 100000
rect 26422 99200 26478 100000
rect 27342 99200 27398 100000
rect 28170 99200 28226 100000
rect 28998 99200 29054 100000
rect 29918 99200 29974 100000
rect 30746 99200 30802 100000
rect 31666 99200 31722 100000
rect 32494 99200 32550 100000
rect 33414 99200 33470 100000
rect 34242 99200 34298 100000
rect 35162 99200 35218 100000
rect 35990 99200 36046 100000
rect 36818 99200 36874 100000
rect 37738 99200 37794 100000
rect 38566 99200 38622 100000
rect 39486 99200 39542 100000
rect 40314 99200 40370 100000
rect 41234 99200 41290 100000
rect 42062 99200 42118 100000
rect 42982 99200 43038 100000
rect 43810 99200 43866 100000
rect 44730 99200 44786 100000
rect 45558 99200 45614 100000
rect 46386 99200 46442 100000
rect 47306 99200 47362 100000
rect 48134 99200 48190 100000
rect 49054 99200 49110 100000
rect 49882 99200 49938 100000
rect 50802 99200 50858 100000
rect 51630 99200 51686 100000
rect 52550 99200 52606 100000
rect 53378 99200 53434 100000
rect 54298 99200 54354 100000
rect 55126 99200 55182 100000
rect 55954 99200 56010 100000
rect 56874 99200 56930 100000
rect 57702 99200 57758 100000
rect 58622 99200 58678 100000
rect 59450 99200 59506 100000
rect 60370 99200 60426 100000
rect 61198 99200 61254 100000
rect 62118 99200 62174 100000
rect 62946 99200 63002 100000
rect 63866 99200 63922 100000
rect 64694 99200 64750 100000
rect 65522 99200 65578 100000
rect 66442 99200 66498 100000
rect 67270 99200 67326 100000
rect 68190 99200 68246 100000
rect 69018 99200 69074 100000
rect 69938 99200 69994 100000
rect 70766 99200 70822 100000
rect 71686 99200 71742 100000
rect 72514 99200 72570 100000
rect 73342 99200 73398 100000
rect 74262 99200 74318 100000
rect 75090 99200 75146 100000
rect 76010 99200 76066 100000
rect 76838 99200 76894 100000
rect 77758 99200 77814 100000
rect 78586 99200 78642 100000
rect 79506 99200 79562 100000
rect 80334 99200 80390 100000
rect 81254 99200 81310 100000
rect 82082 99200 82138 100000
rect 82910 99200 82966 100000
rect 83830 99200 83886 100000
rect 84658 99200 84714 100000
rect 85578 99200 85634 100000
rect 86406 99200 86462 100000
rect 87326 99200 87382 100000
rect 88154 99200 88210 100000
rect 89074 99200 89130 100000
rect 89902 99200 89958 100000
rect 90822 99200 90878 100000
rect 91650 99200 91706 100000
rect 92478 99200 92534 100000
rect 93398 99200 93454 100000
rect 94226 99200 94282 100000
rect 95146 99200 95202 100000
rect 95974 99200 96030 100000
rect 96894 99200 96950 100000
rect 97722 99200 97778 100000
rect 98642 99200 98698 100000
rect 99470 99200 99526 100000
rect 400 97170 428 99200
rect 1228 97306 1256 99200
rect 1216 97300 1268 97306
rect 1216 97242 1268 97248
rect 388 97164 440 97170
rect 388 97106 440 97112
rect 1584 96960 1636 96966
rect 1584 96902 1636 96908
rect 1596 54194 1624 96902
rect 2056 96626 2084 99200
rect 2976 97238 3004 99200
rect 3804 97306 3832 99200
rect 3792 97300 3844 97306
rect 3792 97242 3844 97248
rect 2964 97232 3016 97238
rect 2964 97174 3016 97180
rect 2504 97164 2556 97170
rect 2504 97106 2556 97112
rect 2044 96620 2096 96626
rect 2044 96562 2096 96568
rect 2136 96484 2188 96490
rect 2136 96426 2188 96432
rect 2148 96218 2176 96426
rect 2136 96212 2188 96218
rect 2136 96154 2188 96160
rect 2044 94784 2096 94790
rect 2044 94726 2096 94732
rect 1952 87168 2004 87174
rect 1952 87110 2004 87116
rect 1964 72282 1992 87110
rect 1952 72276 2004 72282
rect 1952 72218 2004 72224
rect 1768 54868 1820 54874
rect 1768 54810 1820 54816
rect 1584 54188 1636 54194
rect 1584 54130 1636 54136
rect 1124 50924 1176 50930
rect 1124 50866 1176 50872
rect 480 5024 532 5030
rect 480 4966 532 4972
rect 112 3732 164 3738
rect 112 3674 164 3680
rect 124 800 152 3674
rect 296 2508 348 2514
rect 296 2450 348 2456
rect 308 800 336 2450
rect 492 800 520 4966
rect 848 4684 900 4690
rect 848 4626 900 4632
rect 664 4072 716 4078
rect 664 4014 716 4020
rect 676 800 704 4014
rect 860 800 888 4626
rect 1136 3738 1164 50866
rect 1398 50008 1454 50017
rect 1398 49943 1454 49952
rect 1412 49774 1440 49943
rect 1400 49768 1452 49774
rect 1400 49710 1452 49716
rect 1676 44736 1728 44742
rect 1676 44678 1728 44684
rect 1688 21418 1716 44678
rect 1676 21412 1728 21418
rect 1676 21354 1728 21360
rect 1780 4758 1808 54810
rect 2056 50182 2084 94726
rect 2320 87304 2372 87310
rect 2320 87246 2372 87252
rect 2136 71120 2188 71126
rect 2136 71062 2188 71068
rect 2044 50176 2096 50182
rect 2044 50118 2096 50124
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 9722 1992 10542
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1768 4752 1820 4758
rect 1768 4694 1820 4700
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1124 3732 1176 3738
rect 1124 3674 1176 3680
rect 1124 3596 1176 3602
rect 1124 3538 1176 3544
rect 1136 800 1164 3538
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 1320 800 1348 2382
rect 1504 800 1532 4014
rect 1768 3936 1820 3942
rect 1688 3896 1768 3924
rect 1688 800 1716 3896
rect 1768 3878 1820 3884
rect 1872 800 1900 5102
rect 2148 2582 2176 71062
rect 2332 65686 2360 87246
rect 2412 87236 2464 87242
rect 2412 87178 2464 87184
rect 2320 65680 2372 65686
rect 2320 65622 2372 65628
rect 2424 27674 2452 87178
rect 2412 27668 2464 27674
rect 2412 27610 2464 27616
rect 2516 15978 2544 97106
rect 3056 96960 3108 96966
rect 3056 96902 3108 96908
rect 2596 94988 2648 94994
rect 2596 94930 2648 94936
rect 2608 94858 2636 94930
rect 2596 94852 2648 94858
rect 2596 94794 2648 94800
rect 2608 94586 2636 94794
rect 2596 94580 2648 94586
rect 2596 94522 2648 94528
rect 2596 88936 2648 88942
rect 2596 88878 2648 88884
rect 2608 88466 2636 88878
rect 2596 88460 2648 88466
rect 2596 88402 2648 88408
rect 2872 74792 2924 74798
rect 2872 74734 2924 74740
rect 2884 30666 2912 74734
rect 3068 45558 3096 96902
rect 4220 96860 4516 96880
rect 4276 96858 4300 96860
rect 4356 96858 4380 96860
rect 4436 96858 4460 96860
rect 4298 96806 4300 96858
rect 4362 96806 4374 96858
rect 4436 96806 4438 96858
rect 4276 96804 4300 96806
rect 4356 96804 4380 96806
rect 4436 96804 4460 96806
rect 4220 96784 4516 96804
rect 4724 96626 4752 99200
rect 5552 97170 5580 99200
rect 6472 97306 6500 99200
rect 6460 97300 6512 97306
rect 6460 97242 6512 97248
rect 6184 97232 6236 97238
rect 6184 97174 6236 97180
rect 5540 97164 5592 97170
rect 5540 97106 5592 97112
rect 5724 97096 5776 97102
rect 5724 97038 5776 97044
rect 4896 97028 4948 97034
rect 4896 96970 4948 96976
rect 4712 96620 4764 96626
rect 4712 96562 4764 96568
rect 4804 96484 4856 96490
rect 4804 96426 4856 96432
rect 4220 95772 4516 95792
rect 4276 95770 4300 95772
rect 4356 95770 4380 95772
rect 4436 95770 4460 95772
rect 4298 95718 4300 95770
rect 4362 95718 4374 95770
rect 4436 95718 4438 95770
rect 4276 95716 4300 95718
rect 4356 95716 4380 95718
rect 4436 95716 4460 95718
rect 4220 95696 4516 95716
rect 4220 94684 4516 94704
rect 4276 94682 4300 94684
rect 4356 94682 4380 94684
rect 4436 94682 4460 94684
rect 4298 94630 4300 94682
rect 4362 94630 4374 94682
rect 4436 94630 4438 94682
rect 4276 94628 4300 94630
rect 4356 94628 4380 94630
rect 4436 94628 4460 94630
rect 4220 94608 4516 94628
rect 4220 93596 4516 93616
rect 4276 93594 4300 93596
rect 4356 93594 4380 93596
rect 4436 93594 4460 93596
rect 4298 93542 4300 93594
rect 4362 93542 4374 93594
rect 4436 93542 4438 93594
rect 4276 93540 4300 93542
rect 4356 93540 4380 93542
rect 4436 93540 4460 93542
rect 4220 93520 4516 93540
rect 4220 92508 4516 92528
rect 4276 92506 4300 92508
rect 4356 92506 4380 92508
rect 4436 92506 4460 92508
rect 4298 92454 4300 92506
rect 4362 92454 4374 92506
rect 4436 92454 4438 92506
rect 4276 92452 4300 92454
rect 4356 92452 4380 92454
rect 4436 92452 4460 92454
rect 4220 92432 4516 92452
rect 4220 91420 4516 91440
rect 4276 91418 4300 91420
rect 4356 91418 4380 91420
rect 4436 91418 4460 91420
rect 4298 91366 4300 91418
rect 4362 91366 4374 91418
rect 4436 91366 4438 91418
rect 4276 91364 4300 91366
rect 4356 91364 4380 91366
rect 4436 91364 4460 91366
rect 4220 91344 4516 91364
rect 4220 90332 4516 90352
rect 4276 90330 4300 90332
rect 4356 90330 4380 90332
rect 4436 90330 4460 90332
rect 4298 90278 4300 90330
rect 4362 90278 4374 90330
rect 4436 90278 4438 90330
rect 4276 90276 4300 90278
rect 4356 90276 4380 90278
rect 4436 90276 4460 90278
rect 4220 90256 4516 90276
rect 4068 89888 4120 89894
rect 4068 89830 4120 89836
rect 4080 88942 4108 89830
rect 4220 89244 4516 89264
rect 4276 89242 4300 89244
rect 4356 89242 4380 89244
rect 4436 89242 4460 89244
rect 4298 89190 4300 89242
rect 4362 89190 4374 89242
rect 4436 89190 4438 89242
rect 4276 89188 4300 89190
rect 4356 89188 4380 89190
rect 4436 89188 4460 89190
rect 4220 89168 4516 89188
rect 4068 88936 4120 88942
rect 4068 88878 4120 88884
rect 4220 88156 4516 88176
rect 4276 88154 4300 88156
rect 4356 88154 4380 88156
rect 4436 88154 4460 88156
rect 4298 88102 4300 88154
rect 4362 88102 4374 88154
rect 4436 88102 4438 88154
rect 4276 88100 4300 88102
rect 4356 88100 4380 88102
rect 4436 88100 4460 88102
rect 4220 88080 4516 88100
rect 4220 87068 4516 87088
rect 4276 87066 4300 87068
rect 4356 87066 4380 87068
rect 4436 87066 4460 87068
rect 4298 87014 4300 87066
rect 4362 87014 4374 87066
rect 4436 87014 4438 87066
rect 4276 87012 4300 87014
rect 4356 87012 4380 87014
rect 4436 87012 4460 87014
rect 4220 86992 4516 87012
rect 4220 85980 4516 86000
rect 4276 85978 4300 85980
rect 4356 85978 4380 85980
rect 4436 85978 4460 85980
rect 4298 85926 4300 85978
rect 4362 85926 4374 85978
rect 4436 85926 4438 85978
rect 4276 85924 4300 85926
rect 4356 85924 4380 85926
rect 4436 85924 4460 85926
rect 4220 85904 4516 85924
rect 4220 84892 4516 84912
rect 4276 84890 4300 84892
rect 4356 84890 4380 84892
rect 4436 84890 4460 84892
rect 4298 84838 4300 84890
rect 4362 84838 4374 84890
rect 4436 84838 4438 84890
rect 4276 84836 4300 84838
rect 4356 84836 4380 84838
rect 4436 84836 4460 84838
rect 4220 84816 4516 84836
rect 4220 83804 4516 83824
rect 4276 83802 4300 83804
rect 4356 83802 4380 83804
rect 4436 83802 4460 83804
rect 4298 83750 4300 83802
rect 4362 83750 4374 83802
rect 4436 83750 4438 83802
rect 4276 83748 4300 83750
rect 4356 83748 4380 83750
rect 4436 83748 4460 83750
rect 4220 83728 4516 83748
rect 4220 82716 4516 82736
rect 4276 82714 4300 82716
rect 4356 82714 4380 82716
rect 4436 82714 4460 82716
rect 4298 82662 4300 82714
rect 4362 82662 4374 82714
rect 4436 82662 4438 82714
rect 4276 82660 4300 82662
rect 4356 82660 4380 82662
rect 4436 82660 4460 82662
rect 4220 82640 4516 82660
rect 4220 81628 4516 81648
rect 4276 81626 4300 81628
rect 4356 81626 4380 81628
rect 4436 81626 4460 81628
rect 4298 81574 4300 81626
rect 4362 81574 4374 81626
rect 4436 81574 4438 81626
rect 4276 81572 4300 81574
rect 4356 81572 4380 81574
rect 4436 81572 4460 81574
rect 4220 81552 4516 81572
rect 4220 80540 4516 80560
rect 4276 80538 4300 80540
rect 4356 80538 4380 80540
rect 4436 80538 4460 80540
rect 4298 80486 4300 80538
rect 4362 80486 4374 80538
rect 4436 80486 4438 80538
rect 4276 80484 4300 80486
rect 4356 80484 4380 80486
rect 4436 80484 4460 80486
rect 4220 80464 4516 80484
rect 3976 79552 4028 79558
rect 3976 79494 4028 79500
rect 3988 79150 4016 79494
rect 4220 79452 4516 79472
rect 4276 79450 4300 79452
rect 4356 79450 4380 79452
rect 4436 79450 4460 79452
rect 4298 79398 4300 79450
rect 4362 79398 4374 79450
rect 4436 79398 4438 79450
rect 4276 79396 4300 79398
rect 4356 79396 4380 79398
rect 4436 79396 4460 79398
rect 4220 79376 4516 79396
rect 3976 79144 4028 79150
rect 3976 79086 4028 79092
rect 4528 79144 4580 79150
rect 4712 79144 4764 79150
rect 4580 79092 4660 79098
rect 4528 79086 4660 79092
rect 4712 79086 4764 79092
rect 4540 79070 4660 79086
rect 3884 78532 3936 78538
rect 3884 78474 3936 78480
rect 3332 76492 3384 76498
rect 3332 76434 3384 76440
rect 3056 45552 3108 45558
rect 3056 45494 3108 45500
rect 3344 36922 3372 76434
rect 3700 49156 3752 49162
rect 3700 49098 3752 49104
rect 3332 36916 3384 36922
rect 3332 36858 3384 36864
rect 3516 34196 3568 34202
rect 3516 34138 3568 34144
rect 3056 32360 3108 32366
rect 3056 32302 3108 32308
rect 2872 30660 2924 30666
rect 2872 30602 2924 30608
rect 2504 15972 2556 15978
rect 2504 15914 2556 15920
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2136 2576 2188 2582
rect 2136 2518 2188 2524
rect 2240 1850 2268 3538
rect 2148 1822 2268 1850
rect 2148 800 2176 1822
rect 2332 800 2360 4626
rect 2424 3058 2452 15846
rect 3068 12170 3096 32302
rect 3424 23044 3476 23050
rect 3424 22986 3476 22992
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 3436 11898 3464 22986
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2608 4146 2636 6938
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2516 800 2544 3946
rect 2700 800 2728 5714
rect 2976 3738 3004 7754
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2884 800 2912 2926
rect 3160 800 3188 2926
rect 3252 2582 3280 9114
rect 3528 5522 3556 34138
rect 3712 11762 3740 49098
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3896 10674 3924 78474
rect 4220 78364 4516 78384
rect 4276 78362 4300 78364
rect 4356 78362 4380 78364
rect 4436 78362 4460 78364
rect 4298 78310 4300 78362
rect 4362 78310 4374 78362
rect 4436 78310 4438 78362
rect 4276 78308 4300 78310
rect 4356 78308 4380 78310
rect 4436 78308 4460 78310
rect 4220 78288 4516 78308
rect 4220 77276 4516 77296
rect 4276 77274 4300 77276
rect 4356 77274 4380 77276
rect 4436 77274 4460 77276
rect 4298 77222 4300 77274
rect 4362 77222 4374 77274
rect 4436 77222 4438 77274
rect 4276 77220 4300 77222
rect 4356 77220 4380 77222
rect 4436 77220 4460 77222
rect 4220 77200 4516 77220
rect 4220 76188 4516 76208
rect 4276 76186 4300 76188
rect 4356 76186 4380 76188
rect 4436 76186 4460 76188
rect 4298 76134 4300 76186
rect 4362 76134 4374 76186
rect 4436 76134 4438 76186
rect 4276 76132 4300 76134
rect 4356 76132 4380 76134
rect 4436 76132 4460 76134
rect 4220 76112 4516 76132
rect 4220 75100 4516 75120
rect 4276 75098 4300 75100
rect 4356 75098 4380 75100
rect 4436 75098 4460 75100
rect 4298 75046 4300 75098
rect 4362 75046 4374 75098
rect 4436 75046 4438 75098
rect 4276 75044 4300 75046
rect 4356 75044 4380 75046
rect 4436 75044 4460 75046
rect 4220 75024 4516 75044
rect 4220 74012 4516 74032
rect 4276 74010 4300 74012
rect 4356 74010 4380 74012
rect 4436 74010 4460 74012
rect 4298 73958 4300 74010
rect 4362 73958 4374 74010
rect 4436 73958 4438 74010
rect 4276 73956 4300 73958
rect 4356 73956 4380 73958
rect 4436 73956 4460 73958
rect 4220 73936 4516 73956
rect 4220 72924 4516 72944
rect 4276 72922 4300 72924
rect 4356 72922 4380 72924
rect 4436 72922 4460 72924
rect 4298 72870 4300 72922
rect 4362 72870 4374 72922
rect 4436 72870 4438 72922
rect 4276 72868 4300 72870
rect 4356 72868 4380 72870
rect 4436 72868 4460 72870
rect 4220 72848 4516 72868
rect 4220 71836 4516 71856
rect 4276 71834 4300 71836
rect 4356 71834 4380 71836
rect 4436 71834 4460 71836
rect 4298 71782 4300 71834
rect 4362 71782 4374 71834
rect 4436 71782 4438 71834
rect 4276 71780 4300 71782
rect 4356 71780 4380 71782
rect 4436 71780 4460 71782
rect 4220 71760 4516 71780
rect 4220 70748 4516 70768
rect 4276 70746 4300 70748
rect 4356 70746 4380 70748
rect 4436 70746 4460 70748
rect 4298 70694 4300 70746
rect 4362 70694 4374 70746
rect 4436 70694 4438 70746
rect 4276 70692 4300 70694
rect 4356 70692 4380 70694
rect 4436 70692 4460 70694
rect 4220 70672 4516 70692
rect 4220 69660 4516 69680
rect 4276 69658 4300 69660
rect 4356 69658 4380 69660
rect 4436 69658 4460 69660
rect 4298 69606 4300 69658
rect 4362 69606 4374 69658
rect 4436 69606 4438 69658
rect 4276 69604 4300 69606
rect 4356 69604 4380 69606
rect 4436 69604 4460 69606
rect 4220 69584 4516 69604
rect 4220 68572 4516 68592
rect 4276 68570 4300 68572
rect 4356 68570 4380 68572
rect 4436 68570 4460 68572
rect 4298 68518 4300 68570
rect 4362 68518 4374 68570
rect 4436 68518 4438 68570
rect 4276 68516 4300 68518
rect 4356 68516 4380 68518
rect 4436 68516 4460 68518
rect 4220 68496 4516 68516
rect 4220 67484 4516 67504
rect 4276 67482 4300 67484
rect 4356 67482 4380 67484
rect 4436 67482 4460 67484
rect 4298 67430 4300 67482
rect 4362 67430 4374 67482
rect 4436 67430 4438 67482
rect 4276 67428 4300 67430
rect 4356 67428 4380 67430
rect 4436 67428 4460 67430
rect 4220 67408 4516 67428
rect 4068 67380 4120 67386
rect 4068 67322 4120 67328
rect 4080 67182 4108 67322
rect 4252 67312 4304 67318
rect 4172 67260 4252 67266
rect 4172 67254 4304 67260
rect 4172 67250 4292 67254
rect 4160 67244 4292 67250
rect 4212 67238 4292 67244
rect 4160 67186 4212 67192
rect 3976 67176 4028 67182
rect 3974 67144 3976 67153
rect 4068 67176 4120 67182
rect 4028 67144 4030 67153
rect 4436 67176 4488 67182
rect 4068 67118 4120 67124
rect 4172 67114 4384 67130
rect 4528 67176 4580 67182
rect 4488 67124 4528 67130
rect 4436 67118 4580 67124
rect 3974 67079 4030 67088
rect 4160 67108 4396 67114
rect 4212 67102 4344 67108
rect 4160 67050 4212 67056
rect 4448 67102 4568 67118
rect 4344 67050 4396 67056
rect 4220 66396 4516 66416
rect 4276 66394 4300 66396
rect 4356 66394 4380 66396
rect 4436 66394 4460 66396
rect 4298 66342 4300 66394
rect 4362 66342 4374 66394
rect 4436 66342 4438 66394
rect 4276 66340 4300 66342
rect 4356 66340 4380 66342
rect 4436 66340 4460 66342
rect 4220 66320 4516 66340
rect 4220 65308 4516 65328
rect 4276 65306 4300 65308
rect 4356 65306 4380 65308
rect 4436 65306 4460 65308
rect 4298 65254 4300 65306
rect 4362 65254 4374 65306
rect 4436 65254 4438 65306
rect 4276 65252 4300 65254
rect 4356 65252 4380 65254
rect 4436 65252 4460 65254
rect 4220 65232 4516 65252
rect 4220 64220 4516 64240
rect 4276 64218 4300 64220
rect 4356 64218 4380 64220
rect 4436 64218 4460 64220
rect 4298 64166 4300 64218
rect 4362 64166 4374 64218
rect 4436 64166 4438 64218
rect 4276 64164 4300 64166
rect 4356 64164 4380 64166
rect 4436 64164 4460 64166
rect 4220 64144 4516 64164
rect 4220 63132 4516 63152
rect 4276 63130 4300 63132
rect 4356 63130 4380 63132
rect 4436 63130 4460 63132
rect 4298 63078 4300 63130
rect 4362 63078 4374 63130
rect 4436 63078 4438 63130
rect 4276 63076 4300 63078
rect 4356 63076 4380 63078
rect 4436 63076 4460 63078
rect 4220 63056 4516 63076
rect 4220 62044 4516 62064
rect 4276 62042 4300 62044
rect 4356 62042 4380 62044
rect 4436 62042 4460 62044
rect 4298 61990 4300 62042
rect 4362 61990 4374 62042
rect 4436 61990 4438 62042
rect 4276 61988 4300 61990
rect 4356 61988 4380 61990
rect 4436 61988 4460 61990
rect 4220 61968 4516 61988
rect 4220 60956 4516 60976
rect 4276 60954 4300 60956
rect 4356 60954 4380 60956
rect 4436 60954 4460 60956
rect 4298 60902 4300 60954
rect 4362 60902 4374 60954
rect 4436 60902 4438 60954
rect 4276 60900 4300 60902
rect 4356 60900 4380 60902
rect 4436 60900 4460 60902
rect 4220 60880 4516 60900
rect 4220 59868 4516 59888
rect 4276 59866 4300 59868
rect 4356 59866 4380 59868
rect 4436 59866 4460 59868
rect 4298 59814 4300 59866
rect 4362 59814 4374 59866
rect 4436 59814 4438 59866
rect 4276 59812 4300 59814
rect 4356 59812 4380 59814
rect 4436 59812 4460 59814
rect 4220 59792 4516 59812
rect 4220 58780 4516 58800
rect 4276 58778 4300 58780
rect 4356 58778 4380 58780
rect 4436 58778 4460 58780
rect 4298 58726 4300 58778
rect 4362 58726 4374 58778
rect 4436 58726 4438 58778
rect 4276 58724 4300 58726
rect 4356 58724 4380 58726
rect 4436 58724 4460 58726
rect 4220 58704 4516 58724
rect 4220 57692 4516 57712
rect 4276 57690 4300 57692
rect 4356 57690 4380 57692
rect 4436 57690 4460 57692
rect 4298 57638 4300 57690
rect 4362 57638 4374 57690
rect 4436 57638 4438 57690
rect 4276 57636 4300 57638
rect 4356 57636 4380 57638
rect 4436 57636 4460 57638
rect 4220 57616 4516 57636
rect 4220 56604 4516 56624
rect 4276 56602 4300 56604
rect 4356 56602 4380 56604
rect 4436 56602 4460 56604
rect 4298 56550 4300 56602
rect 4362 56550 4374 56602
rect 4436 56550 4438 56602
rect 4276 56548 4300 56550
rect 4356 56548 4380 56550
rect 4436 56548 4460 56550
rect 4220 56528 4516 56548
rect 4220 55516 4516 55536
rect 4276 55514 4300 55516
rect 4356 55514 4380 55516
rect 4436 55514 4460 55516
rect 4298 55462 4300 55514
rect 4362 55462 4374 55514
rect 4436 55462 4438 55514
rect 4276 55460 4300 55462
rect 4356 55460 4380 55462
rect 4436 55460 4460 55462
rect 4220 55440 4516 55460
rect 4220 54428 4516 54448
rect 4276 54426 4300 54428
rect 4356 54426 4380 54428
rect 4436 54426 4460 54428
rect 4298 54374 4300 54426
rect 4362 54374 4374 54426
rect 4436 54374 4438 54426
rect 4276 54372 4300 54374
rect 4356 54372 4380 54374
rect 4436 54372 4460 54374
rect 4220 54352 4516 54372
rect 4220 53340 4516 53360
rect 4276 53338 4300 53340
rect 4356 53338 4380 53340
rect 4436 53338 4460 53340
rect 4298 53286 4300 53338
rect 4362 53286 4374 53338
rect 4436 53286 4438 53338
rect 4276 53284 4300 53286
rect 4356 53284 4380 53286
rect 4436 53284 4460 53286
rect 4220 53264 4516 53284
rect 4436 53168 4488 53174
rect 4436 53110 4488 53116
rect 3976 52896 4028 52902
rect 3976 52838 4028 52844
rect 3988 52698 4016 52838
rect 3976 52692 4028 52698
rect 3976 52634 4028 52640
rect 4448 52562 4476 53110
rect 4436 52556 4488 52562
rect 4436 52498 4488 52504
rect 4220 52252 4516 52272
rect 4276 52250 4300 52252
rect 4356 52250 4380 52252
rect 4436 52250 4460 52252
rect 4298 52198 4300 52250
rect 4362 52198 4374 52250
rect 4436 52198 4438 52250
rect 4276 52196 4300 52198
rect 4356 52196 4380 52198
rect 4436 52196 4460 52198
rect 4220 52176 4516 52196
rect 4220 51164 4516 51184
rect 4276 51162 4300 51164
rect 4356 51162 4380 51164
rect 4436 51162 4460 51164
rect 4298 51110 4300 51162
rect 4362 51110 4374 51162
rect 4436 51110 4438 51162
rect 4276 51108 4300 51110
rect 4356 51108 4380 51110
rect 4436 51108 4460 51110
rect 4220 51088 4516 51108
rect 4220 50076 4516 50096
rect 4276 50074 4300 50076
rect 4356 50074 4380 50076
rect 4436 50074 4460 50076
rect 4298 50022 4300 50074
rect 4362 50022 4374 50074
rect 4436 50022 4438 50074
rect 4276 50020 4300 50022
rect 4356 50020 4380 50022
rect 4436 50020 4460 50022
rect 4220 50000 4516 50020
rect 4220 48988 4516 49008
rect 4276 48986 4300 48988
rect 4356 48986 4380 48988
rect 4436 48986 4460 48988
rect 4298 48934 4300 48986
rect 4362 48934 4374 48986
rect 4436 48934 4438 48986
rect 4276 48932 4300 48934
rect 4356 48932 4380 48934
rect 4436 48932 4460 48934
rect 4220 48912 4516 48932
rect 4220 47900 4516 47920
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4298 47846 4300 47898
rect 4362 47846 4374 47898
rect 4436 47846 4438 47898
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4220 47824 4516 47844
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4632 44810 4660 79070
rect 4724 78810 4752 79086
rect 4712 78804 4764 78810
rect 4712 78746 4764 78752
rect 4712 67720 4764 67726
rect 4712 67662 4764 67668
rect 4724 67318 4752 67662
rect 4712 67312 4764 67318
rect 4712 67254 4764 67260
rect 4816 45014 4844 96426
rect 4908 48210 4936 96970
rect 5448 94988 5500 94994
rect 5448 94930 5500 94936
rect 5172 94784 5224 94790
rect 5172 94726 5224 94732
rect 5080 89072 5132 89078
rect 5080 89014 5132 89020
rect 5092 85202 5120 89014
rect 5080 85196 5132 85202
rect 5080 85138 5132 85144
rect 5080 75880 5132 75886
rect 5080 75822 5132 75828
rect 5092 69494 5120 75822
rect 5080 69488 5132 69494
rect 5080 69430 5132 69436
rect 4988 67584 5040 67590
rect 4988 67526 5040 67532
rect 5000 55214 5028 67526
rect 5092 60178 5120 69430
rect 5184 67726 5212 94726
rect 5356 76016 5408 76022
rect 5356 75958 5408 75964
rect 5264 69284 5316 69290
rect 5264 69226 5316 69232
rect 5172 67720 5224 67726
rect 5172 67662 5224 67668
rect 5276 67590 5304 69226
rect 5368 69018 5396 75958
rect 5356 69012 5408 69018
rect 5356 68954 5408 68960
rect 5264 67584 5316 67590
rect 5264 67526 5316 67532
rect 5172 67244 5224 67250
rect 5172 67186 5224 67192
rect 5184 67153 5212 67186
rect 5170 67144 5226 67153
rect 5170 67079 5226 67088
rect 5080 60172 5132 60178
rect 5080 60114 5132 60120
rect 5356 57452 5408 57458
rect 5356 57394 5408 57400
rect 5000 55186 5304 55214
rect 4988 52896 5040 52902
rect 4988 52838 5040 52844
rect 5000 52562 5028 52838
rect 5080 52692 5132 52698
rect 5080 52634 5132 52640
rect 4988 52556 5040 52562
rect 4988 52498 5040 52504
rect 4896 48204 4948 48210
rect 4896 48146 4948 48152
rect 4804 45008 4856 45014
rect 4804 44950 4856 44956
rect 4620 44804 4672 44810
rect 4620 44746 4672 44752
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 5092 39506 5120 52634
rect 5080 39500 5132 39506
rect 5080 39442 5132 39448
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4344 32224 4396 32230
rect 4344 32166 4396 32172
rect 4356 32026 4384 32166
rect 4344 32020 4396 32026
rect 4344 31962 4396 31968
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 5276 20398 5304 55186
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3988 11694 4016 18906
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 4816 10198 4844 20334
rect 4988 17264 5040 17270
rect 4988 17206 5040 17212
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3436 5494 3556 5522
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 3344 800 3372 5034
rect 3436 4146 3464 5494
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3528 800 3556 5170
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3620 4282 3648 5034
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3988 4010 4016 8978
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4816 8634 4844 10134
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 4080 3670 4108 8298
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3712 800 3740 2926
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3896 800 3924 2450
rect 3988 1358 4016 2858
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4632 1986 4660 4422
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4172 1958 4660 1986
rect 3976 1352 4028 1358
rect 3976 1294 4028 1300
rect 4172 800 4200 1958
rect 4344 1896 4396 1902
rect 4344 1838 4396 1844
rect 4356 800 4384 1838
rect 4528 1420 4580 1426
rect 4528 1362 4580 1368
rect 4540 800 4568 1362
rect 4724 800 4752 3538
rect 4816 1902 4844 5102
rect 5000 2582 5028 17206
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 4758 5212 4966
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 5092 2258 5120 4422
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5000 2230 5120 2258
rect 4804 1896 4856 1902
rect 4804 1838 4856 1844
rect 5000 800 5028 2230
rect 5184 800 5212 4014
rect 5368 3942 5396 57394
rect 5460 37670 5488 94930
rect 5540 52692 5592 52698
rect 5540 52634 5592 52640
rect 5552 52494 5580 52634
rect 5540 52488 5592 52494
rect 5540 52430 5592 52436
rect 5736 47802 5764 97038
rect 6000 60104 6052 60110
rect 6000 60046 6052 60052
rect 5816 52964 5868 52970
rect 5816 52906 5868 52912
rect 5828 52630 5856 52906
rect 5816 52624 5868 52630
rect 5816 52566 5868 52572
rect 5724 47796 5776 47802
rect 5724 47738 5776 47744
rect 5448 37664 5500 37670
rect 5448 37606 5500 37612
rect 6012 36786 6040 60046
rect 6196 54126 6224 97174
rect 7012 97164 7064 97170
rect 7012 97106 7064 97112
rect 6920 88800 6972 88806
rect 6920 88742 6972 88748
rect 6460 85128 6512 85134
rect 6460 85070 6512 85076
rect 6276 79212 6328 79218
rect 6276 79154 6328 79160
rect 6184 54120 6236 54126
rect 6184 54062 6236 54068
rect 6184 53168 6236 53174
rect 6184 53110 6236 53116
rect 6196 39642 6224 53110
rect 6184 39636 6236 39642
rect 6184 39578 6236 39584
rect 6092 39432 6144 39438
rect 6092 39374 6144 39380
rect 6104 37806 6132 39374
rect 6092 37800 6144 37806
rect 6092 37742 6144 37748
rect 6000 36780 6052 36786
rect 6000 36722 6052 36728
rect 5908 25764 5960 25770
rect 5908 25706 5960 25712
rect 5724 23724 5776 23730
rect 5724 23666 5776 23672
rect 5736 11150 5764 23666
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5736 10810 5764 11086
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5920 4758 5948 25706
rect 6092 12912 6144 12918
rect 6092 12854 6144 12860
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 2774 5488 3538
rect 5368 2746 5488 2774
rect 5368 800 5396 2746
rect 5552 800 5580 4558
rect 6104 4010 6132 12854
rect 6196 10674 6224 39578
rect 6288 16726 6316 79154
rect 6368 66632 6420 66638
rect 6368 66574 6420 66580
rect 6380 32434 6408 66574
rect 6472 62286 6500 85070
rect 6932 82346 6960 88742
rect 6920 82340 6972 82346
rect 6920 82282 6972 82288
rect 7024 81394 7052 97106
rect 7300 96626 7328 99200
rect 7656 97504 7708 97510
rect 7656 97446 7708 97452
rect 7288 96620 7340 96626
rect 7288 96562 7340 96568
rect 7104 96416 7156 96422
rect 7104 96358 7156 96364
rect 7012 81388 7064 81394
rect 7012 81330 7064 81336
rect 6828 79348 6880 79354
rect 6828 79290 6880 79296
rect 6460 62280 6512 62286
rect 6460 62222 6512 62228
rect 6460 59560 6512 59566
rect 6460 59502 6512 59508
rect 6472 52698 6500 59502
rect 6552 58948 6604 58954
rect 6552 58890 6604 58896
rect 6460 52692 6512 52698
rect 6460 52634 6512 52640
rect 6564 52494 6592 58890
rect 6552 52488 6604 52494
rect 6552 52430 6604 52436
rect 6644 45416 6696 45422
rect 6644 45358 6696 45364
rect 6656 44742 6684 45358
rect 6644 44736 6696 44742
rect 6644 44678 6696 44684
rect 6460 36644 6512 36650
rect 6460 36586 6512 36592
rect 6368 32428 6420 32434
rect 6368 32370 6420 32376
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 6380 12434 6408 22714
rect 6288 12406 6408 12434
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5644 1426 5672 2450
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5632 1420 5684 1426
rect 5632 1362 5684 1368
rect 5736 800 5764 2382
rect 6012 800 6040 2858
rect 6196 800 6224 4558
rect 6288 3670 6316 12406
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6380 800 6408 4014
rect 6472 3670 6500 36586
rect 6656 10606 6684 44678
rect 6736 37800 6788 37806
rect 6736 37742 6788 37748
rect 6748 32366 6776 37742
rect 6736 32360 6788 32366
rect 6736 32302 6788 32308
rect 6840 12918 6868 79290
rect 7012 68264 7064 68270
rect 7012 68206 7064 68212
rect 7024 55894 7052 68206
rect 7012 55888 7064 55894
rect 7012 55830 7064 55836
rect 7116 47734 7144 96358
rect 7564 88936 7616 88942
rect 7564 88878 7616 88884
rect 7576 80054 7604 88878
rect 7484 80026 7604 80054
rect 7380 65612 7432 65618
rect 7380 65554 7432 65560
rect 7392 60790 7420 65554
rect 7380 60784 7432 60790
rect 7380 60726 7432 60732
rect 7196 57384 7248 57390
rect 7196 57326 7248 57332
rect 7104 47728 7156 47734
rect 7104 47670 7156 47676
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6656 4758 6684 5306
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6564 800 6592 2450
rect 6748 800 6776 3946
rect 7024 800 7052 5102
rect 7208 3942 7236 57326
rect 7484 47598 7512 80026
rect 7564 52964 7616 52970
rect 7564 52906 7616 52912
rect 7472 47592 7524 47598
rect 7472 47534 7524 47540
rect 7576 39030 7604 52906
rect 7668 52630 7696 97446
rect 8220 97170 8248 99200
rect 9048 97306 9076 99200
rect 9036 97300 9088 97306
rect 9036 97242 9088 97248
rect 8208 97164 8260 97170
rect 8208 97106 8260 97112
rect 8760 97096 8812 97102
rect 8760 97038 8812 97044
rect 8300 90636 8352 90642
rect 8300 90578 8352 90584
rect 7748 88936 7800 88942
rect 7748 88878 7800 88884
rect 7760 88534 7788 88878
rect 7748 88528 7800 88534
rect 7748 88470 7800 88476
rect 8312 87854 8340 90578
rect 8300 87848 8352 87854
rect 8300 87790 8352 87796
rect 8208 81388 8260 81394
rect 8208 81330 8260 81336
rect 8220 80306 8248 81330
rect 8208 80300 8260 80306
rect 8208 80242 8260 80248
rect 7840 53236 7892 53242
rect 7840 53178 7892 53184
rect 7852 52698 7880 53178
rect 7840 52692 7892 52698
rect 7840 52634 7892 52640
rect 7656 52624 7708 52630
rect 7656 52566 7708 52572
rect 7852 52562 7880 52634
rect 7840 52556 7892 52562
rect 7840 52498 7892 52504
rect 8116 52488 8168 52494
rect 8116 52430 8168 52436
rect 7656 45348 7708 45354
rect 7656 45290 7708 45296
rect 7668 44946 7696 45290
rect 8128 45082 8156 52430
rect 8220 47258 8248 80242
rect 8312 74534 8340 87790
rect 8312 74506 8432 74534
rect 8300 63912 8352 63918
rect 8300 63854 8352 63860
rect 8312 50250 8340 63854
rect 8404 63442 8432 74506
rect 8668 64048 8720 64054
rect 8668 63990 8720 63996
rect 8392 63436 8444 63442
rect 8392 63378 8444 63384
rect 8484 57316 8536 57322
rect 8484 57258 8536 57264
rect 8300 50244 8352 50250
rect 8300 50186 8352 50192
rect 8300 48068 8352 48074
rect 8300 48010 8352 48016
rect 8392 48068 8444 48074
rect 8392 48010 8444 48016
rect 8208 47252 8260 47258
rect 8208 47194 8260 47200
rect 8116 45076 8168 45082
rect 8116 45018 8168 45024
rect 7656 44940 7708 44946
rect 7656 44882 7708 44888
rect 7656 43444 7708 43450
rect 7656 43386 7708 43392
rect 7564 39024 7616 39030
rect 7564 38966 7616 38972
rect 7472 27668 7524 27674
rect 7472 27610 7524 27616
rect 7484 26926 7512 27610
rect 7472 26920 7524 26926
rect 7472 26862 7524 26868
rect 7576 26234 7604 38966
rect 7392 26206 7604 26234
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7392 3670 7420 26206
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 4758 7512 5170
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7208 800 7236 3538
rect 7484 2258 7512 4422
rect 7392 2230 7512 2258
rect 7392 800 7420 2230
rect 7576 800 7604 4626
rect 7668 4078 7696 43386
rect 7748 39908 7800 39914
rect 7748 39850 7800 39856
rect 7760 35894 7788 39850
rect 8220 36718 8248 47194
rect 8312 41070 8340 48010
rect 8404 47802 8432 48010
rect 8392 47796 8444 47802
rect 8392 47738 8444 47744
rect 8300 41064 8352 41070
rect 8300 41006 8352 41012
rect 8208 36712 8260 36718
rect 8208 36654 8260 36660
rect 7760 35866 8156 35894
rect 8128 27878 8156 35866
rect 8208 28008 8260 28014
rect 8208 27950 8260 27956
rect 8116 27872 8168 27878
rect 8116 27814 8168 27820
rect 8128 26926 8156 27814
rect 8220 27674 8248 27950
rect 8208 27668 8260 27674
rect 8208 27610 8260 27616
rect 8116 26920 8168 26926
rect 8116 26862 8168 26868
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7760 3924 7788 25842
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8404 4078 8432 6122
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 7668 3896 7788 3924
rect 8024 3936 8076 3942
rect 7668 2582 7696 3896
rect 8024 3878 8076 3884
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7760 800 7788 3538
rect 8036 800 8064 3878
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8220 800 8248 2926
rect 8404 800 8432 2926
rect 8496 2650 8524 57258
rect 8680 50726 8708 63990
rect 8668 50720 8720 50726
rect 8668 50662 8720 50668
rect 8576 36576 8628 36582
rect 8576 36518 8628 36524
rect 8588 16726 8616 36518
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8772 11286 8800 97038
rect 9876 96626 9904 99200
rect 10796 97238 10824 99200
rect 11624 97306 11652 99200
rect 11612 97300 11664 97306
rect 11612 97242 11664 97248
rect 10784 97232 10836 97238
rect 10784 97174 10836 97180
rect 12348 97164 12400 97170
rect 12348 97106 12400 97112
rect 11060 96960 11112 96966
rect 11060 96902 11112 96908
rect 9864 96620 9916 96626
rect 9864 96562 9916 96568
rect 9956 96484 10008 96490
rect 9956 96426 10008 96432
rect 9864 94920 9916 94926
rect 9864 94862 9916 94868
rect 9876 93362 9904 94862
rect 9864 93356 9916 93362
rect 9864 93298 9916 93304
rect 9680 90432 9732 90438
rect 9680 90374 9732 90380
rect 9588 85128 9640 85134
rect 9588 85070 9640 85076
rect 8944 76288 8996 76294
rect 8944 76230 8996 76236
rect 8956 64122 8984 76230
rect 9496 72140 9548 72146
rect 9496 72082 9548 72088
rect 9404 66496 9456 66502
rect 9404 66438 9456 66444
rect 8944 64116 8996 64122
rect 8944 64058 8996 64064
rect 9416 61266 9444 66438
rect 9404 61260 9456 61266
rect 9404 61202 9456 61208
rect 9036 61056 9088 61062
rect 9036 60998 9088 61004
rect 8944 54120 8996 54126
rect 8944 54062 8996 54068
rect 8956 19378 8984 54062
rect 9048 35494 9076 60998
rect 9220 57588 9272 57594
rect 9220 57530 9272 57536
rect 9036 35488 9088 35494
rect 9036 35430 9088 35436
rect 9036 32564 9088 32570
rect 9036 32506 9088 32512
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8956 16658 8984 19314
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 3670 8616 10610
rect 9048 7834 9076 32506
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 9140 24410 9168 24550
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 8680 7806 9076 7834
rect 8576 3664 8628 3670
rect 8576 3606 8628 3612
rect 8680 2990 8708 7806
rect 9140 7750 9168 24346
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 8772 3058 8800 7686
rect 9232 7290 9260 57530
rect 9508 56302 9536 72082
rect 9496 56296 9548 56302
rect 9496 56238 9548 56244
rect 9404 37800 9456 37806
rect 9404 37742 9456 37748
rect 9416 27946 9444 37742
rect 9600 33522 9628 85070
rect 9692 75818 9720 90374
rect 9680 75812 9732 75818
rect 9680 75754 9732 75760
rect 9692 74534 9720 75754
rect 9692 74506 9904 74534
rect 9680 71936 9732 71942
rect 9680 71878 9732 71884
rect 9692 46102 9720 71878
rect 9772 68264 9824 68270
rect 9772 68206 9824 68212
rect 9784 64938 9812 68206
rect 9772 64932 9824 64938
rect 9772 64874 9824 64880
rect 9876 51950 9904 74506
rect 9864 51944 9916 51950
rect 9864 51886 9916 51892
rect 9968 46918 9996 96426
rect 10876 95396 10928 95402
rect 10876 95338 10928 95344
rect 10692 93832 10744 93838
rect 10692 93774 10744 93780
rect 10704 93362 10732 93774
rect 10692 93356 10744 93362
rect 10692 93298 10744 93304
rect 10140 87236 10192 87242
rect 10140 87178 10192 87184
rect 10046 85232 10102 85241
rect 10046 85167 10048 85176
rect 10100 85167 10102 85176
rect 10048 85138 10100 85144
rect 10048 68332 10100 68338
rect 10048 68274 10100 68280
rect 9956 46912 10008 46918
rect 9956 46854 10008 46860
rect 9680 46096 9732 46102
rect 9680 46038 9732 46044
rect 10060 39914 10088 68274
rect 10152 61266 10180 87178
rect 10508 85332 10560 85338
rect 10508 85274 10560 85280
rect 10520 85202 10548 85274
rect 10600 85264 10652 85270
rect 10600 85206 10652 85212
rect 10508 85196 10560 85202
rect 10508 85138 10560 85144
rect 10232 85128 10284 85134
rect 10232 85070 10284 85076
rect 10324 85128 10376 85134
rect 10324 85070 10376 85076
rect 10244 80646 10272 85070
rect 10232 80640 10284 80646
rect 10232 80582 10284 80588
rect 10336 79286 10364 85070
rect 10612 84998 10640 85206
rect 10600 84992 10652 84998
rect 10600 84934 10652 84940
rect 10324 79280 10376 79286
rect 10324 79222 10376 79228
rect 10140 61260 10192 61266
rect 10140 61202 10192 61208
rect 10336 45490 10364 79222
rect 10704 68270 10732 93298
rect 10784 87440 10836 87446
rect 10784 87382 10836 87388
rect 10692 68264 10744 68270
rect 10692 68206 10744 68212
rect 10508 67040 10560 67046
rect 10508 66982 10560 66988
rect 10324 45484 10376 45490
rect 10324 45426 10376 45432
rect 10416 43988 10468 43994
rect 10416 43930 10468 43936
rect 10048 39908 10100 39914
rect 10048 39850 10100 39856
rect 9956 36780 10008 36786
rect 9956 36722 10008 36728
rect 9588 33516 9640 33522
rect 9588 33458 9640 33464
rect 9968 30802 9996 36722
rect 10048 35284 10100 35290
rect 10048 35226 10100 35232
rect 9956 30796 10008 30802
rect 9956 30738 10008 30744
rect 9772 30660 9824 30666
rect 9772 30602 9824 30608
rect 9404 27940 9456 27946
rect 9404 27882 9456 27888
rect 9784 23866 9812 30602
rect 9956 24880 10008 24886
rect 9956 24822 10008 24828
rect 9968 24274 9996 24822
rect 10060 24818 10088 35226
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 8956 7262 9260 7290
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8588 800 8616 2246
rect 8864 800 8892 4014
rect 8956 2378 8984 7262
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 9140 1850 9168 3538
rect 9324 3194 9352 13262
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9048 1822 9168 1850
rect 9048 800 9076 1822
rect 9232 800 9260 2790
rect 9416 800 9444 4014
rect 9784 3670 9812 9046
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9876 2990 9904 16050
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9600 800 9628 2450
rect 9864 2372 9916 2378
rect 9864 2314 9916 2320
rect 9876 800 9904 2314
rect 10060 800 10088 4626
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10244 800 10272 3538
rect 10428 2582 10456 43930
rect 10520 38350 10548 66982
rect 10692 57248 10744 57254
rect 10692 57190 10744 57196
rect 10704 57050 10732 57190
rect 10692 57044 10744 57050
rect 10692 56986 10744 56992
rect 10600 52080 10652 52086
rect 10600 52022 10652 52028
rect 10612 51882 10640 52022
rect 10600 51876 10652 51882
rect 10600 51818 10652 51824
rect 10508 38344 10560 38350
rect 10508 38286 10560 38292
rect 10612 30802 10640 51818
rect 10600 30796 10652 30802
rect 10600 30738 10652 30744
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10508 25696 10560 25702
rect 10508 25638 10560 25644
rect 10520 24818 10548 25638
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10612 24698 10640 25978
rect 10520 24670 10640 24698
rect 10520 4078 10548 24670
rect 10600 24608 10652 24614
rect 10600 24550 10652 24556
rect 10612 23798 10640 24550
rect 10600 23792 10652 23798
rect 10600 23734 10652 23740
rect 10796 20534 10824 87382
rect 10888 39982 10916 95338
rect 11072 55690 11100 96902
rect 11704 93152 11756 93158
rect 11704 93094 11756 93100
rect 11612 79008 11664 79014
rect 11612 78950 11664 78956
rect 11520 78668 11572 78674
rect 11520 78610 11572 78616
rect 11532 78198 11560 78610
rect 11520 78192 11572 78198
rect 11520 78134 11572 78140
rect 11336 69896 11388 69902
rect 11336 69838 11388 69844
rect 11152 56160 11204 56166
rect 11152 56102 11204 56108
rect 11060 55684 11112 55690
rect 11060 55626 11112 55632
rect 10876 39976 10928 39982
rect 10876 39918 10928 39924
rect 10968 38412 11020 38418
rect 10968 38354 11020 38360
rect 10876 38208 10928 38214
rect 10876 38150 10928 38156
rect 10888 33658 10916 38150
rect 10980 37874 11008 38354
rect 10968 37868 11020 37874
rect 10968 37810 11020 37816
rect 10876 33652 10928 33658
rect 10876 33594 10928 33600
rect 11060 24132 11112 24138
rect 11060 24074 11112 24080
rect 11072 23594 11100 24074
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 10784 20528 10836 20534
rect 10784 20470 10836 20476
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 10520 1986 10548 3878
rect 10428 1958 10548 1986
rect 10428 800 10456 1958
rect 10612 800 10640 5102
rect 10796 3670 10824 20470
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 10980 3058 11008 13466
rect 11164 4758 11192 56102
rect 11244 46164 11296 46170
rect 11244 46106 11296 46112
rect 11256 38282 11284 46106
rect 11348 38486 11376 69838
rect 11624 60734 11652 78950
rect 11532 60706 11652 60734
rect 11428 52896 11480 52902
rect 11428 52838 11480 52844
rect 11336 38480 11388 38486
rect 11336 38422 11388 38428
rect 11244 38276 11296 38282
rect 11244 38218 11296 38224
rect 11244 38004 11296 38010
rect 11244 37946 11296 37952
rect 11256 37330 11284 37946
rect 11244 37324 11296 37330
rect 11244 37266 11296 37272
rect 11440 13394 11468 52838
rect 11532 37330 11560 60706
rect 11612 55956 11664 55962
rect 11612 55898 11664 55904
rect 11624 46170 11652 55898
rect 11612 46164 11664 46170
rect 11612 46106 11664 46112
rect 11520 37324 11572 37330
rect 11520 37266 11572 37272
rect 11716 27062 11744 93094
rect 11796 91792 11848 91798
rect 11796 91734 11848 91740
rect 11808 48006 11836 91734
rect 12072 86760 12124 86766
rect 12072 86702 12124 86708
rect 12084 86358 12112 86702
rect 12072 86352 12124 86358
rect 12072 86294 12124 86300
rect 11888 64932 11940 64938
rect 11888 64874 11940 64880
rect 11796 48000 11848 48006
rect 11796 47942 11848 47948
rect 11900 46714 11928 64874
rect 11980 63232 12032 63238
rect 11980 63174 12032 63180
rect 11888 46708 11940 46714
rect 11888 46650 11940 46656
rect 11888 40928 11940 40934
rect 11888 40870 11940 40876
rect 11796 35624 11848 35630
rect 11796 35566 11848 35572
rect 11704 27056 11756 27062
rect 11704 26998 11756 27004
rect 11808 26234 11836 35566
rect 11900 30870 11928 40870
rect 11888 30864 11940 30870
rect 11888 30806 11940 30812
rect 11808 26206 11928 26234
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11348 4758 11376 10474
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10888 800 10916 2926
rect 11072 800 11100 3946
rect 11428 2916 11480 2922
rect 11428 2858 11480 2864
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 11256 800 11284 2790
rect 11440 800 11468 2858
rect 11624 800 11652 4422
rect 11716 2582 11744 8570
rect 11808 4758 11836 24074
rect 11900 16574 11928 26206
rect 11992 21690 12020 63174
rect 12164 51808 12216 51814
rect 12164 51750 12216 51756
rect 12072 42764 12124 42770
rect 12072 42706 12124 42712
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11900 16546 12020 16574
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 11900 800 11928 5102
rect 11992 4146 12020 16546
rect 12084 11694 12112 42706
rect 12176 32366 12204 51750
rect 12256 49768 12308 49774
rect 12256 49710 12308 49716
rect 12268 42770 12296 49710
rect 12256 42764 12308 42770
rect 12256 42706 12308 42712
rect 12360 41274 12388 97106
rect 12544 96626 12572 99200
rect 13372 97170 13400 99200
rect 14292 97238 14320 99200
rect 14280 97232 14332 97238
rect 14280 97174 14332 97180
rect 13360 97164 13412 97170
rect 13360 97106 13412 97112
rect 15016 97164 15068 97170
rect 15016 97106 15068 97112
rect 14832 97096 14884 97102
rect 14832 97038 14884 97044
rect 14464 96688 14516 96694
rect 14464 96630 14516 96636
rect 12532 96620 12584 96626
rect 12532 96562 12584 96568
rect 12624 96484 12676 96490
rect 12624 96426 12676 96432
rect 12532 86896 12584 86902
rect 12532 86838 12584 86844
rect 12440 75404 12492 75410
rect 12440 75346 12492 75352
rect 12452 74662 12480 75346
rect 12440 74656 12492 74662
rect 12440 74598 12492 74604
rect 12544 64874 12572 86838
rect 12636 75410 12664 96426
rect 13820 88868 13872 88874
rect 13820 88810 13872 88816
rect 13832 88466 13860 88810
rect 13820 88460 13872 88466
rect 13820 88402 13872 88408
rect 12808 86760 12860 86766
rect 12808 86702 12860 86708
rect 12820 83638 12848 86702
rect 12808 83632 12860 83638
rect 12808 83574 12860 83580
rect 12900 80640 12952 80646
rect 12900 80582 12952 80588
rect 12912 79218 12940 80582
rect 12900 79212 12952 79218
rect 12900 79154 12952 79160
rect 12624 75404 12676 75410
rect 12624 75346 12676 75352
rect 12452 64846 12572 64874
rect 12348 41268 12400 41274
rect 12348 41210 12400 41216
rect 12360 40934 12388 41210
rect 12348 40928 12400 40934
rect 12348 40870 12400 40876
rect 12452 37806 12480 64846
rect 12440 37800 12492 37806
rect 12440 37742 12492 37748
rect 12164 32360 12216 32366
rect 12164 32302 12216 32308
rect 12348 32020 12400 32026
rect 12348 31962 12400 31968
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12268 18698 12296 19246
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12176 13394 12204 13806
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 12084 800 12112 3538
rect 12268 2582 12296 18634
rect 12360 8634 12388 31962
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12624 27056 12676 27062
rect 12624 26998 12676 27004
rect 12636 26858 12664 26998
rect 12624 26852 12676 26858
rect 12624 26794 12676 26800
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12544 13326 12572 13398
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 12360 1986 12388 3878
rect 12268 1958 12388 1986
rect 12268 800 12296 1958
rect 12452 800 12480 4558
rect 12544 2854 12572 4626
rect 12636 3924 12664 26794
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12728 23730 12756 24686
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12728 4078 12756 21422
rect 12820 20262 12848 27474
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12912 10674 12940 79154
rect 13820 76424 13872 76430
rect 13820 76366 13872 76372
rect 13832 75834 13860 76366
rect 13740 75806 13860 75834
rect 13740 74866 13768 75806
rect 13728 74860 13780 74866
rect 13728 74802 13780 74808
rect 13740 72690 13768 74802
rect 13728 72684 13780 72690
rect 13728 72626 13780 72632
rect 13544 72616 13596 72622
rect 13544 72558 13596 72564
rect 13556 67114 13584 72558
rect 13636 72480 13688 72486
rect 13636 72422 13688 72428
rect 13648 67250 13676 72422
rect 13636 67244 13688 67250
rect 13636 67186 13688 67192
rect 13544 67108 13596 67114
rect 13544 67050 13596 67056
rect 13740 66502 13768 72626
rect 13728 66496 13780 66502
rect 13728 66438 13780 66444
rect 14280 64048 14332 64054
rect 14280 63990 14332 63996
rect 12992 62756 13044 62762
rect 12992 62698 13044 62704
rect 13004 62354 13032 62698
rect 12992 62348 13044 62354
rect 12992 62290 13044 62296
rect 13176 62348 13228 62354
rect 13176 62290 13228 62296
rect 12992 49768 13044 49774
rect 12992 49710 13044 49716
rect 13004 49162 13032 49710
rect 12992 49156 13044 49162
rect 12992 49098 13044 49104
rect 12992 40044 13044 40050
rect 12992 39986 13044 39992
rect 13004 37398 13032 39986
rect 12992 37392 13044 37398
rect 12992 37334 13044 37340
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 13188 10470 13216 62290
rect 14004 57384 14056 57390
rect 14004 57326 14056 57332
rect 13452 50788 13504 50794
rect 13452 50730 13504 50736
rect 13464 49978 13492 50730
rect 13452 49972 13504 49978
rect 13452 49914 13504 49920
rect 13636 46368 13688 46374
rect 13636 46310 13688 46316
rect 13648 46034 13676 46310
rect 13636 46028 13688 46034
rect 13636 45970 13688 45976
rect 14016 32842 14044 57326
rect 14004 32836 14056 32842
rect 14004 32778 14056 32784
rect 13268 25968 13320 25974
rect 13268 25910 13320 25916
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12636 3896 12756 3924
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12636 800 12664 3538
rect 12728 3058 12756 3896
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 13004 1986 13032 4082
rect 12912 1958 13032 1986
rect 12912 800 12940 1958
rect 13096 800 13124 5102
rect 13188 2990 13216 9522
rect 13280 3670 13308 25910
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13648 15434 13676 15914
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13648 14958 13676 15370
rect 14004 15156 14056 15162
rect 14004 15098 14056 15104
rect 14016 14958 14044 15098
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 3738 13400 7142
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13372 3126 13400 3674
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13280 800 13308 2450
rect 13464 800 13492 3878
rect 13556 2582 13584 14418
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13740 4078 13768 5510
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 13648 2122 13676 3946
rect 13832 2582 13860 14826
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 13924 3058 13952 6870
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14016 2990 14044 6258
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13648 2094 13768 2122
rect 13740 800 13768 2094
rect 13924 800 13952 2858
rect 14108 800 14136 3062
rect 14200 3058 14228 6394
rect 14292 5574 14320 63990
rect 14372 41132 14424 41138
rect 14372 41074 14424 41080
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14292 800 14320 5102
rect 14384 4078 14412 41074
rect 14476 10742 14504 96630
rect 14556 96212 14608 96218
rect 14556 96154 14608 96160
rect 14568 16590 14596 96154
rect 14740 91520 14792 91526
rect 14740 91462 14792 91468
rect 14648 85332 14700 85338
rect 14648 85274 14700 85280
rect 14660 85241 14688 85274
rect 14646 85232 14702 85241
rect 14646 85167 14702 85176
rect 14648 82272 14700 82278
rect 14648 82214 14700 82220
rect 14660 40050 14688 82214
rect 14752 62966 14780 91462
rect 14740 62960 14792 62966
rect 14740 62902 14792 62908
rect 14740 61192 14792 61198
rect 14740 61134 14792 61140
rect 14752 53650 14780 61134
rect 14844 55078 14872 97038
rect 14924 94988 14976 94994
rect 14924 94930 14976 94936
rect 14832 55072 14884 55078
rect 14832 55014 14884 55020
rect 14740 53644 14792 53650
rect 14740 53586 14792 53592
rect 14752 47122 14780 53586
rect 14936 51066 14964 94930
rect 15028 75886 15056 97106
rect 15120 96626 15148 99200
rect 16040 97238 16068 99200
rect 16304 97640 16356 97646
rect 16304 97582 16356 97588
rect 16028 97232 16080 97238
rect 16028 97174 16080 97180
rect 16212 96960 16264 96966
rect 16212 96902 16264 96908
rect 15108 96620 15160 96626
rect 15108 96562 15160 96568
rect 15384 94988 15436 94994
rect 15384 94930 15436 94936
rect 15108 88868 15160 88874
rect 15108 88810 15160 88816
rect 15120 76430 15148 88810
rect 15108 76424 15160 76430
rect 15108 76366 15160 76372
rect 15016 75880 15068 75886
rect 15016 75822 15068 75828
rect 15028 57322 15056 75822
rect 15108 62144 15160 62150
rect 15108 62086 15160 62092
rect 15016 57316 15068 57322
rect 15016 57258 15068 57264
rect 15120 55418 15148 62086
rect 15108 55412 15160 55418
rect 15108 55354 15160 55360
rect 15016 53576 15068 53582
rect 15016 53518 15068 53524
rect 14924 51060 14976 51066
rect 14924 51002 14976 51008
rect 15028 49298 15056 53518
rect 15108 49904 15160 49910
rect 15108 49846 15160 49852
rect 15016 49292 15068 49298
rect 15016 49234 15068 49240
rect 14740 47116 14792 47122
rect 14740 47058 14792 47064
rect 14832 46708 14884 46714
rect 14832 46650 14884 46656
rect 14844 46510 14872 46650
rect 14740 46504 14792 46510
rect 14740 46446 14792 46452
rect 14832 46504 14884 46510
rect 14832 46446 14884 46452
rect 14752 46170 14780 46446
rect 14740 46164 14792 46170
rect 14740 46106 14792 46112
rect 14844 41002 14872 46446
rect 15120 45286 15148 49846
rect 15396 48754 15424 94930
rect 15476 94784 15528 94790
rect 15476 94726 15528 94732
rect 15488 63306 15516 94726
rect 16120 88596 16172 88602
rect 16120 88538 16172 88544
rect 15844 88460 15896 88466
rect 15844 88402 15896 88408
rect 15752 87780 15804 87786
rect 15752 87722 15804 87728
rect 15764 64874 15792 87722
rect 15856 74534 15884 88402
rect 15856 74506 16068 74534
rect 15936 69828 15988 69834
rect 15936 69770 15988 69776
rect 15948 68882 15976 69770
rect 15936 68876 15988 68882
rect 15936 68818 15988 68824
rect 15948 68338 15976 68818
rect 15936 68332 15988 68338
rect 15936 68274 15988 68280
rect 15672 64846 15792 64874
rect 15476 63300 15528 63306
rect 15476 63242 15528 63248
rect 15672 62898 15700 64846
rect 16040 64530 16068 74506
rect 16132 68202 16160 88538
rect 16224 71194 16252 96902
rect 16316 96762 16344 97582
rect 16868 97306 16896 99200
rect 16856 97300 16908 97306
rect 16856 97242 16908 97248
rect 17684 97164 17736 97170
rect 17684 97106 17736 97112
rect 16304 96756 16356 96762
rect 16304 96698 16356 96704
rect 16304 88936 16356 88942
rect 16304 88878 16356 88884
rect 16316 88602 16344 88878
rect 16304 88596 16356 88602
rect 16304 88538 16356 88544
rect 17592 78736 17644 78742
rect 17420 78684 17592 78690
rect 17420 78678 17644 78684
rect 17040 78668 17092 78674
rect 17040 78610 17092 78616
rect 17132 78668 17184 78674
rect 17132 78610 17184 78616
rect 17420 78662 17632 78678
rect 17052 78470 17080 78610
rect 17040 78464 17092 78470
rect 17040 78406 17092 78412
rect 17052 78130 17080 78406
rect 17040 78124 17092 78130
rect 17040 78066 17092 78072
rect 16304 73908 16356 73914
rect 16304 73850 16356 73856
rect 16212 71188 16264 71194
rect 16212 71130 16264 71136
rect 16120 68196 16172 68202
rect 16120 68138 16172 68144
rect 16132 67794 16160 68138
rect 16120 67788 16172 67794
rect 16120 67730 16172 67736
rect 16028 64524 16080 64530
rect 16028 64466 16080 64472
rect 15660 62892 15712 62898
rect 15660 62834 15712 62840
rect 15476 62756 15528 62762
rect 15476 62698 15528 62704
rect 15488 58886 15516 62698
rect 15672 59158 15700 62834
rect 15844 62348 15896 62354
rect 15844 62290 15896 62296
rect 15660 59152 15712 59158
rect 15660 59094 15712 59100
rect 15476 58880 15528 58886
rect 15476 58822 15528 58828
rect 15384 48748 15436 48754
rect 15384 48690 15436 48696
rect 15108 45280 15160 45286
rect 15108 45222 15160 45228
rect 14832 40996 14884 41002
rect 14832 40938 14884 40944
rect 14648 40044 14700 40050
rect 14648 39986 14700 39992
rect 15200 30796 15252 30802
rect 15200 30738 15252 30744
rect 14924 27464 14976 27470
rect 14924 27406 14976 27412
rect 14936 24750 14964 27406
rect 14924 24744 14976 24750
rect 14924 24686 14976 24692
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14568 15162 14596 16526
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14476 800 14504 3538
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14752 800 14780 2382
rect 14936 800 14964 3674
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15028 1850 15056 3538
rect 15120 3058 15148 22578
rect 15212 4826 15240 30738
rect 15488 28626 15516 58822
rect 15672 28626 15700 59094
rect 15476 28620 15528 28626
rect 15476 28562 15528 28568
rect 15660 28620 15712 28626
rect 15660 28562 15712 28568
rect 15488 27538 15516 28562
rect 15476 27532 15528 27538
rect 15476 27474 15528 27480
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15396 3670 15424 21490
rect 15856 20398 15884 62290
rect 15936 54256 15988 54262
rect 15936 54198 15988 54204
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 15028 1822 15148 1850
rect 15120 800 15148 1822
rect 15304 800 15332 2314
rect 15488 800 15516 5102
rect 15580 2582 15608 15098
rect 15948 15026 15976 54198
rect 16040 38418 16068 64466
rect 16120 49088 16172 49094
rect 16120 49030 16172 49036
rect 16028 38412 16080 38418
rect 16028 38354 16080 38360
rect 16040 36718 16068 38354
rect 16028 36712 16080 36718
rect 16028 36654 16080 36660
rect 16028 27600 16080 27606
rect 16028 27542 16080 27548
rect 16040 27130 16068 27542
rect 16028 27124 16080 27130
rect 16028 27066 16080 27072
rect 16028 24880 16080 24886
rect 16028 24822 16080 24828
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15764 3738 15792 4626
rect 16040 4078 16068 24822
rect 16132 23322 16160 49030
rect 16212 42084 16264 42090
rect 16212 42026 16264 42032
rect 16224 32570 16252 42026
rect 16212 32564 16264 32570
rect 16212 32506 16264 32512
rect 16212 29708 16264 29714
rect 16212 29650 16264 29656
rect 16224 29034 16252 29650
rect 16212 29028 16264 29034
rect 16212 28970 16264 28976
rect 16120 23316 16172 23322
rect 16120 23258 16172 23264
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16132 6934 16160 19994
rect 16224 12434 16252 28970
rect 16316 13870 16344 73850
rect 16488 68808 16540 68814
rect 16488 68750 16540 68756
rect 16500 46374 16528 68750
rect 16948 67720 17000 67726
rect 16948 67662 17000 67668
rect 16488 46368 16540 46374
rect 16488 46310 16540 46316
rect 16500 43382 16528 46310
rect 16960 46170 16988 67662
rect 16948 46164 17000 46170
rect 16948 46106 17000 46112
rect 16488 43376 16540 43382
rect 16488 43318 16540 43324
rect 16960 42158 16988 46106
rect 16948 42152 17000 42158
rect 16948 42094 17000 42100
rect 17040 37800 17092 37806
rect 17040 37742 17092 37748
rect 16488 29028 16540 29034
rect 16488 28970 16540 28976
rect 16396 23180 16448 23186
rect 16396 23122 16448 23128
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16224 12406 16344 12434
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15752 2984 15804 2990
rect 15752 2926 15804 2932
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 15764 800 15792 2926
rect 15948 800 15976 3878
rect 16132 800 16160 4626
rect 16224 2922 16252 7482
rect 16316 5302 16344 12406
rect 16408 7206 16436 23122
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16304 5296 16356 5302
rect 16304 5238 16356 5244
rect 16316 4622 16344 5238
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16316 800 16344 3538
rect 16408 1986 16436 3878
rect 16500 3670 16528 28970
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16960 10810 16988 13126
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 16684 2582 16712 9318
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16868 2666 16896 5102
rect 16960 4622 16988 5170
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 17052 3058 17080 37742
rect 17144 27538 17172 78610
rect 17420 78606 17448 78662
rect 17408 78600 17460 78606
rect 17408 78542 17460 78548
rect 17224 78464 17276 78470
rect 17224 78406 17276 78412
rect 17132 27532 17184 27538
rect 17132 27474 17184 27480
rect 17236 26450 17264 78406
rect 17696 66570 17724 97106
rect 17788 96626 17816 99200
rect 18616 97238 18644 99200
rect 19444 97306 19472 99200
rect 19580 97404 19876 97424
rect 19636 97402 19660 97404
rect 19716 97402 19740 97404
rect 19796 97402 19820 97404
rect 19658 97350 19660 97402
rect 19722 97350 19734 97402
rect 19796 97350 19798 97402
rect 19636 97348 19660 97350
rect 19716 97348 19740 97350
rect 19796 97348 19820 97350
rect 19580 97328 19876 97348
rect 20364 97322 20392 99200
rect 19432 97300 19484 97306
rect 20364 97294 20484 97322
rect 19432 97242 19484 97248
rect 18604 97232 18656 97238
rect 18604 97174 18656 97180
rect 20352 97164 20404 97170
rect 20352 97106 20404 97112
rect 18788 96960 18840 96966
rect 18788 96902 18840 96908
rect 17776 96620 17828 96626
rect 17776 96562 17828 96568
rect 17868 96484 17920 96490
rect 17868 96426 17920 96432
rect 17776 78668 17828 78674
rect 17776 78610 17828 78616
rect 17788 75342 17816 78610
rect 17776 75336 17828 75342
rect 17776 75278 17828 75284
rect 17880 73914 17908 96426
rect 17960 88936 18012 88942
rect 17960 88878 18012 88884
rect 17868 73908 17920 73914
rect 17868 73850 17920 73856
rect 17684 66564 17736 66570
rect 17684 66506 17736 66512
rect 17408 49768 17460 49774
rect 17408 49710 17460 49716
rect 17316 45484 17368 45490
rect 17316 45426 17368 45432
rect 17328 45014 17356 45426
rect 17316 45008 17368 45014
rect 17316 44950 17368 44956
rect 17420 42838 17448 49710
rect 17696 45554 17724 66506
rect 17868 52692 17920 52698
rect 17868 52634 17920 52640
rect 17880 49978 17908 52634
rect 17868 49972 17920 49978
rect 17868 49914 17920 49920
rect 17512 45526 17724 45554
rect 17408 42832 17460 42838
rect 17408 42774 17460 42780
rect 17224 26444 17276 26450
rect 17224 26386 17276 26392
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17144 17202 17172 17478
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17236 9994 17264 14826
rect 17224 9988 17276 9994
rect 17224 9930 17276 9936
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17144 4690 17172 5170
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17236 4826 17264 4966
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16776 2638 16896 2666
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 16408 1958 16528 1986
rect 16500 800 16528 1958
rect 16776 800 16804 2638
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 16960 800 16988 2450
rect 17144 800 17172 4422
rect 17328 800 17356 4626
rect 17420 4078 17448 42774
rect 17512 37942 17540 45526
rect 17972 45098 18000 88878
rect 18696 63232 18748 63238
rect 18696 63174 18748 63180
rect 18144 59560 18196 59566
rect 18144 59502 18196 59508
rect 18156 45354 18184 59502
rect 18604 59424 18656 59430
rect 18604 59366 18656 59372
rect 18616 48822 18644 59366
rect 18708 53038 18736 63174
rect 18800 57526 18828 96902
rect 19580 96316 19876 96336
rect 19636 96314 19660 96316
rect 19716 96314 19740 96316
rect 19796 96314 19820 96316
rect 19658 96262 19660 96314
rect 19722 96262 19734 96314
rect 19796 96262 19798 96314
rect 19636 96260 19660 96262
rect 19716 96260 19740 96262
rect 19796 96260 19820 96262
rect 19580 96240 19876 96260
rect 19580 95228 19876 95248
rect 19636 95226 19660 95228
rect 19716 95226 19740 95228
rect 19796 95226 19820 95228
rect 19658 95174 19660 95226
rect 19722 95174 19734 95226
rect 19796 95174 19798 95226
rect 19636 95172 19660 95174
rect 19716 95172 19740 95174
rect 19796 95172 19820 95174
rect 19580 95152 19876 95172
rect 19580 94140 19876 94160
rect 19636 94138 19660 94140
rect 19716 94138 19740 94140
rect 19796 94138 19820 94140
rect 19658 94086 19660 94138
rect 19722 94086 19734 94138
rect 19796 94086 19798 94138
rect 19636 94084 19660 94086
rect 19716 94084 19740 94086
rect 19796 94084 19820 94086
rect 19580 94064 19876 94084
rect 19580 93052 19876 93072
rect 19636 93050 19660 93052
rect 19716 93050 19740 93052
rect 19796 93050 19820 93052
rect 19658 92998 19660 93050
rect 19722 92998 19734 93050
rect 19796 92998 19798 93050
rect 19636 92996 19660 92998
rect 19716 92996 19740 92998
rect 19796 92996 19820 92998
rect 19580 92976 19876 92996
rect 19580 91964 19876 91984
rect 19636 91962 19660 91964
rect 19716 91962 19740 91964
rect 19796 91962 19820 91964
rect 19658 91910 19660 91962
rect 19722 91910 19734 91962
rect 19796 91910 19798 91962
rect 19636 91908 19660 91910
rect 19716 91908 19740 91910
rect 19796 91908 19820 91910
rect 19580 91888 19876 91908
rect 19580 90876 19876 90896
rect 19636 90874 19660 90876
rect 19716 90874 19740 90876
rect 19796 90874 19820 90876
rect 19658 90822 19660 90874
rect 19722 90822 19734 90874
rect 19796 90822 19798 90874
rect 19636 90820 19660 90822
rect 19716 90820 19740 90822
rect 19796 90820 19820 90822
rect 19580 90800 19876 90820
rect 19580 89788 19876 89808
rect 19636 89786 19660 89788
rect 19716 89786 19740 89788
rect 19796 89786 19820 89788
rect 19658 89734 19660 89786
rect 19722 89734 19734 89786
rect 19796 89734 19798 89786
rect 19636 89732 19660 89734
rect 19716 89732 19740 89734
rect 19796 89732 19820 89734
rect 19580 89712 19876 89732
rect 19064 88800 19116 88806
rect 19064 88742 19116 88748
rect 18788 57520 18840 57526
rect 18788 57462 18840 57468
rect 18696 53032 18748 53038
rect 18696 52974 18748 52980
rect 18972 51060 19024 51066
rect 18972 51002 19024 51008
rect 18788 50380 18840 50386
rect 18788 50322 18840 50328
rect 18604 48816 18656 48822
rect 18604 48758 18656 48764
rect 18420 46640 18472 46646
rect 18420 46582 18472 46588
rect 18144 45348 18196 45354
rect 18144 45290 18196 45296
rect 17972 45070 18184 45098
rect 17960 44940 18012 44946
rect 17960 44882 18012 44888
rect 17972 44810 18000 44882
rect 17960 44804 18012 44810
rect 17960 44746 18012 44752
rect 17684 44328 17736 44334
rect 17684 44270 17736 44276
rect 17696 38010 17724 44270
rect 17684 38004 17736 38010
rect 17684 37946 17736 37952
rect 17500 37936 17552 37942
rect 17500 37878 17552 37884
rect 17696 34066 17724 37946
rect 17868 37936 17920 37942
rect 17868 37878 17920 37884
rect 17880 37806 17908 37878
rect 17868 37800 17920 37806
rect 17868 37742 17920 37748
rect 17972 37466 18000 44746
rect 18156 41546 18184 45070
rect 18236 44940 18288 44946
rect 18236 44882 18288 44888
rect 18248 44742 18276 44882
rect 18236 44736 18288 44742
rect 18236 44678 18288 44684
rect 18144 41540 18196 41546
rect 18144 41482 18196 41488
rect 18236 38956 18288 38962
rect 18236 38898 18288 38904
rect 17960 37460 18012 37466
rect 17960 37402 18012 37408
rect 17776 37324 17828 37330
rect 17776 37266 17828 37272
rect 17684 34060 17736 34066
rect 17684 34002 17736 34008
rect 17696 29306 17724 34002
rect 17684 29300 17736 29306
rect 17684 29242 17736 29248
rect 17696 26314 17724 29242
rect 17684 26308 17736 26314
rect 17684 26250 17736 26256
rect 17788 15978 17816 37266
rect 17868 28416 17920 28422
rect 17868 28358 17920 28364
rect 17880 26994 17908 28358
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17776 15972 17828 15978
rect 17776 15914 17828 15920
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17972 11626 18000 11698
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17696 9926 17724 9998
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 7410 17908 9862
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17972 4842 18000 11562
rect 17972 4814 18092 4842
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 17604 800 17632 2450
rect 17788 800 17816 3878
rect 17972 800 18000 4626
rect 18064 4078 18092 4814
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18248 3670 18276 38898
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 18156 800 18184 3538
rect 18340 800 18368 3878
rect 18432 2582 18460 46582
rect 18616 44878 18644 48758
rect 18696 46504 18748 46510
rect 18696 46446 18748 46452
rect 18708 46102 18736 46446
rect 18696 46096 18748 46102
rect 18696 46038 18748 46044
rect 18800 45914 18828 50322
rect 18984 48686 19012 51002
rect 18972 48680 19024 48686
rect 18972 48622 19024 48628
rect 18708 45886 18828 45914
rect 18604 44872 18656 44878
rect 18604 44814 18656 44820
rect 18512 37664 18564 37670
rect 18512 37606 18564 37612
rect 18524 37398 18552 37606
rect 18512 37392 18564 37398
rect 18512 37334 18564 37340
rect 18604 37324 18656 37330
rect 18604 37266 18656 37272
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 18524 14618 18552 37198
rect 18616 18154 18644 37266
rect 18604 18148 18656 18154
rect 18604 18090 18656 18096
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18616 12434 18644 18090
rect 18708 15094 18736 45886
rect 19076 45554 19104 88742
rect 19580 88700 19876 88720
rect 19636 88698 19660 88700
rect 19716 88698 19740 88700
rect 19796 88698 19820 88700
rect 19658 88646 19660 88698
rect 19722 88646 19734 88698
rect 19796 88646 19798 88698
rect 19636 88644 19660 88646
rect 19716 88644 19740 88646
rect 19796 88644 19820 88646
rect 19580 88624 19876 88644
rect 19580 87612 19876 87632
rect 19636 87610 19660 87612
rect 19716 87610 19740 87612
rect 19796 87610 19820 87612
rect 19658 87558 19660 87610
rect 19722 87558 19734 87610
rect 19796 87558 19798 87610
rect 19636 87556 19660 87558
rect 19716 87556 19740 87558
rect 19796 87556 19820 87558
rect 19580 87536 19876 87556
rect 19580 86524 19876 86544
rect 19636 86522 19660 86524
rect 19716 86522 19740 86524
rect 19796 86522 19820 86524
rect 19658 86470 19660 86522
rect 19722 86470 19734 86522
rect 19796 86470 19798 86522
rect 19636 86468 19660 86470
rect 19716 86468 19740 86470
rect 19796 86468 19820 86470
rect 19580 86448 19876 86468
rect 19580 85436 19876 85456
rect 19636 85434 19660 85436
rect 19716 85434 19740 85436
rect 19796 85434 19820 85436
rect 19658 85382 19660 85434
rect 19722 85382 19734 85434
rect 19796 85382 19798 85434
rect 19636 85380 19660 85382
rect 19716 85380 19740 85382
rect 19796 85380 19820 85382
rect 19580 85360 19876 85380
rect 19580 84348 19876 84368
rect 19636 84346 19660 84348
rect 19716 84346 19740 84348
rect 19796 84346 19820 84348
rect 19658 84294 19660 84346
rect 19722 84294 19734 84346
rect 19796 84294 19798 84346
rect 19636 84292 19660 84294
rect 19716 84292 19740 84294
rect 19796 84292 19820 84294
rect 19580 84272 19876 84292
rect 20364 83570 20392 97106
rect 20456 96558 20484 97294
rect 21192 97170 21220 99200
rect 22112 97306 22140 99200
rect 22100 97300 22152 97306
rect 22100 97242 22152 97248
rect 21456 97232 21508 97238
rect 21456 97174 21508 97180
rect 22836 97232 22888 97238
rect 22836 97174 22888 97180
rect 21180 97164 21232 97170
rect 21180 97106 21232 97112
rect 21364 97096 21416 97102
rect 21364 97038 21416 97044
rect 21376 96762 21404 97038
rect 21364 96756 21416 96762
rect 21364 96698 21416 96704
rect 20444 96552 20496 96558
rect 20444 96494 20496 96500
rect 20444 96416 20496 96422
rect 20444 96358 20496 96364
rect 20352 83564 20404 83570
rect 20352 83506 20404 83512
rect 19580 83260 19876 83280
rect 19636 83258 19660 83260
rect 19716 83258 19740 83260
rect 19796 83258 19820 83260
rect 19658 83206 19660 83258
rect 19722 83206 19734 83258
rect 19796 83206 19798 83258
rect 19636 83204 19660 83206
rect 19716 83204 19740 83206
rect 19796 83204 19820 83206
rect 19580 83184 19876 83204
rect 19580 82172 19876 82192
rect 19636 82170 19660 82172
rect 19716 82170 19740 82172
rect 19796 82170 19820 82172
rect 19658 82118 19660 82170
rect 19722 82118 19734 82170
rect 19796 82118 19798 82170
rect 19636 82116 19660 82118
rect 19716 82116 19740 82118
rect 19796 82116 19820 82118
rect 19580 82096 19876 82116
rect 19580 81084 19876 81104
rect 19636 81082 19660 81084
rect 19716 81082 19740 81084
rect 19796 81082 19820 81084
rect 19658 81030 19660 81082
rect 19722 81030 19734 81082
rect 19796 81030 19798 81082
rect 19636 81028 19660 81030
rect 19716 81028 19740 81030
rect 19796 81028 19820 81030
rect 19580 81008 19876 81028
rect 19580 79996 19876 80016
rect 19636 79994 19660 79996
rect 19716 79994 19740 79996
rect 19796 79994 19820 79996
rect 19658 79942 19660 79994
rect 19722 79942 19734 79994
rect 19796 79942 19798 79994
rect 19636 79940 19660 79942
rect 19716 79940 19740 79942
rect 19796 79940 19820 79942
rect 19580 79920 19876 79940
rect 19580 78908 19876 78928
rect 19636 78906 19660 78908
rect 19716 78906 19740 78908
rect 19796 78906 19820 78908
rect 19658 78854 19660 78906
rect 19722 78854 19734 78906
rect 19796 78854 19798 78906
rect 19636 78852 19660 78854
rect 19716 78852 19740 78854
rect 19796 78852 19820 78854
rect 19580 78832 19876 78852
rect 19580 77820 19876 77840
rect 19636 77818 19660 77820
rect 19716 77818 19740 77820
rect 19796 77818 19820 77820
rect 19658 77766 19660 77818
rect 19722 77766 19734 77818
rect 19796 77766 19798 77818
rect 19636 77764 19660 77766
rect 19716 77764 19740 77766
rect 19796 77764 19820 77766
rect 19580 77744 19876 77764
rect 19580 76732 19876 76752
rect 19636 76730 19660 76732
rect 19716 76730 19740 76732
rect 19796 76730 19820 76732
rect 19658 76678 19660 76730
rect 19722 76678 19734 76730
rect 19796 76678 19798 76730
rect 19636 76676 19660 76678
rect 19716 76676 19740 76678
rect 19796 76676 19820 76678
rect 19580 76656 19876 76676
rect 19580 75644 19876 75664
rect 19636 75642 19660 75644
rect 19716 75642 19740 75644
rect 19796 75642 19820 75644
rect 19658 75590 19660 75642
rect 19722 75590 19734 75642
rect 19796 75590 19798 75642
rect 19636 75588 19660 75590
rect 19716 75588 19740 75590
rect 19796 75588 19820 75590
rect 19580 75568 19876 75588
rect 19580 74556 19876 74576
rect 19636 74554 19660 74556
rect 19716 74554 19740 74556
rect 19796 74554 19820 74556
rect 19658 74502 19660 74554
rect 19722 74502 19734 74554
rect 19796 74502 19798 74554
rect 19636 74500 19660 74502
rect 19716 74500 19740 74502
rect 19796 74500 19820 74502
rect 19580 74480 19876 74500
rect 19580 73468 19876 73488
rect 19636 73466 19660 73468
rect 19716 73466 19740 73468
rect 19796 73466 19820 73468
rect 19658 73414 19660 73466
rect 19722 73414 19734 73466
rect 19796 73414 19798 73466
rect 19636 73412 19660 73414
rect 19716 73412 19740 73414
rect 19796 73412 19820 73414
rect 19580 73392 19876 73412
rect 19580 72380 19876 72400
rect 19636 72378 19660 72380
rect 19716 72378 19740 72380
rect 19796 72378 19820 72380
rect 19658 72326 19660 72378
rect 19722 72326 19734 72378
rect 19796 72326 19798 72378
rect 19636 72324 19660 72326
rect 19716 72324 19740 72326
rect 19796 72324 19820 72326
rect 19580 72304 19876 72324
rect 19580 71292 19876 71312
rect 19636 71290 19660 71292
rect 19716 71290 19740 71292
rect 19796 71290 19820 71292
rect 19658 71238 19660 71290
rect 19722 71238 19734 71290
rect 19796 71238 19798 71290
rect 19636 71236 19660 71238
rect 19716 71236 19740 71238
rect 19796 71236 19820 71238
rect 19580 71216 19876 71236
rect 19580 70204 19876 70224
rect 19636 70202 19660 70204
rect 19716 70202 19740 70204
rect 19796 70202 19820 70204
rect 19658 70150 19660 70202
rect 19722 70150 19734 70202
rect 19796 70150 19798 70202
rect 19636 70148 19660 70150
rect 19716 70148 19740 70150
rect 19796 70148 19820 70150
rect 19580 70128 19876 70148
rect 19580 69116 19876 69136
rect 19636 69114 19660 69116
rect 19716 69114 19740 69116
rect 19796 69114 19820 69116
rect 19658 69062 19660 69114
rect 19722 69062 19734 69114
rect 19796 69062 19798 69114
rect 19636 69060 19660 69062
rect 19716 69060 19740 69062
rect 19796 69060 19820 69062
rect 19580 69040 19876 69060
rect 19580 68028 19876 68048
rect 19636 68026 19660 68028
rect 19716 68026 19740 68028
rect 19796 68026 19820 68028
rect 19658 67974 19660 68026
rect 19722 67974 19734 68026
rect 19796 67974 19798 68026
rect 19636 67972 19660 67974
rect 19716 67972 19740 67974
rect 19796 67972 19820 67974
rect 19580 67952 19876 67972
rect 19432 67244 19484 67250
rect 19432 67186 19484 67192
rect 19340 63436 19392 63442
rect 19340 63378 19392 63384
rect 19352 58682 19380 63378
rect 19340 58676 19392 58682
rect 19340 58618 19392 58624
rect 19248 49156 19300 49162
rect 19248 49098 19300 49104
rect 19260 48686 19288 49098
rect 19248 48680 19300 48686
rect 19248 48622 19300 48628
rect 19248 46572 19300 46578
rect 19248 46514 19300 46520
rect 18800 45526 19104 45554
rect 18800 41478 18828 45526
rect 19260 44946 19288 46514
rect 19248 44940 19300 44946
rect 19248 44882 19300 44888
rect 18788 41472 18840 41478
rect 18788 41414 18840 41420
rect 18800 24886 18828 41414
rect 18972 39976 19024 39982
rect 18972 39918 19024 39924
rect 18984 38962 19012 39918
rect 18972 38956 19024 38962
rect 18972 38898 19024 38904
rect 18788 24880 18840 24886
rect 18788 24822 18840 24828
rect 19156 24744 19208 24750
rect 19156 24686 19208 24692
rect 19168 22574 19196 24686
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 18696 15088 18748 15094
rect 18696 15030 18748 15036
rect 19076 12782 19104 19926
rect 19352 18222 19380 58618
rect 19444 36650 19472 67186
rect 20456 67182 20484 96358
rect 21088 83632 21140 83638
rect 21088 83574 21140 83580
rect 20720 78804 20772 78810
rect 20720 78746 20772 78752
rect 20732 77654 20760 78746
rect 20720 77648 20772 77654
rect 20720 77590 20772 77596
rect 20732 77110 20760 77590
rect 20720 77104 20772 77110
rect 20720 77046 20772 77052
rect 20628 67244 20680 67250
rect 20628 67186 20680 67192
rect 20260 67176 20312 67182
rect 20260 67118 20312 67124
rect 20444 67176 20496 67182
rect 20444 67118 20496 67124
rect 20076 67040 20128 67046
rect 20076 66982 20128 66988
rect 19580 66940 19876 66960
rect 19636 66938 19660 66940
rect 19716 66938 19740 66940
rect 19796 66938 19820 66940
rect 19658 66886 19660 66938
rect 19722 66886 19734 66938
rect 19796 66886 19798 66938
rect 19636 66884 19660 66886
rect 19716 66884 19740 66886
rect 19796 66884 19820 66886
rect 19580 66864 19876 66884
rect 19580 65852 19876 65872
rect 19636 65850 19660 65852
rect 19716 65850 19740 65852
rect 19796 65850 19820 65852
rect 19658 65798 19660 65850
rect 19722 65798 19734 65850
rect 19796 65798 19798 65850
rect 19636 65796 19660 65798
rect 19716 65796 19740 65798
rect 19796 65796 19820 65798
rect 19580 65776 19876 65796
rect 19580 64764 19876 64784
rect 19636 64762 19660 64764
rect 19716 64762 19740 64764
rect 19796 64762 19820 64764
rect 19658 64710 19660 64762
rect 19722 64710 19734 64762
rect 19796 64710 19798 64762
rect 19636 64708 19660 64710
rect 19716 64708 19740 64710
rect 19796 64708 19820 64710
rect 19580 64688 19876 64708
rect 19580 63676 19876 63696
rect 19636 63674 19660 63676
rect 19716 63674 19740 63676
rect 19796 63674 19820 63676
rect 19658 63622 19660 63674
rect 19722 63622 19734 63674
rect 19796 63622 19798 63674
rect 19636 63620 19660 63622
rect 19716 63620 19740 63622
rect 19796 63620 19820 63622
rect 19580 63600 19876 63620
rect 19580 62588 19876 62608
rect 19636 62586 19660 62588
rect 19716 62586 19740 62588
rect 19796 62586 19820 62588
rect 19658 62534 19660 62586
rect 19722 62534 19734 62586
rect 19796 62534 19798 62586
rect 19636 62532 19660 62534
rect 19716 62532 19740 62534
rect 19796 62532 19820 62534
rect 19580 62512 19876 62532
rect 19580 61500 19876 61520
rect 19636 61498 19660 61500
rect 19716 61498 19740 61500
rect 19796 61498 19820 61500
rect 19658 61446 19660 61498
rect 19722 61446 19734 61498
rect 19796 61446 19798 61498
rect 19636 61444 19660 61446
rect 19716 61444 19740 61446
rect 19796 61444 19820 61446
rect 19580 61424 19876 61444
rect 19580 60412 19876 60432
rect 19636 60410 19660 60412
rect 19716 60410 19740 60412
rect 19796 60410 19820 60412
rect 19658 60358 19660 60410
rect 19722 60358 19734 60410
rect 19796 60358 19798 60410
rect 19636 60356 19660 60358
rect 19716 60356 19740 60358
rect 19796 60356 19820 60358
rect 19580 60336 19876 60356
rect 19580 59324 19876 59344
rect 19636 59322 19660 59324
rect 19716 59322 19740 59324
rect 19796 59322 19820 59324
rect 19658 59270 19660 59322
rect 19722 59270 19734 59322
rect 19796 59270 19798 59322
rect 19636 59268 19660 59270
rect 19716 59268 19740 59270
rect 19796 59268 19820 59270
rect 19580 59248 19876 59268
rect 19580 58236 19876 58256
rect 19636 58234 19660 58236
rect 19716 58234 19740 58236
rect 19796 58234 19820 58236
rect 19658 58182 19660 58234
rect 19722 58182 19734 58234
rect 19796 58182 19798 58234
rect 19636 58180 19660 58182
rect 19716 58180 19740 58182
rect 19796 58180 19820 58182
rect 19580 58160 19876 58180
rect 19580 57148 19876 57168
rect 19636 57146 19660 57148
rect 19716 57146 19740 57148
rect 19796 57146 19820 57148
rect 19658 57094 19660 57146
rect 19722 57094 19734 57146
rect 19796 57094 19798 57146
rect 19636 57092 19660 57094
rect 19716 57092 19740 57094
rect 19796 57092 19820 57094
rect 19580 57072 19876 57092
rect 19580 56060 19876 56080
rect 19636 56058 19660 56060
rect 19716 56058 19740 56060
rect 19796 56058 19820 56060
rect 19658 56006 19660 56058
rect 19722 56006 19734 56058
rect 19796 56006 19798 56058
rect 19636 56004 19660 56006
rect 19716 56004 19740 56006
rect 19796 56004 19820 56006
rect 19580 55984 19876 56004
rect 19580 54972 19876 54992
rect 19636 54970 19660 54972
rect 19716 54970 19740 54972
rect 19796 54970 19820 54972
rect 19658 54918 19660 54970
rect 19722 54918 19734 54970
rect 19796 54918 19798 54970
rect 19636 54916 19660 54918
rect 19716 54916 19740 54918
rect 19796 54916 19820 54918
rect 19580 54896 19876 54916
rect 19580 53884 19876 53904
rect 19636 53882 19660 53884
rect 19716 53882 19740 53884
rect 19796 53882 19820 53884
rect 19658 53830 19660 53882
rect 19722 53830 19734 53882
rect 19796 53830 19798 53882
rect 19636 53828 19660 53830
rect 19716 53828 19740 53830
rect 19796 53828 19820 53830
rect 19580 53808 19876 53828
rect 19892 52964 19944 52970
rect 19892 52906 19944 52912
rect 19580 52796 19876 52816
rect 19636 52794 19660 52796
rect 19716 52794 19740 52796
rect 19796 52794 19820 52796
rect 19658 52742 19660 52794
rect 19722 52742 19734 52794
rect 19796 52742 19798 52794
rect 19636 52740 19660 52742
rect 19716 52740 19740 52742
rect 19796 52740 19820 52742
rect 19580 52720 19876 52740
rect 19580 51708 19876 51728
rect 19636 51706 19660 51708
rect 19716 51706 19740 51708
rect 19796 51706 19820 51708
rect 19658 51654 19660 51706
rect 19722 51654 19734 51706
rect 19796 51654 19798 51706
rect 19636 51652 19660 51654
rect 19716 51652 19740 51654
rect 19796 51652 19820 51654
rect 19580 51632 19876 51652
rect 19580 50620 19876 50640
rect 19636 50618 19660 50620
rect 19716 50618 19740 50620
rect 19796 50618 19820 50620
rect 19658 50566 19660 50618
rect 19722 50566 19734 50618
rect 19796 50566 19798 50618
rect 19636 50564 19660 50566
rect 19716 50564 19740 50566
rect 19796 50564 19820 50566
rect 19580 50544 19876 50564
rect 19904 50386 19932 52906
rect 19892 50380 19944 50386
rect 19892 50322 19944 50328
rect 19524 50244 19576 50250
rect 19524 50186 19576 50192
rect 19536 49774 19564 50186
rect 19524 49768 19576 49774
rect 19524 49710 19576 49716
rect 19580 49532 19876 49552
rect 19636 49530 19660 49532
rect 19716 49530 19740 49532
rect 19796 49530 19820 49532
rect 19658 49478 19660 49530
rect 19722 49478 19734 49530
rect 19796 49478 19798 49530
rect 19636 49476 19660 49478
rect 19716 49476 19740 49478
rect 19796 49476 19820 49478
rect 19580 49456 19876 49476
rect 19580 48444 19876 48464
rect 19636 48442 19660 48444
rect 19716 48442 19740 48444
rect 19796 48442 19820 48444
rect 19658 48390 19660 48442
rect 19722 48390 19734 48442
rect 19796 48390 19798 48442
rect 19636 48388 19660 48390
rect 19716 48388 19740 48390
rect 19796 48388 19820 48390
rect 19580 48368 19876 48388
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 20088 45554 20116 66982
rect 20272 45554 20300 67118
rect 20456 62898 20484 67118
rect 20640 62966 20668 67186
rect 20628 62960 20680 62966
rect 20628 62902 20680 62908
rect 20444 62892 20496 62898
rect 20444 62834 20496 62840
rect 20996 59084 21048 59090
rect 20996 59026 21048 59032
rect 20536 48544 20588 48550
rect 20536 48486 20588 48492
rect 19996 45526 20116 45554
rect 20180 45526 20300 45554
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 19996 40730 20024 45526
rect 20180 40746 20208 45526
rect 19984 40724 20036 40730
rect 19984 40666 20036 40672
rect 20088 40718 20208 40746
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 19892 37800 19944 37806
rect 19892 37742 19944 37748
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19432 36644 19484 36650
rect 19432 36586 19484 36592
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19904 34542 19932 37742
rect 19996 37330 20024 40666
rect 19984 37324 20036 37330
rect 19984 37266 20036 37272
rect 19892 34536 19944 34542
rect 19892 34478 19944 34484
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 20088 30394 20116 40718
rect 20168 38344 20220 38350
rect 20168 38286 20220 38292
rect 20076 30388 20128 30394
rect 20076 30330 20128 30336
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19432 26308 19484 26314
rect 19432 26250 19484 26256
rect 19444 24750 19472 26250
rect 20088 26234 20116 30330
rect 19996 26206 20116 26234
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19432 24744 19484 24750
rect 19432 24686 19484 24692
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19444 22234 19472 22510
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19444 18290 19472 20334
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19076 12434 19104 12718
rect 18524 12406 18644 12434
rect 18984 12406 19104 12434
rect 18524 4554 18552 12406
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18512 4548 18564 4554
rect 18512 4490 18564 4496
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18616 800 18644 5102
rect 18892 4078 18920 8026
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 18984 3194 19012 12406
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18800 800 18828 2926
rect 19076 2774 19104 3878
rect 18984 2746 19104 2774
rect 18984 800 19012 2746
rect 19168 2582 19196 10950
rect 19260 3058 19288 15982
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 19156 2576 19208 2582
rect 19156 2518 19208 2524
rect 19260 2394 19288 2858
rect 19168 2366 19288 2394
rect 19168 800 19196 2366
rect 19352 800 19380 2926
rect 19444 2922 19472 4626
rect 19904 4078 19932 18226
rect 19996 13462 20024 26206
rect 20076 24744 20128 24750
rect 20076 24686 20128 24692
rect 20088 24070 20116 24686
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 19984 13456 20036 13462
rect 19984 13398 20036 13404
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19984 3936 20036 3942
rect 19904 3896 19984 3924
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19904 1986 19932 3896
rect 19984 3878 20036 3884
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19628 1958 19932 1986
rect 19628 800 19656 1958
rect 19800 1896 19852 1902
rect 19800 1838 19852 1844
rect 19812 800 19840 1838
rect 19996 800 20024 3538
rect 20088 1902 20116 4014
rect 20180 3670 20208 38286
rect 20548 26926 20576 48486
rect 21008 37466 21036 59026
rect 21100 53446 21128 83574
rect 21364 76900 21416 76906
rect 21364 76842 21416 76848
rect 21272 76832 21324 76838
rect 21272 76774 21324 76780
rect 21180 53644 21232 53650
rect 21180 53586 21232 53592
rect 21088 53440 21140 53446
rect 21088 53382 21140 53388
rect 20720 37460 20772 37466
rect 20720 37402 20772 37408
rect 20996 37460 21048 37466
rect 20996 37402 21048 37408
rect 20628 36644 20680 36650
rect 20628 36586 20680 36592
rect 20640 36378 20668 36586
rect 20628 36372 20680 36378
rect 20628 36314 20680 36320
rect 20732 36174 20760 37402
rect 20720 36168 20772 36174
rect 20720 36110 20772 36116
rect 20536 26920 20588 26926
rect 20536 26862 20588 26868
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 21100 26382 21128 26862
rect 21088 26376 21140 26382
rect 21088 26318 21140 26324
rect 21100 26042 21128 26318
rect 21088 26036 21140 26042
rect 21088 25978 21140 25984
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 18698 20760 20742
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20168 3664 20220 3670
rect 20168 3606 20220 3612
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20076 1896 20128 1902
rect 20076 1838 20128 1844
rect 20180 800 20208 3334
rect 20272 3058 20300 16594
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20640 10266 20668 11766
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20352 4684 20404 4690
rect 20352 4626 20404 4632
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20364 800 20392 4626
rect 20548 2582 20576 9386
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 4010 20668 8230
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20732 4622 20760 6054
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20628 4004 20680 4010
rect 20628 3946 20680 3952
rect 21008 3670 21036 19246
rect 21192 16998 21220 53586
rect 21284 29782 21312 76774
rect 21376 76498 21404 76842
rect 21364 76492 21416 76498
rect 21364 76434 21416 76440
rect 21468 65618 21496 97174
rect 22100 87780 22152 87786
rect 22100 87722 22152 87728
rect 22112 87446 22140 87722
rect 22100 87440 22152 87446
rect 22100 87382 22152 87388
rect 21456 65612 21508 65618
rect 21456 65554 21508 65560
rect 21468 64874 21496 65554
rect 21468 64846 21772 64874
rect 21548 53644 21600 53650
rect 21548 53586 21600 53592
rect 21364 53576 21416 53582
rect 21364 53518 21416 53524
rect 21376 53446 21404 53518
rect 21364 53440 21416 53446
rect 21364 53382 21416 53388
rect 21376 52018 21404 53382
rect 21364 52012 21416 52018
rect 21364 51954 21416 51960
rect 21364 45280 21416 45286
rect 21364 45222 21416 45228
rect 21376 45014 21404 45222
rect 21364 45008 21416 45014
rect 21364 44950 21416 44956
rect 21560 42702 21588 53586
rect 21640 53440 21692 53446
rect 21640 53382 21692 53388
rect 21652 51814 21680 53382
rect 21640 51808 21692 51814
rect 21640 51750 21692 51756
rect 21548 42696 21600 42702
rect 21548 42638 21600 42644
rect 21560 42090 21588 42638
rect 21548 42084 21600 42090
rect 21548 42026 21600 42032
rect 21744 34134 21772 64846
rect 22100 63028 22152 63034
rect 22100 62970 22152 62976
rect 21824 47592 21876 47598
rect 21824 47534 21876 47540
rect 21732 34128 21784 34134
rect 21732 34070 21784 34076
rect 21364 30728 21416 30734
rect 21364 30670 21416 30676
rect 21272 29776 21324 29782
rect 21272 29718 21324 29724
rect 21376 28422 21404 30670
rect 21364 28416 21416 28422
rect 21364 28358 21416 28364
rect 21376 26858 21404 28358
rect 21732 27532 21784 27538
rect 21732 27474 21784 27480
rect 21364 26852 21416 26858
rect 21364 26794 21416 26800
rect 21744 26586 21772 27474
rect 21732 26580 21784 26586
rect 21732 26522 21784 26528
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21284 24342 21312 24550
rect 21272 24336 21324 24342
rect 21272 24278 21324 24284
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 20996 3664 21048 3670
rect 20996 3606 21048 3612
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20536 2576 20588 2582
rect 20536 2518 20588 2524
rect 20640 800 20668 2994
rect 20824 800 20852 3402
rect 21100 2394 21128 4626
rect 21376 3534 21404 16934
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21468 3058 21496 7958
rect 21744 6118 21772 26522
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21640 2916 21692 2922
rect 21640 2858 21692 2864
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21008 2366 21128 2394
rect 21008 800 21036 2366
rect 21192 800 21220 2450
rect 21376 800 21404 2790
rect 21652 800 21680 2858
rect 21836 2582 21864 47534
rect 21916 29708 21968 29714
rect 21916 29650 21968 29656
rect 21928 20806 21956 29650
rect 22112 22506 22140 62970
rect 22744 57452 22796 57458
rect 22744 57394 22796 57400
rect 22468 50992 22520 50998
rect 22468 50934 22520 50940
rect 22480 50318 22508 50934
rect 22468 50312 22520 50318
rect 22468 50254 22520 50260
rect 22652 50244 22704 50250
rect 22652 50186 22704 50192
rect 22284 50176 22336 50182
rect 22284 50118 22336 50124
rect 22296 30734 22324 50118
rect 22664 49774 22692 50186
rect 22652 49768 22704 49774
rect 22652 49710 22704 49716
rect 22376 49632 22428 49638
rect 22376 49574 22428 49580
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 22284 29504 22336 29510
rect 22284 29446 22336 29452
rect 22204 29238 22232 29446
rect 22192 29232 22244 29238
rect 22192 29174 22244 29180
rect 22296 29102 22324 29446
rect 22284 29096 22336 29102
rect 22284 29038 22336 29044
rect 22100 22500 22152 22506
rect 22100 22442 22152 22448
rect 22388 21622 22416 49574
rect 22652 49088 22704 49094
rect 22652 49030 22704 49036
rect 22664 48822 22692 49030
rect 22652 48816 22704 48822
rect 22652 48758 22704 48764
rect 22652 26036 22704 26042
rect 22652 25978 22704 25984
rect 22376 21616 22428 21622
rect 22376 21558 22428 21564
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 21928 3670 21956 20538
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 22112 8022 22140 14282
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 21916 3664 21968 3670
rect 21916 3606 21968 3612
rect 21824 2576 21876 2582
rect 21824 2518 21876 2524
rect 21824 2372 21876 2378
rect 21824 2314 21876 2320
rect 21836 800 21864 2314
rect 22020 800 22048 4014
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22204 800 22232 3538
rect 22664 2990 22692 25978
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 22756 2650 22784 57394
rect 22848 48618 22876 97174
rect 22940 96626 22968 99200
rect 23112 97164 23164 97170
rect 23112 97106 23164 97112
rect 22928 96620 22980 96626
rect 22928 96562 22980 96568
rect 23020 96484 23072 96490
rect 23020 96426 23072 96432
rect 23032 53174 23060 96426
rect 23124 61402 23152 97106
rect 23572 96960 23624 96966
rect 23572 96902 23624 96908
rect 23584 96558 23612 96902
rect 23860 96558 23888 99200
rect 23940 97572 23992 97578
rect 23940 97514 23992 97520
rect 23952 97238 23980 97514
rect 24688 97238 24716 99200
rect 23940 97232 23992 97238
rect 23940 97174 23992 97180
rect 24676 97232 24728 97238
rect 24676 97174 24728 97180
rect 24492 97164 24544 97170
rect 24492 97106 24544 97112
rect 24504 96966 24532 97106
rect 24492 96960 24544 96966
rect 24492 96902 24544 96908
rect 23572 96552 23624 96558
rect 23572 96494 23624 96500
rect 23848 96552 23900 96558
rect 23848 96494 23900 96500
rect 24032 96416 24084 96422
rect 24032 96358 24084 96364
rect 23480 92132 23532 92138
rect 23480 92074 23532 92080
rect 23664 92132 23716 92138
rect 23664 92074 23716 92080
rect 23388 87780 23440 87786
rect 23388 87722 23440 87728
rect 23400 80054 23428 87722
rect 23216 80026 23428 80054
rect 23216 72010 23244 80026
rect 23388 77512 23440 77518
rect 23388 77454 23440 77460
rect 23400 77178 23428 77454
rect 23388 77172 23440 77178
rect 23388 77114 23440 77120
rect 23204 72004 23256 72010
rect 23204 71946 23256 71952
rect 23112 61396 23164 61402
rect 23112 61338 23164 61344
rect 23020 53168 23072 53174
rect 23020 53110 23072 53116
rect 23112 51808 23164 51814
rect 23112 51750 23164 51756
rect 22928 49972 22980 49978
rect 22928 49914 22980 49920
rect 23020 49972 23072 49978
rect 23020 49914 23072 49920
rect 22940 49774 22968 49914
rect 23032 49774 23060 49914
rect 22928 49768 22980 49774
rect 22928 49710 22980 49716
rect 23020 49768 23072 49774
rect 23020 49710 23072 49716
rect 23032 49638 23060 49710
rect 23020 49632 23072 49638
rect 23020 49574 23072 49580
rect 22836 48612 22888 48618
rect 22836 48554 22888 48560
rect 23124 45554 23152 51750
rect 22940 45526 23152 45554
rect 22836 21616 22888 21622
rect 22836 21558 22888 21564
rect 22848 8090 22876 21558
rect 22940 8294 22968 45526
rect 23216 28694 23244 71946
rect 23492 67590 23520 92074
rect 23676 85610 23704 92074
rect 23664 85604 23716 85610
rect 23664 85546 23716 85552
rect 23676 85270 23704 85546
rect 23664 85264 23716 85270
rect 23664 85206 23716 85212
rect 24044 78674 24072 96358
rect 24216 86692 24268 86698
rect 24216 86634 24268 86640
rect 24032 78668 24084 78674
rect 24032 78610 24084 78616
rect 23664 78056 23716 78062
rect 23664 77998 23716 78004
rect 23676 69766 23704 77998
rect 24124 76356 24176 76362
rect 24124 76298 24176 76304
rect 24032 71392 24084 71398
rect 24032 71334 24084 71340
rect 24044 71126 24072 71334
rect 24032 71120 24084 71126
rect 24032 71062 24084 71068
rect 23664 69760 23716 69766
rect 23664 69702 23716 69708
rect 23480 67584 23532 67590
rect 23480 67526 23532 67532
rect 23756 67584 23808 67590
rect 23756 67526 23808 67532
rect 23768 66706 23796 67526
rect 23756 66700 23808 66706
rect 23756 66642 23808 66648
rect 24136 63850 24164 76298
rect 24228 73778 24256 86634
rect 24400 85604 24452 85610
rect 24400 85546 24452 85552
rect 24216 73772 24268 73778
rect 24216 73714 24268 73720
rect 24124 63844 24176 63850
rect 24124 63786 24176 63792
rect 23940 53712 23992 53718
rect 23940 53654 23992 53660
rect 23296 50720 23348 50726
rect 23296 50662 23348 50668
rect 23308 49774 23336 50662
rect 23848 50176 23900 50182
rect 23848 50118 23900 50124
rect 23860 49774 23888 50118
rect 23296 49768 23348 49774
rect 23296 49710 23348 49716
rect 23848 49768 23900 49774
rect 23848 49710 23900 49716
rect 23308 45286 23336 49710
rect 23952 48618 23980 53654
rect 24032 49904 24084 49910
rect 24032 49846 24084 49852
rect 24044 49434 24072 49846
rect 24032 49428 24084 49434
rect 24032 49370 24084 49376
rect 24136 48770 24164 63786
rect 24228 53718 24256 73714
rect 24216 53712 24268 53718
rect 24216 53654 24268 53660
rect 24216 51944 24268 51950
rect 24216 51886 24268 51892
rect 24044 48742 24164 48770
rect 24228 48770 24256 51886
rect 24308 49088 24360 49094
rect 24308 49030 24360 49036
rect 24320 48890 24348 49030
rect 24308 48884 24360 48890
rect 24308 48826 24360 48832
rect 24228 48742 24348 48770
rect 23940 48612 23992 48618
rect 23940 48554 23992 48560
rect 24044 45642 24072 48742
rect 24216 48612 24268 48618
rect 24216 48554 24268 48560
rect 24044 45614 24164 45642
rect 23296 45280 23348 45286
rect 23296 45222 23348 45228
rect 23572 44328 23624 44334
rect 23572 44270 23624 44276
rect 23584 36106 23612 44270
rect 23572 36100 23624 36106
rect 23572 36042 23624 36048
rect 23940 35556 23992 35562
rect 23940 35498 23992 35504
rect 23204 28688 23256 28694
rect 23204 28630 23256 28636
rect 23020 26852 23072 26858
rect 23020 26794 23072 26800
rect 23032 14550 23060 26794
rect 23112 22500 23164 22506
rect 23112 22442 23164 22448
rect 23020 14544 23072 14550
rect 23020 14486 23072 14492
rect 23124 12782 23152 22442
rect 23952 20398 23980 35498
rect 24136 32502 24164 45614
rect 24228 39302 24256 48554
rect 24216 39296 24268 39302
rect 24216 39238 24268 39244
rect 24124 32496 24176 32502
rect 24124 32438 24176 32444
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 24136 19310 24164 32438
rect 24216 31136 24268 31142
rect 24216 31078 24268 31084
rect 24228 20602 24256 31078
rect 24216 20596 24268 20602
rect 24216 20538 24268 20544
rect 24320 20466 24348 48742
rect 24412 38214 24440 85546
rect 24504 76634 24532 96902
rect 25608 96626 25636 99200
rect 26436 97238 26464 99200
rect 27356 97306 27384 99200
rect 27344 97300 27396 97306
rect 27344 97242 27396 97248
rect 26424 97232 26476 97238
rect 26424 97174 26476 97180
rect 26056 97164 26108 97170
rect 26056 97106 26108 97112
rect 25596 96620 25648 96626
rect 25596 96562 25648 96568
rect 25688 96484 25740 96490
rect 25688 96426 25740 96432
rect 25504 94240 25556 94246
rect 25504 94182 25556 94188
rect 24492 76628 24544 76634
rect 24492 76570 24544 76576
rect 25044 74112 25096 74118
rect 25044 74054 25096 74060
rect 25056 73914 25084 74054
rect 25044 73908 25096 73914
rect 25044 73850 25096 73856
rect 25320 71936 25372 71942
rect 25320 71878 25372 71884
rect 24492 50380 24544 50386
rect 24492 50322 24544 50328
rect 24504 43790 24532 50322
rect 24860 44192 24912 44198
rect 24860 44134 24912 44140
rect 24584 43852 24636 43858
rect 24584 43794 24636 43800
rect 24492 43784 24544 43790
rect 24492 43726 24544 43732
rect 24400 38208 24452 38214
rect 24400 38150 24452 38156
rect 24308 20460 24360 20466
rect 24308 20402 24360 20408
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24228 19990 24256 20334
rect 24320 20058 24348 20402
rect 24492 20392 24544 20398
rect 24492 20334 24544 20340
rect 24504 20262 24532 20334
rect 24492 20256 24544 20262
rect 24492 20198 24544 20204
rect 24308 20052 24360 20058
rect 24308 19994 24360 20000
rect 24216 19984 24268 19990
rect 24216 19926 24268 19932
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 24308 16720 24360 16726
rect 24308 16662 24360 16668
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23216 9518 23244 13806
rect 24320 10606 24348 16662
rect 24032 10600 24084 10606
rect 24032 10542 24084 10548
rect 24308 10600 24360 10606
rect 24308 10542 24360 10548
rect 24044 9926 24072 10542
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24400 9920 24452 9926
rect 24400 9862 24452 9868
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 22836 4072 22888 4078
rect 23296 4072 23348 4078
rect 22836 4014 22888 4020
rect 23216 4032 23296 4060
rect 22744 2644 22796 2650
rect 22744 2586 22796 2592
rect 22468 2304 22520 2310
rect 22468 2246 22520 2252
rect 22480 800 22508 2246
rect 22848 2122 22876 4014
rect 22928 2916 22980 2922
rect 22928 2858 22980 2864
rect 22664 2094 22876 2122
rect 22664 800 22692 2094
rect 22940 1578 22968 2858
rect 23020 2372 23072 2378
rect 23020 2314 23072 2320
rect 22848 1550 22968 1578
rect 22848 800 22876 1550
rect 23032 800 23060 2314
rect 23216 800 23244 4032
rect 23296 4014 23348 4020
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 23492 800 23520 3538
rect 23860 2582 23888 8230
rect 24412 5166 24440 9862
rect 24492 7812 24544 7818
rect 24492 7754 24544 7760
rect 24400 5160 24452 5166
rect 24400 5102 24452 5108
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23848 2576 23900 2582
rect 23848 2518 23900 2524
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 23676 800 23704 2382
rect 23952 2122 23980 4014
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 23860 2094 23980 2122
rect 23860 800 23888 2094
rect 24044 800 24072 2926
rect 24504 2582 24532 7754
rect 24596 5030 24624 43794
rect 24872 41274 24900 44134
rect 24860 41268 24912 41274
rect 24860 41210 24912 41216
rect 24872 40934 24900 41210
rect 24860 40928 24912 40934
rect 24860 40870 24912 40876
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24872 19990 24900 20334
rect 24860 19984 24912 19990
rect 24860 19926 24912 19932
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 24780 16726 24808 17546
rect 24768 16720 24820 16726
rect 24768 16662 24820 16668
rect 24584 5024 24636 5030
rect 24584 4966 24636 4972
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 24584 4072 24636 4078
rect 24584 4014 24636 4020
rect 24492 2576 24544 2582
rect 24492 2518 24544 2524
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 24228 800 24256 2450
rect 24596 2122 24624 4014
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24504 2094 24624 2122
rect 24504 800 24532 2094
rect 24688 800 24716 3538
rect 24860 2372 24912 2378
rect 24860 2314 24912 2320
rect 24872 800 24900 2314
rect 25056 800 25084 4626
rect 25228 3460 25280 3466
rect 25228 3402 25280 3408
rect 25240 800 25268 3402
rect 25332 3194 25360 71878
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 25424 8974 25452 27406
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25516 8294 25544 94182
rect 25700 80054 25728 96426
rect 25872 94376 25924 94382
rect 25872 94318 25924 94324
rect 25700 80026 25820 80054
rect 25792 78810 25820 80026
rect 25780 78804 25832 78810
rect 25780 78746 25832 78752
rect 25688 70848 25740 70854
rect 25688 70790 25740 70796
rect 25700 70650 25728 70790
rect 25688 70644 25740 70650
rect 25688 70586 25740 70592
rect 25792 70394 25820 78746
rect 25884 75206 25912 94318
rect 25964 77580 26016 77586
rect 25964 77522 26016 77528
rect 25872 75200 25924 75206
rect 25872 75142 25924 75148
rect 25700 70366 25820 70394
rect 25596 54120 25648 54126
rect 25596 54062 25648 54068
rect 25608 41206 25636 54062
rect 25700 53514 25728 70366
rect 25976 65550 26004 77522
rect 26068 73846 26096 97106
rect 28184 97102 28212 99200
rect 29012 97238 29040 99200
rect 29932 97306 29960 99200
rect 30760 97306 30788 99200
rect 31680 97866 31708 99200
rect 31680 97838 31800 97866
rect 29920 97300 29972 97306
rect 29920 97242 29972 97248
rect 30748 97300 30800 97306
rect 30748 97242 30800 97248
rect 31772 97238 31800 97838
rect 32508 97306 32536 99200
rect 32496 97300 32548 97306
rect 32496 97242 32548 97248
rect 29000 97232 29052 97238
rect 29000 97174 29052 97180
rect 31760 97232 31812 97238
rect 31760 97174 31812 97180
rect 28264 97164 28316 97170
rect 28264 97106 28316 97112
rect 29828 97164 29880 97170
rect 29828 97106 29880 97112
rect 31024 97164 31076 97170
rect 31024 97106 31076 97112
rect 32496 97164 32548 97170
rect 32496 97106 32548 97112
rect 28172 97096 28224 97102
rect 28172 97038 28224 97044
rect 26608 96960 26660 96966
rect 26608 96902 26660 96908
rect 26620 83026 26648 96902
rect 26884 96008 26936 96014
rect 26884 95950 26936 95956
rect 26608 83020 26660 83026
rect 26608 82962 26660 82968
rect 26148 77580 26200 77586
rect 26148 77522 26200 77528
rect 26516 77580 26568 77586
rect 26516 77522 26568 77528
rect 26056 73840 26108 73846
rect 26056 73782 26108 73788
rect 25964 65544 26016 65550
rect 25964 65486 26016 65492
rect 25688 53508 25740 53514
rect 25688 53450 25740 53456
rect 25700 46714 25728 53450
rect 25872 49156 25924 49162
rect 25872 49098 25924 49104
rect 25688 46708 25740 46714
rect 25688 46650 25740 46656
rect 25596 41200 25648 41206
rect 25596 41142 25648 41148
rect 25688 34536 25740 34542
rect 25688 34478 25740 34484
rect 25700 29186 25728 34478
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 25792 29306 25820 30194
rect 25780 29300 25832 29306
rect 25780 29242 25832 29248
rect 25700 29158 25820 29186
rect 25686 29064 25742 29073
rect 25686 28999 25688 29008
rect 25740 28999 25742 29008
rect 25688 28970 25740 28976
rect 25504 8288 25556 8294
rect 25504 8230 25556 8236
rect 25688 4684 25740 4690
rect 25688 4626 25740 4632
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 25332 2990 25360 3130
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 25516 800 25544 2858
rect 25700 800 25728 4626
rect 25792 2582 25820 29158
rect 25884 19990 25912 49098
rect 26056 30184 26108 30190
rect 26056 30126 26108 30132
rect 26068 29102 26096 30126
rect 26160 29782 26188 77522
rect 26424 77376 26476 77382
rect 26528 77330 26556 77522
rect 26476 77324 26556 77330
rect 26424 77318 26556 77324
rect 26608 77376 26660 77382
rect 26608 77318 26660 77324
rect 26436 77302 26556 77318
rect 26424 71188 26476 71194
rect 26424 71130 26476 71136
rect 26436 71097 26464 71130
rect 26422 71088 26478 71097
rect 26332 71052 26384 71058
rect 26422 71023 26478 71032
rect 26332 70994 26384 71000
rect 26344 56234 26372 70994
rect 26424 64320 26476 64326
rect 26424 64262 26476 64268
rect 26332 56228 26384 56234
rect 26332 56170 26384 56176
rect 26436 51074 26464 64262
rect 26528 56166 26556 77302
rect 26620 56234 26648 77318
rect 26792 74112 26844 74118
rect 26792 74054 26844 74060
rect 26804 71126 26832 74054
rect 26792 71120 26844 71126
rect 26698 71088 26754 71097
rect 26792 71062 26844 71068
rect 26698 71023 26700 71032
rect 26752 71023 26754 71032
rect 26700 70994 26752 71000
rect 26792 70984 26844 70990
rect 26792 70926 26844 70932
rect 26804 69358 26832 70926
rect 26792 69352 26844 69358
rect 26792 69294 26844 69300
rect 26896 68270 26924 95950
rect 27068 91656 27120 91662
rect 27068 91598 27120 91604
rect 26976 71392 27028 71398
rect 26976 71334 27028 71340
rect 26988 71194 27016 71334
rect 26976 71188 27028 71194
rect 26976 71130 27028 71136
rect 27080 70922 27108 91598
rect 28276 89962 28304 97106
rect 29184 96960 29236 96966
rect 29184 96902 29236 96908
rect 28264 89956 28316 89962
rect 28264 89898 28316 89904
rect 28276 89714 28304 89898
rect 28184 89686 28304 89714
rect 28184 89010 28212 89686
rect 28172 89004 28224 89010
rect 28172 88946 28224 88952
rect 27896 87372 27948 87378
rect 27896 87314 27948 87320
rect 27620 81184 27672 81190
rect 27620 81126 27672 81132
rect 27160 71528 27212 71534
rect 27160 71470 27212 71476
rect 27172 70990 27200 71470
rect 27160 70984 27212 70990
rect 27160 70926 27212 70932
rect 27068 70916 27120 70922
rect 27068 70858 27120 70864
rect 26884 68264 26936 68270
rect 26884 68206 26936 68212
rect 27528 67176 27580 67182
rect 27528 67118 27580 67124
rect 27540 66842 27568 67118
rect 27252 66836 27304 66842
rect 27252 66778 27304 66784
rect 27528 66836 27580 66842
rect 27528 66778 27580 66784
rect 27264 63306 27292 66778
rect 27344 65680 27396 65686
rect 27344 65622 27396 65628
rect 27356 65006 27384 65622
rect 27344 65000 27396 65006
rect 27344 64942 27396 64948
rect 27356 64666 27384 64942
rect 27344 64660 27396 64666
rect 27344 64602 27396 64608
rect 27252 63300 27304 63306
rect 27252 63242 27304 63248
rect 27160 56296 27212 56302
rect 27160 56238 27212 56244
rect 26608 56228 26660 56234
rect 26608 56170 26660 56176
rect 26516 56160 26568 56166
rect 26516 56102 26568 56108
rect 26976 56160 27028 56166
rect 26976 56102 27028 56108
rect 26436 51046 26556 51074
rect 26240 38208 26292 38214
rect 26240 38150 26292 38156
rect 26252 38010 26280 38150
rect 26240 38004 26292 38010
rect 26240 37946 26292 37952
rect 26332 37800 26384 37806
rect 26332 37742 26384 37748
rect 26148 29776 26200 29782
rect 26148 29718 26200 29724
rect 26240 29300 26292 29306
rect 26240 29242 26292 29248
rect 26252 29102 26280 29242
rect 26056 29096 26108 29102
rect 26056 29038 26108 29044
rect 26240 29096 26292 29102
rect 26240 29038 26292 29044
rect 26068 28966 26096 29038
rect 26056 28960 26108 28966
rect 26056 28902 26108 28908
rect 25872 19984 25924 19990
rect 25872 19926 25924 19932
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25976 16250 26004 17478
rect 26344 17338 26372 37742
rect 26528 34474 26556 51046
rect 26884 45416 26936 45422
rect 26884 45358 26936 45364
rect 26516 34468 26568 34474
rect 26516 34410 26568 34416
rect 26516 30932 26568 30938
rect 26516 30874 26568 30880
rect 26424 29572 26476 29578
rect 26424 29514 26476 29520
rect 26436 29306 26464 29514
rect 26424 29300 26476 29306
rect 26424 29242 26476 29248
rect 26528 29102 26556 30874
rect 26700 30048 26752 30054
rect 26700 29990 26752 29996
rect 26712 29102 26740 29990
rect 26792 29708 26844 29714
rect 26792 29650 26844 29656
rect 26804 29306 26832 29650
rect 26792 29300 26844 29306
rect 26792 29242 26844 29248
rect 26516 29096 26568 29102
rect 26514 29064 26516 29073
rect 26700 29096 26752 29102
rect 26568 29064 26570 29073
rect 26700 29038 26752 29044
rect 26514 28999 26570 29008
rect 26792 21888 26844 21894
rect 26792 21830 26844 21836
rect 26804 21486 26832 21830
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 26332 17332 26384 17338
rect 26332 17274 26384 17280
rect 25964 16244 26016 16250
rect 25964 16186 26016 16192
rect 26896 6914 26924 45358
rect 26988 41138 27016 56102
rect 27172 53582 27200 56238
rect 27160 53576 27212 53582
rect 27160 53518 27212 53524
rect 27068 46980 27120 46986
rect 27068 46922 27120 46928
rect 26976 41132 27028 41138
rect 26976 41074 27028 41080
rect 26976 21480 27028 21486
rect 26976 21422 27028 21428
rect 26804 6886 26924 6914
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 25780 2576 25832 2582
rect 25780 2518 25832 2524
rect 25884 800 25912 4014
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 26344 2990 26372 3334
rect 26332 2984 26384 2990
rect 26332 2926 26384 2932
rect 26056 2848 26108 2854
rect 26056 2790 26108 2796
rect 26068 800 26096 2790
rect 26436 2394 26464 4626
rect 26516 4072 26568 4078
rect 26516 4014 26568 4020
rect 26344 2366 26464 2394
rect 26344 800 26372 2366
rect 26528 800 26556 4014
rect 26700 3460 26752 3466
rect 26700 3402 26752 3408
rect 26712 800 26740 3402
rect 26804 2650 26832 6886
rect 26884 4684 26936 4690
rect 26884 4626 26936 4632
rect 26792 2644 26844 2650
rect 26792 2586 26844 2592
rect 26896 800 26924 4626
rect 26988 3670 27016 21422
rect 27080 9586 27108 46922
rect 27172 11218 27200 53518
rect 27528 47660 27580 47666
rect 27528 47602 27580 47608
rect 27540 47462 27568 47602
rect 27528 47456 27580 47462
rect 27528 47398 27580 47404
rect 27540 46986 27568 47398
rect 27528 46980 27580 46986
rect 27528 46922 27580 46928
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 27068 9580 27120 9586
rect 27068 9522 27120 9528
rect 27632 6914 27660 81126
rect 27908 78606 27936 87314
rect 28448 87304 28500 87310
rect 28448 87246 28500 87252
rect 27896 78600 27948 78606
rect 27896 78542 27948 78548
rect 27908 73234 27936 78542
rect 28460 77722 28488 87246
rect 29196 79762 29224 96902
rect 29276 90024 29328 90030
rect 29276 89966 29328 89972
rect 29460 90024 29512 90030
rect 29460 89966 29512 89972
rect 29288 87718 29316 89966
rect 29276 87712 29328 87718
rect 29276 87654 29328 87660
rect 29288 87378 29316 87654
rect 29276 87372 29328 87378
rect 29276 87314 29328 87320
rect 29368 86964 29420 86970
rect 29368 86906 29420 86912
rect 29380 86766 29408 86906
rect 29368 86760 29420 86766
rect 29368 86702 29420 86708
rect 29380 80102 29408 86702
rect 29368 80096 29420 80102
rect 29368 80038 29420 80044
rect 29184 79756 29236 79762
rect 29184 79698 29236 79704
rect 29184 79552 29236 79558
rect 29184 79494 29236 79500
rect 28540 79144 28592 79150
rect 28540 79086 28592 79092
rect 28448 77716 28500 77722
rect 28448 77658 28500 77664
rect 27896 73228 27948 73234
rect 27896 73170 27948 73176
rect 28264 69352 28316 69358
rect 28264 69294 28316 69300
rect 27712 60172 27764 60178
rect 27712 60114 27764 60120
rect 27724 59022 27752 60114
rect 27712 59016 27764 59022
rect 27712 58958 27764 58964
rect 28172 59016 28224 59022
rect 28172 58958 28224 58964
rect 27712 53712 27764 53718
rect 27712 53654 27764 53660
rect 27724 12442 27752 53654
rect 27804 50380 27856 50386
rect 27804 50322 27856 50328
rect 27816 29714 27844 50322
rect 28184 47666 28212 58958
rect 28276 53718 28304 69294
rect 28460 64874 28488 77658
rect 28552 75274 28580 79086
rect 29196 76974 29224 79494
rect 28816 76968 28868 76974
rect 28816 76910 28868 76916
rect 29184 76968 29236 76974
rect 29184 76910 29236 76916
rect 29368 76968 29420 76974
rect 29368 76910 29420 76916
rect 28540 75268 28592 75274
rect 28540 75210 28592 75216
rect 28632 64932 28684 64938
rect 28632 64874 28684 64880
rect 28368 64846 28488 64874
rect 28368 63578 28396 64846
rect 28356 63572 28408 63578
rect 28356 63514 28408 63520
rect 28356 63436 28408 63442
rect 28356 63378 28408 63384
rect 28264 53712 28316 53718
rect 28264 53654 28316 53660
rect 28276 53174 28304 53654
rect 28264 53168 28316 53174
rect 28264 53110 28316 53116
rect 28368 50726 28396 63378
rect 28356 50720 28408 50726
rect 28356 50662 28408 50668
rect 28368 50386 28396 50662
rect 28356 50380 28408 50386
rect 28356 50322 28408 50328
rect 28448 49360 28500 49366
rect 28448 49302 28500 49308
rect 28460 47802 28488 49302
rect 28448 47796 28500 47802
rect 28448 47738 28500 47744
rect 28172 47660 28224 47666
rect 28172 47602 28224 47608
rect 27988 47592 28040 47598
rect 27988 47534 28040 47540
rect 28000 29714 28028 47534
rect 28264 39840 28316 39846
rect 28264 39782 28316 39788
rect 28276 39642 28304 39782
rect 28264 39636 28316 39642
rect 28264 39578 28316 39584
rect 27804 29708 27856 29714
rect 27804 29650 27856 29656
rect 27988 29708 28040 29714
rect 27988 29650 28040 29656
rect 28000 26234 28028 29650
rect 28644 27674 28672 64874
rect 28828 47802 28856 76910
rect 29276 67584 29328 67590
rect 29276 67526 29328 67532
rect 29288 67114 29316 67526
rect 29276 67108 29328 67114
rect 29276 67050 29328 67056
rect 28816 47796 28868 47802
rect 28816 47738 28868 47744
rect 29288 41682 29316 67050
rect 29276 41676 29328 41682
rect 29276 41618 29328 41624
rect 28724 39976 28776 39982
rect 28724 39918 28776 39924
rect 28632 27668 28684 27674
rect 28632 27610 28684 27616
rect 28736 26234 28764 39918
rect 29000 34944 29052 34950
rect 29000 34886 29052 34892
rect 29012 34746 29040 34886
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 28908 27668 28960 27674
rect 28908 27610 28960 27616
rect 28920 27062 28948 27610
rect 28908 27056 28960 27062
rect 28908 26998 28960 27004
rect 28000 26206 28304 26234
rect 27804 25492 27856 25498
rect 27804 25434 27856 25440
rect 27712 12436 27764 12442
rect 27712 12378 27764 12384
rect 27712 11620 27764 11626
rect 27712 11562 27764 11568
rect 27724 11218 27752 11562
rect 27712 11212 27764 11218
rect 27712 11154 27764 11160
rect 27448 6886 27660 6914
rect 26976 3664 27028 3670
rect 26976 3606 27028 3612
rect 27068 3596 27120 3602
rect 27068 3538 27120 3544
rect 27080 800 27108 3538
rect 27344 2848 27396 2854
rect 27344 2790 27396 2796
rect 27356 800 27384 2790
rect 27448 2514 27476 6886
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 27540 800 27568 4014
rect 27816 3194 27844 25434
rect 28276 21554 28304 26206
rect 28552 26206 28764 26234
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 28356 21548 28408 21554
rect 28356 21490 28408 21496
rect 28172 20256 28224 20262
rect 28172 20198 28224 20204
rect 28184 19922 28212 20198
rect 28172 19916 28224 19922
rect 28172 19858 28224 19864
rect 28368 18290 28396 21490
rect 28552 19174 28580 26206
rect 28816 21684 28868 21690
rect 28816 21626 28868 21632
rect 28632 21412 28684 21418
rect 28632 21354 28684 21360
rect 28540 19168 28592 19174
rect 28540 19110 28592 19116
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 27988 12436 28040 12442
rect 27988 12378 28040 12384
rect 28000 11286 28028 12378
rect 27988 11280 28040 11286
rect 27988 11222 28040 11228
rect 28080 3596 28132 3602
rect 28080 3538 28132 3544
rect 27804 3188 27856 3194
rect 27804 3130 27856 3136
rect 27816 2990 27844 3130
rect 27804 2984 27856 2990
rect 27804 2926 27856 2932
rect 27712 2916 27764 2922
rect 27712 2858 27764 2864
rect 27724 800 27752 2858
rect 27896 2372 27948 2378
rect 27896 2314 27948 2320
rect 27908 800 27936 2314
rect 28092 800 28120 3538
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 28368 800 28396 2790
rect 28644 2650 28672 21354
rect 28724 4072 28776 4078
rect 28724 4014 28776 4020
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 28540 2372 28592 2378
rect 28540 2314 28592 2320
rect 28552 800 28580 2314
rect 28736 800 28764 4014
rect 28828 2650 28856 21626
rect 29000 18896 29052 18902
rect 29000 18838 29052 18844
rect 29012 16114 29040 18838
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29380 13802 29408 76910
rect 29472 59770 29500 89966
rect 29736 86760 29788 86766
rect 29736 86702 29788 86708
rect 29644 80232 29696 80238
rect 29644 80174 29696 80180
rect 29656 80054 29684 80174
rect 29564 80026 29684 80054
rect 29564 64394 29592 80026
rect 29644 76832 29696 76838
rect 29644 76774 29696 76780
rect 29552 64388 29604 64394
rect 29552 64330 29604 64336
rect 29460 59764 29512 59770
rect 29460 59706 29512 59712
rect 29552 52012 29604 52018
rect 29552 51954 29604 51960
rect 29564 39506 29592 51954
rect 29552 39500 29604 39506
rect 29552 39442 29604 39448
rect 29552 23112 29604 23118
rect 29552 23054 29604 23060
rect 29368 13796 29420 13802
rect 29368 13738 29420 13744
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 28920 8090 28948 13126
rect 28908 8084 28960 8090
rect 28908 8026 28960 8032
rect 29564 6914 29592 23054
rect 29656 7206 29684 76774
rect 29748 60518 29776 86702
rect 29736 60512 29788 60518
rect 29736 60454 29788 60460
rect 29840 43314 29868 97106
rect 30380 96484 30432 96490
rect 30380 96426 30432 96432
rect 30288 96076 30340 96082
rect 30288 96018 30340 96024
rect 30300 90030 30328 96018
rect 30392 96014 30420 96426
rect 30380 96008 30432 96014
rect 30380 95950 30432 95956
rect 30288 90024 30340 90030
rect 30288 89966 30340 89972
rect 30300 89714 30328 89966
rect 30208 89686 30328 89714
rect 30208 86970 30236 89686
rect 30196 86964 30248 86970
rect 30196 86906 30248 86912
rect 30392 85542 30420 95950
rect 30656 95940 30708 95946
rect 30656 95882 30708 95888
rect 30380 85536 30432 85542
rect 30380 85478 30432 85484
rect 30012 85264 30064 85270
rect 30012 85206 30064 85212
rect 29920 81184 29972 81190
rect 29920 81126 29972 81132
rect 29932 67590 29960 81126
rect 29920 67584 29972 67590
rect 29920 67526 29972 67532
rect 29920 51400 29972 51406
rect 29920 51342 29972 51348
rect 29828 43308 29880 43314
rect 29828 43250 29880 43256
rect 29736 39840 29788 39846
rect 29736 39782 29788 39788
rect 29748 18902 29776 39782
rect 29736 18896 29788 18902
rect 29736 18838 29788 18844
rect 29736 13796 29788 13802
rect 29736 13738 29788 13744
rect 29748 12646 29776 13738
rect 29736 12640 29788 12646
rect 29736 12582 29788 12588
rect 29644 7200 29696 7206
rect 29644 7142 29696 7148
rect 29564 6886 29684 6914
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28816 2644 28868 2650
rect 28816 2586 28868 2592
rect 28920 800 28948 3538
rect 29092 2372 29144 2378
rect 29092 2314 29144 2320
rect 29104 800 29132 2314
rect 29380 800 29408 4014
rect 29552 2984 29604 2990
rect 29552 2926 29604 2932
rect 29564 800 29592 2926
rect 29656 2650 29684 6886
rect 29748 4282 29776 12582
rect 29932 7750 29960 51342
rect 30024 30938 30052 85206
rect 30392 85134 30420 85478
rect 30380 85128 30432 85134
rect 30380 85070 30432 85076
rect 30472 79688 30524 79694
rect 30472 79630 30524 79636
rect 30380 79552 30432 79558
rect 30380 79494 30432 79500
rect 30392 79286 30420 79494
rect 30380 79280 30432 79286
rect 30380 79222 30432 79228
rect 30392 78606 30420 79222
rect 30484 79218 30512 79630
rect 30472 79212 30524 79218
rect 30472 79154 30524 79160
rect 30484 78674 30512 79154
rect 30472 78668 30524 78674
rect 30472 78610 30524 78616
rect 30380 78600 30432 78606
rect 30380 78542 30432 78548
rect 30564 76492 30616 76498
rect 30564 76434 30616 76440
rect 30576 75818 30604 76434
rect 30564 75812 30616 75818
rect 30564 75754 30616 75760
rect 30668 61810 30696 95882
rect 30748 90024 30800 90030
rect 30748 89966 30800 89972
rect 30656 61804 30708 61810
rect 30656 61746 30708 61752
rect 30288 59764 30340 59770
rect 30288 59706 30340 59712
rect 30196 52420 30248 52426
rect 30196 52362 30248 52368
rect 30104 48884 30156 48890
rect 30104 48826 30156 48832
rect 30012 30932 30064 30938
rect 30012 30874 30064 30880
rect 30116 10470 30144 48826
rect 30208 20466 30236 52362
rect 30300 32570 30328 59706
rect 30380 50312 30432 50318
rect 30380 50254 30432 50260
rect 30392 49774 30420 50254
rect 30380 49768 30432 49774
rect 30380 49710 30432 49716
rect 30564 49768 30616 49774
rect 30564 49710 30616 49716
rect 30380 34468 30432 34474
rect 30380 34410 30432 34416
rect 30288 32564 30340 32570
rect 30288 32506 30340 32512
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 30196 18216 30248 18222
rect 30196 18158 30248 18164
rect 30208 11898 30236 18158
rect 30196 11892 30248 11898
rect 30196 11834 30248 11840
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 29920 7744 29972 7750
rect 29920 7686 29972 7692
rect 29736 4276 29788 4282
rect 29736 4218 29788 4224
rect 29920 3596 29972 3602
rect 29920 3538 29972 3544
rect 29644 2644 29696 2650
rect 29644 2586 29696 2592
rect 29828 2372 29880 2378
rect 29828 2314 29880 2320
rect 29840 1170 29868 2314
rect 29748 1142 29868 1170
rect 29748 800 29776 1142
rect 29932 800 29960 3538
rect 30104 2984 30156 2990
rect 30104 2926 30156 2932
rect 30116 800 30144 2926
rect 30392 2650 30420 34410
rect 30576 24818 30604 49710
rect 30760 32366 30788 89966
rect 30840 80164 30892 80170
rect 30840 80106 30892 80112
rect 30852 72078 30880 80106
rect 31036 79898 31064 97106
rect 31852 96960 31904 96966
rect 31852 96902 31904 96908
rect 31392 95396 31444 95402
rect 31392 95338 31444 95344
rect 31116 89548 31168 89554
rect 31116 89490 31168 89496
rect 31024 79892 31076 79898
rect 31024 79834 31076 79840
rect 31128 78470 31156 89490
rect 31300 85536 31352 85542
rect 31300 85478 31352 85484
rect 31208 83564 31260 83570
rect 31208 83506 31260 83512
rect 31116 78464 31168 78470
rect 31116 78406 31168 78412
rect 31116 76424 31168 76430
rect 31116 76366 31168 76372
rect 30840 72072 30892 72078
rect 30840 72014 30892 72020
rect 30852 67318 30880 72014
rect 30840 67312 30892 67318
rect 30840 67254 30892 67260
rect 30840 61736 30892 61742
rect 30840 61678 30892 61684
rect 30852 61334 30880 61678
rect 30840 61328 30892 61334
rect 30840 61270 30892 61276
rect 31024 43784 31076 43790
rect 31024 43726 31076 43732
rect 31036 39914 31064 43726
rect 31024 39908 31076 39914
rect 31024 39850 31076 39856
rect 31036 38350 31064 39850
rect 31128 39642 31156 76366
rect 31116 39636 31168 39642
rect 31116 39578 31168 39584
rect 31024 38344 31076 38350
rect 31024 38286 31076 38292
rect 31036 35086 31064 38286
rect 31024 35080 31076 35086
rect 31024 35022 31076 35028
rect 31036 33454 31064 35022
rect 31128 33930 31156 39578
rect 31116 33924 31168 33930
rect 31116 33866 31168 33872
rect 31024 33448 31076 33454
rect 31024 33390 31076 33396
rect 31220 33318 31248 83506
rect 31312 70394 31340 85478
rect 31404 80646 31432 95338
rect 31864 85338 31892 96902
rect 31944 89888 31996 89894
rect 31944 89830 31996 89836
rect 31852 85332 31904 85338
rect 31852 85274 31904 85280
rect 31392 80640 31444 80646
rect 31392 80582 31444 80588
rect 31404 76498 31432 80582
rect 31392 76492 31444 76498
rect 31392 76434 31444 76440
rect 31312 70366 31432 70394
rect 31404 68338 31432 70366
rect 31392 68332 31444 68338
rect 31392 68274 31444 68280
rect 31392 61736 31444 61742
rect 31392 61678 31444 61684
rect 31300 41608 31352 41614
rect 31300 41550 31352 41556
rect 31208 33312 31260 33318
rect 31208 33254 31260 33260
rect 30748 32360 30800 32366
rect 30748 32302 30800 32308
rect 31312 30938 31340 41550
rect 31404 35086 31432 61678
rect 31668 61600 31720 61606
rect 31668 61542 31720 61548
rect 31576 49632 31628 49638
rect 31576 49574 31628 49580
rect 31588 49366 31616 49574
rect 31576 49360 31628 49366
rect 31576 49302 31628 49308
rect 31484 47252 31536 47258
rect 31484 47194 31536 47200
rect 31496 38350 31524 47194
rect 31576 39500 31628 39506
rect 31576 39442 31628 39448
rect 31484 38344 31536 38350
rect 31484 38286 31536 38292
rect 31484 35488 31536 35494
rect 31484 35430 31536 35436
rect 31392 35080 31444 35086
rect 31392 35022 31444 35028
rect 31116 30932 31168 30938
rect 31116 30874 31168 30880
rect 31300 30932 31352 30938
rect 31300 30874 31352 30880
rect 31128 26234 31156 30874
rect 31036 26206 31156 26234
rect 30564 24812 30616 24818
rect 30564 24754 30616 24760
rect 31036 13394 31064 26206
rect 31404 24138 31432 35022
rect 31392 24132 31444 24138
rect 31392 24074 31444 24080
rect 31116 17536 31168 17542
rect 31116 17478 31168 17484
rect 31024 13388 31076 13394
rect 31024 13330 31076 13336
rect 31128 7818 31156 17478
rect 31116 7812 31168 7818
rect 31116 7754 31168 7760
rect 30564 4072 30616 4078
rect 30564 4014 30616 4020
rect 31208 4072 31260 4078
rect 31208 4014 31260 4020
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 30392 800 30420 2382
rect 30576 800 30604 4014
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 30760 800 30788 2926
rect 31024 2372 31076 2378
rect 31024 2314 31076 2320
rect 31036 1170 31064 2314
rect 30944 1142 31064 1170
rect 30944 800 30972 1142
rect 31220 800 31248 4014
rect 31392 2984 31444 2990
rect 31392 2926 31444 2932
rect 31404 800 31432 2926
rect 31496 2650 31524 35430
rect 31588 3670 31616 39442
rect 31680 23662 31708 61542
rect 31760 60648 31812 60654
rect 31760 60590 31812 60596
rect 31772 56506 31800 60590
rect 31760 56500 31812 56506
rect 31760 56442 31812 56448
rect 31760 49768 31812 49774
rect 31760 49710 31812 49716
rect 31772 40594 31800 49710
rect 31760 40588 31812 40594
rect 31760 40530 31812 40536
rect 31956 33114 31984 89830
rect 32508 87922 32536 97106
rect 33428 96626 33456 99200
rect 34256 97170 34284 99200
rect 35176 97306 35204 99200
rect 35164 97300 35216 97306
rect 35164 97242 35216 97248
rect 34244 97164 34296 97170
rect 34244 97106 34296 97112
rect 34796 97164 34848 97170
rect 34796 97106 34848 97112
rect 34612 96756 34664 96762
rect 34612 96698 34664 96704
rect 33416 96620 33468 96626
rect 33416 96562 33468 96568
rect 34520 93220 34572 93226
rect 34520 93162 34572 93168
rect 32496 87916 32548 87922
rect 32496 87858 32548 87864
rect 32508 84194 32536 87858
rect 34532 86834 34560 93162
rect 34520 86828 34572 86834
rect 34520 86770 34572 86776
rect 32588 85196 32640 85202
rect 32588 85138 32640 85144
rect 32416 84166 32536 84194
rect 32416 62422 32444 84166
rect 32600 81258 32628 85138
rect 34152 84992 34204 84998
rect 34152 84934 34204 84940
rect 32496 81252 32548 81258
rect 32496 81194 32548 81200
rect 32588 81252 32640 81258
rect 32588 81194 32640 81200
rect 32508 74458 32536 81194
rect 32600 76906 32628 81194
rect 32588 76900 32640 76906
rect 32588 76842 32640 76848
rect 32496 74452 32548 74458
rect 32496 74394 32548 74400
rect 32404 62416 32456 62422
rect 32404 62358 32456 62364
rect 32404 53984 32456 53990
rect 32404 53926 32456 53932
rect 32220 50312 32272 50318
rect 32220 50254 32272 50260
rect 31944 33108 31996 33114
rect 31944 33050 31996 33056
rect 32232 30870 32260 50254
rect 32416 44878 32444 53926
rect 32404 44872 32456 44878
rect 32404 44814 32456 44820
rect 32404 40588 32456 40594
rect 32404 40530 32456 40536
rect 32220 30864 32272 30870
rect 32220 30806 32272 30812
rect 31668 23656 31720 23662
rect 31668 23598 31720 23604
rect 31668 18216 31720 18222
rect 31668 18158 31720 18164
rect 31680 15434 31708 18158
rect 31668 15428 31720 15434
rect 31668 15370 31720 15376
rect 31680 11558 31708 15370
rect 31668 11552 31720 11558
rect 31668 11494 31720 11500
rect 32416 4826 32444 40530
rect 32508 39438 32536 74394
rect 33876 69352 33928 69358
rect 33876 69294 33928 69300
rect 33784 65544 33836 65550
rect 33784 65486 33836 65492
rect 33796 63850 33824 65486
rect 33784 63844 33836 63850
rect 33784 63786 33836 63792
rect 33796 62830 33824 63786
rect 33784 62824 33836 62830
rect 33784 62766 33836 62772
rect 33692 62688 33744 62694
rect 33692 62630 33744 62636
rect 33704 62490 33732 62630
rect 33692 62484 33744 62490
rect 33692 62426 33744 62432
rect 33784 59968 33836 59974
rect 33784 59910 33836 59916
rect 32588 54528 32640 54534
rect 32588 54470 32640 54476
rect 32496 39432 32548 39438
rect 32496 39374 32548 39380
rect 32508 12850 32536 39374
rect 32600 16574 32628 54470
rect 33796 52494 33824 59910
rect 33784 52488 33836 52494
rect 33784 52430 33836 52436
rect 32956 50720 33008 50726
rect 32956 50662 33008 50668
rect 33600 50720 33652 50726
rect 33600 50662 33652 50668
rect 32968 50454 32996 50662
rect 32956 50448 33008 50454
rect 32956 50390 33008 50396
rect 33612 50386 33640 50662
rect 33600 50380 33652 50386
rect 33600 50322 33652 50328
rect 33416 50176 33468 50182
rect 33416 50118 33468 50124
rect 32864 39840 32916 39846
rect 32864 39782 32916 39788
rect 32876 39370 32904 39782
rect 32956 39500 33008 39506
rect 32956 39442 33008 39448
rect 32864 39364 32916 39370
rect 32864 39306 32916 39312
rect 32600 16546 32720 16574
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 32404 4820 32456 4826
rect 32404 4762 32456 4768
rect 31760 4072 31812 4078
rect 31760 4014 31812 4020
rect 31576 3664 31628 3670
rect 31576 3606 31628 3612
rect 31484 2644 31536 2650
rect 31484 2586 31536 2592
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 31588 800 31616 2246
rect 31772 800 31800 4014
rect 31944 3596 31996 3602
rect 31944 3538 31996 3544
rect 32496 3596 32548 3602
rect 32496 3538 32548 3544
rect 31956 800 31984 3538
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 32232 800 32260 2382
rect 32508 1850 32536 3538
rect 32588 2984 32640 2990
rect 32588 2926 32640 2932
rect 32416 1822 32536 1850
rect 32416 800 32444 1822
rect 32600 800 32628 2926
rect 32692 2582 32720 16546
rect 32876 8498 32904 39306
rect 32968 26586 32996 39442
rect 33048 38820 33100 38826
rect 33048 38762 33100 38768
rect 33060 38554 33088 38762
rect 33048 38548 33100 38554
rect 33048 38490 33100 38496
rect 33324 34536 33376 34542
rect 33324 34478 33376 34484
rect 33048 33856 33100 33862
rect 33048 33798 33100 33804
rect 33060 33454 33088 33798
rect 33336 33454 33364 34478
rect 33048 33448 33100 33454
rect 33048 33390 33100 33396
rect 33324 33448 33376 33454
rect 33324 33390 33376 33396
rect 33428 31142 33456 50118
rect 33692 39636 33744 39642
rect 33692 39578 33744 39584
rect 33600 39500 33652 39506
rect 33600 39442 33652 39448
rect 33508 39432 33560 39438
rect 33508 39374 33560 39380
rect 33520 39098 33548 39374
rect 33508 39092 33560 39098
rect 33508 39034 33560 39040
rect 33612 38962 33640 39442
rect 33704 39438 33732 39578
rect 33692 39432 33744 39438
rect 33692 39374 33744 39380
rect 33600 38956 33652 38962
rect 33600 38898 33652 38904
rect 33704 36854 33732 39374
rect 33692 36848 33744 36854
rect 33692 36790 33744 36796
rect 33416 31136 33468 31142
rect 33416 31078 33468 31084
rect 32956 26580 33008 26586
rect 32956 26522 33008 26528
rect 33784 21956 33836 21962
rect 33784 21898 33836 21904
rect 33692 17196 33744 17202
rect 33692 17138 33744 17144
rect 32864 8492 32916 8498
rect 32864 8434 32916 8440
rect 33600 4072 33652 4078
rect 33600 4014 33652 4020
rect 32956 3528 33008 3534
rect 32956 3470 33008 3476
rect 32680 2576 32732 2582
rect 32680 2518 32732 2524
rect 32772 2372 32824 2378
rect 32772 2314 32824 2320
rect 32784 800 32812 2314
rect 32968 800 32996 3470
rect 33232 2984 33284 2990
rect 33232 2926 33284 2932
rect 33244 800 33272 2926
rect 33416 2508 33468 2514
rect 33416 2450 33468 2456
rect 33428 800 33456 2450
rect 33612 800 33640 4014
rect 33704 2582 33732 17138
rect 33796 11626 33824 21898
rect 33888 21486 33916 69294
rect 33968 67312 34020 67318
rect 33968 67254 34020 67260
rect 33980 60246 34008 67254
rect 34164 66842 34192 84934
rect 34152 66836 34204 66842
rect 34152 66778 34204 66784
rect 34164 64874 34192 66778
rect 34072 64846 34192 64874
rect 33968 60240 34020 60246
rect 33968 60182 34020 60188
rect 33980 56302 34008 60182
rect 33968 56296 34020 56302
rect 33968 56238 34020 56244
rect 33980 54670 34008 56238
rect 33968 54664 34020 54670
rect 33968 54606 34020 54612
rect 33968 52488 34020 52494
rect 33968 52430 34020 52436
rect 33980 39506 34008 52430
rect 34072 48278 34100 64846
rect 34152 64116 34204 64122
rect 34152 64058 34204 64064
rect 34164 63578 34192 64058
rect 34152 63572 34204 63578
rect 34152 63514 34204 63520
rect 34164 62830 34192 63514
rect 34244 63232 34296 63238
rect 34244 63174 34296 63180
rect 34152 62824 34204 62830
rect 34152 62766 34204 62772
rect 34256 62762 34284 63174
rect 34520 62824 34572 62830
rect 34520 62766 34572 62772
rect 34244 62756 34296 62762
rect 34244 62698 34296 62704
rect 34152 62688 34204 62694
rect 34152 62630 34204 62636
rect 34336 62688 34388 62694
rect 34336 62630 34388 62636
rect 34164 62422 34192 62630
rect 34152 62416 34204 62422
rect 34152 62358 34204 62364
rect 34152 60104 34204 60110
rect 34152 60046 34204 60052
rect 34060 48272 34112 48278
rect 34060 48214 34112 48220
rect 34060 39840 34112 39846
rect 34060 39782 34112 39788
rect 34072 39574 34100 39782
rect 34164 39642 34192 60046
rect 34348 55622 34376 62630
rect 34532 62490 34560 62766
rect 34520 62484 34572 62490
rect 34520 62426 34572 62432
rect 34520 60036 34572 60042
rect 34520 59978 34572 59984
rect 34336 55616 34388 55622
rect 34336 55558 34388 55564
rect 34428 54664 34480 54670
rect 34428 54606 34480 54612
rect 34440 50726 34468 54606
rect 34428 50720 34480 50726
rect 34428 50662 34480 50668
rect 34336 46912 34388 46918
rect 34336 46854 34388 46860
rect 34348 46102 34376 46854
rect 34336 46096 34388 46102
rect 34336 46038 34388 46044
rect 34244 40112 34296 40118
rect 34244 40054 34296 40060
rect 34152 39636 34204 39642
rect 34152 39578 34204 39584
rect 34060 39568 34112 39574
rect 34060 39510 34112 39516
rect 33968 39500 34020 39506
rect 33968 39442 34020 39448
rect 34060 38208 34112 38214
rect 34060 38150 34112 38156
rect 33876 21480 33928 21486
rect 33876 21422 33928 21428
rect 33968 21412 34020 21418
rect 33968 21354 34020 21360
rect 33980 14890 34008 21354
rect 34072 17678 34100 38150
rect 34152 32836 34204 32842
rect 34152 32778 34204 32784
rect 34060 17672 34112 17678
rect 34060 17614 34112 17620
rect 33968 14884 34020 14890
rect 33968 14826 34020 14832
rect 33784 11620 33836 11626
rect 33784 11562 33836 11568
rect 33784 2984 33836 2990
rect 33784 2926 33836 2932
rect 33692 2576 33744 2582
rect 33692 2518 33744 2524
rect 33796 800 33824 2926
rect 34164 2650 34192 32778
rect 34256 17542 34284 40054
rect 34348 21962 34376 46038
rect 34428 41200 34480 41206
rect 34428 41142 34480 41148
rect 34440 40458 34468 41142
rect 34428 40452 34480 40458
rect 34428 40394 34480 40400
rect 34440 39982 34468 40394
rect 34428 39976 34480 39982
rect 34428 39918 34480 39924
rect 34532 39098 34560 59978
rect 34624 39982 34652 96698
rect 34808 87786 34836 97106
rect 34940 96860 35236 96880
rect 34996 96858 35020 96860
rect 35076 96858 35100 96860
rect 35156 96858 35180 96860
rect 35018 96806 35020 96858
rect 35082 96806 35094 96858
rect 35156 96806 35158 96858
rect 34996 96804 35020 96806
rect 35076 96804 35100 96806
rect 35156 96804 35180 96806
rect 34940 96784 35236 96804
rect 36004 96626 36032 99200
rect 36832 97238 36860 99200
rect 37752 97306 37780 99200
rect 37740 97300 37792 97306
rect 37740 97242 37792 97248
rect 36820 97232 36872 97238
rect 36820 97174 36872 97180
rect 37832 97164 37884 97170
rect 37832 97106 37884 97112
rect 37096 96960 37148 96966
rect 37096 96902 37148 96908
rect 35992 96620 36044 96626
rect 35992 96562 36044 96568
rect 36084 96484 36136 96490
rect 36084 96426 36136 96432
rect 34940 95772 35236 95792
rect 34996 95770 35020 95772
rect 35076 95770 35100 95772
rect 35156 95770 35180 95772
rect 35018 95718 35020 95770
rect 35082 95718 35094 95770
rect 35156 95718 35158 95770
rect 34996 95716 35020 95718
rect 35076 95716 35100 95718
rect 35156 95716 35180 95718
rect 34940 95696 35236 95716
rect 35348 95464 35400 95470
rect 35348 95406 35400 95412
rect 34940 94684 35236 94704
rect 34996 94682 35020 94684
rect 35076 94682 35100 94684
rect 35156 94682 35180 94684
rect 35018 94630 35020 94682
rect 35082 94630 35094 94682
rect 35156 94630 35158 94682
rect 34996 94628 35020 94630
rect 35076 94628 35100 94630
rect 35156 94628 35180 94630
rect 34940 94608 35236 94628
rect 34940 93596 35236 93616
rect 34996 93594 35020 93596
rect 35076 93594 35100 93596
rect 35156 93594 35180 93596
rect 35018 93542 35020 93594
rect 35082 93542 35094 93594
rect 35156 93542 35158 93594
rect 34996 93540 35020 93542
rect 35076 93540 35100 93542
rect 35156 93540 35180 93542
rect 34940 93520 35236 93540
rect 35360 93226 35388 95406
rect 35348 93220 35400 93226
rect 35348 93162 35400 93168
rect 34940 92508 35236 92528
rect 34996 92506 35020 92508
rect 35076 92506 35100 92508
rect 35156 92506 35180 92508
rect 35018 92454 35020 92506
rect 35082 92454 35094 92506
rect 35156 92454 35158 92506
rect 34996 92452 35020 92454
rect 35076 92452 35100 92454
rect 35156 92452 35180 92454
rect 34940 92432 35236 92452
rect 35440 92132 35492 92138
rect 35440 92074 35492 92080
rect 34940 91420 35236 91440
rect 34996 91418 35020 91420
rect 35076 91418 35100 91420
rect 35156 91418 35180 91420
rect 35018 91366 35020 91418
rect 35082 91366 35094 91418
rect 35156 91366 35158 91418
rect 34996 91364 35020 91366
rect 35076 91364 35100 91366
rect 35156 91364 35180 91366
rect 34940 91344 35236 91364
rect 34940 90332 35236 90352
rect 34996 90330 35020 90332
rect 35076 90330 35100 90332
rect 35156 90330 35180 90332
rect 35018 90278 35020 90330
rect 35082 90278 35094 90330
rect 35156 90278 35158 90330
rect 34996 90276 35020 90278
rect 35076 90276 35100 90278
rect 35156 90276 35180 90278
rect 34940 90256 35236 90276
rect 34940 89244 35236 89264
rect 34996 89242 35020 89244
rect 35076 89242 35100 89244
rect 35156 89242 35180 89244
rect 35018 89190 35020 89242
rect 35082 89190 35094 89242
rect 35156 89190 35158 89242
rect 34996 89188 35020 89190
rect 35076 89188 35100 89190
rect 35156 89188 35180 89190
rect 34940 89168 35236 89188
rect 34940 88156 35236 88176
rect 34996 88154 35020 88156
rect 35076 88154 35100 88156
rect 35156 88154 35180 88156
rect 35018 88102 35020 88154
rect 35082 88102 35094 88154
rect 35156 88102 35158 88154
rect 34996 88100 35020 88102
rect 35076 88100 35100 88102
rect 35156 88100 35180 88102
rect 34940 88080 35236 88100
rect 34796 87780 34848 87786
rect 34796 87722 34848 87728
rect 35256 87168 35308 87174
rect 35256 87110 35308 87116
rect 34940 87068 35236 87088
rect 34996 87066 35020 87068
rect 35076 87066 35100 87068
rect 35156 87066 35180 87068
rect 35018 87014 35020 87066
rect 35082 87014 35094 87066
rect 35156 87014 35158 87066
rect 34996 87012 35020 87014
rect 35076 87012 35100 87014
rect 35156 87012 35180 87014
rect 34940 86992 35236 87012
rect 34940 85980 35236 86000
rect 34996 85978 35020 85980
rect 35076 85978 35100 85980
rect 35156 85978 35180 85980
rect 35018 85926 35020 85978
rect 35082 85926 35094 85978
rect 35156 85926 35158 85978
rect 34996 85924 35020 85926
rect 35076 85924 35100 85926
rect 35156 85924 35180 85926
rect 34940 85904 35236 85924
rect 34940 84892 35236 84912
rect 34996 84890 35020 84892
rect 35076 84890 35100 84892
rect 35156 84890 35180 84892
rect 35018 84838 35020 84890
rect 35082 84838 35094 84890
rect 35156 84838 35158 84890
rect 34996 84836 35020 84838
rect 35076 84836 35100 84838
rect 35156 84836 35180 84838
rect 34940 84816 35236 84836
rect 34940 83804 35236 83824
rect 34996 83802 35020 83804
rect 35076 83802 35100 83804
rect 35156 83802 35180 83804
rect 35018 83750 35020 83802
rect 35082 83750 35094 83802
rect 35156 83750 35158 83802
rect 34996 83748 35020 83750
rect 35076 83748 35100 83750
rect 35156 83748 35180 83750
rect 34940 83728 35236 83748
rect 34940 82716 35236 82736
rect 34996 82714 35020 82716
rect 35076 82714 35100 82716
rect 35156 82714 35180 82716
rect 35018 82662 35020 82714
rect 35082 82662 35094 82714
rect 35156 82662 35158 82714
rect 34996 82660 35020 82662
rect 35076 82660 35100 82662
rect 35156 82660 35180 82662
rect 34940 82640 35236 82660
rect 34940 81628 35236 81648
rect 34996 81626 35020 81628
rect 35076 81626 35100 81628
rect 35156 81626 35180 81628
rect 35018 81574 35020 81626
rect 35082 81574 35094 81626
rect 35156 81574 35158 81626
rect 34996 81572 35020 81574
rect 35076 81572 35100 81574
rect 35156 81572 35180 81574
rect 34940 81552 35236 81572
rect 34940 80540 35236 80560
rect 34996 80538 35020 80540
rect 35076 80538 35100 80540
rect 35156 80538 35180 80540
rect 35018 80486 35020 80538
rect 35082 80486 35094 80538
rect 35156 80486 35158 80538
rect 34996 80484 35020 80486
rect 35076 80484 35100 80486
rect 35156 80484 35180 80486
rect 34940 80464 35236 80484
rect 34940 79452 35236 79472
rect 34996 79450 35020 79452
rect 35076 79450 35100 79452
rect 35156 79450 35180 79452
rect 35018 79398 35020 79450
rect 35082 79398 35094 79450
rect 35156 79398 35158 79450
rect 34996 79396 35020 79398
rect 35076 79396 35100 79398
rect 35156 79396 35180 79398
rect 34940 79376 35236 79396
rect 34940 78364 35236 78384
rect 34996 78362 35020 78364
rect 35076 78362 35100 78364
rect 35156 78362 35180 78364
rect 35018 78310 35020 78362
rect 35082 78310 35094 78362
rect 35156 78310 35158 78362
rect 34996 78308 35020 78310
rect 35076 78308 35100 78310
rect 35156 78308 35180 78310
rect 34940 78288 35236 78308
rect 34940 77276 35236 77296
rect 34996 77274 35020 77276
rect 35076 77274 35100 77276
rect 35156 77274 35180 77276
rect 35018 77222 35020 77274
rect 35082 77222 35094 77274
rect 35156 77222 35158 77274
rect 34996 77220 35020 77222
rect 35076 77220 35100 77222
rect 35156 77220 35180 77222
rect 34940 77200 35236 77220
rect 34940 76188 35236 76208
rect 34996 76186 35020 76188
rect 35076 76186 35100 76188
rect 35156 76186 35180 76188
rect 35018 76134 35020 76186
rect 35082 76134 35094 76186
rect 35156 76134 35158 76186
rect 34996 76132 35020 76134
rect 35076 76132 35100 76134
rect 35156 76132 35180 76134
rect 34940 76112 35236 76132
rect 34940 75100 35236 75120
rect 34996 75098 35020 75100
rect 35076 75098 35100 75100
rect 35156 75098 35180 75100
rect 35018 75046 35020 75098
rect 35082 75046 35094 75098
rect 35156 75046 35158 75098
rect 34996 75044 35020 75046
rect 35076 75044 35100 75046
rect 35156 75044 35180 75046
rect 34940 75024 35236 75044
rect 34940 74012 35236 74032
rect 34996 74010 35020 74012
rect 35076 74010 35100 74012
rect 35156 74010 35180 74012
rect 35018 73958 35020 74010
rect 35082 73958 35094 74010
rect 35156 73958 35158 74010
rect 34996 73956 35020 73958
rect 35076 73956 35100 73958
rect 35156 73956 35180 73958
rect 34940 73936 35236 73956
rect 34940 72924 35236 72944
rect 34996 72922 35020 72924
rect 35076 72922 35100 72924
rect 35156 72922 35180 72924
rect 35018 72870 35020 72922
rect 35082 72870 35094 72922
rect 35156 72870 35158 72922
rect 34996 72868 35020 72870
rect 35076 72868 35100 72870
rect 35156 72868 35180 72870
rect 34940 72848 35236 72868
rect 34940 71836 35236 71856
rect 34996 71834 35020 71836
rect 35076 71834 35100 71836
rect 35156 71834 35180 71836
rect 35018 71782 35020 71834
rect 35082 71782 35094 71834
rect 35156 71782 35158 71834
rect 34996 71780 35020 71782
rect 35076 71780 35100 71782
rect 35156 71780 35180 71782
rect 34940 71760 35236 71780
rect 34940 70748 35236 70768
rect 34996 70746 35020 70748
rect 35076 70746 35100 70748
rect 35156 70746 35180 70748
rect 35018 70694 35020 70746
rect 35082 70694 35094 70746
rect 35156 70694 35158 70746
rect 34996 70692 35020 70694
rect 35076 70692 35100 70694
rect 35156 70692 35180 70694
rect 34940 70672 35236 70692
rect 34940 69660 35236 69680
rect 34996 69658 35020 69660
rect 35076 69658 35100 69660
rect 35156 69658 35180 69660
rect 35018 69606 35020 69658
rect 35082 69606 35094 69658
rect 35156 69606 35158 69658
rect 34996 69604 35020 69606
rect 35076 69604 35100 69606
rect 35156 69604 35180 69606
rect 34940 69584 35236 69604
rect 34940 68572 35236 68592
rect 34996 68570 35020 68572
rect 35076 68570 35100 68572
rect 35156 68570 35180 68572
rect 35018 68518 35020 68570
rect 35082 68518 35094 68570
rect 35156 68518 35158 68570
rect 34996 68516 35020 68518
rect 35076 68516 35100 68518
rect 35156 68516 35180 68518
rect 34940 68496 35236 68516
rect 34940 67484 35236 67504
rect 34996 67482 35020 67484
rect 35076 67482 35100 67484
rect 35156 67482 35180 67484
rect 35018 67430 35020 67482
rect 35082 67430 35094 67482
rect 35156 67430 35158 67482
rect 34996 67428 35020 67430
rect 35076 67428 35100 67430
rect 35156 67428 35180 67430
rect 34940 67408 35236 67428
rect 35268 67250 35296 87110
rect 35452 75886 35480 92074
rect 35440 75880 35492 75886
rect 35440 75822 35492 75828
rect 35256 67244 35308 67250
rect 35256 67186 35308 67192
rect 34940 66396 35236 66416
rect 34996 66394 35020 66396
rect 35076 66394 35100 66396
rect 35156 66394 35180 66396
rect 35018 66342 35020 66394
rect 35082 66342 35094 66394
rect 35156 66342 35158 66394
rect 34996 66340 35020 66342
rect 35076 66340 35100 66342
rect 35156 66340 35180 66342
rect 34940 66320 35236 66340
rect 34940 65308 35236 65328
rect 34996 65306 35020 65308
rect 35076 65306 35100 65308
rect 35156 65306 35180 65308
rect 35018 65254 35020 65306
rect 35082 65254 35094 65306
rect 35156 65254 35158 65306
rect 34996 65252 35020 65254
rect 35076 65252 35100 65254
rect 35156 65252 35180 65254
rect 34940 65232 35236 65252
rect 34940 64220 35236 64240
rect 34996 64218 35020 64220
rect 35076 64218 35100 64220
rect 35156 64218 35180 64220
rect 35018 64166 35020 64218
rect 35082 64166 35094 64218
rect 35156 64166 35158 64218
rect 34996 64164 35020 64166
rect 35076 64164 35100 64166
rect 35156 64164 35180 64166
rect 34940 64144 35236 64164
rect 34940 63132 35236 63152
rect 34996 63130 35020 63132
rect 35076 63130 35100 63132
rect 35156 63130 35180 63132
rect 35018 63078 35020 63130
rect 35082 63078 35094 63130
rect 35156 63078 35158 63130
rect 34996 63076 35020 63078
rect 35076 63076 35100 63078
rect 35156 63076 35180 63078
rect 34940 63056 35236 63076
rect 34796 62416 34848 62422
rect 34796 62358 34848 62364
rect 34808 59226 34836 62358
rect 34940 62044 35236 62064
rect 34996 62042 35020 62044
rect 35076 62042 35100 62044
rect 35156 62042 35180 62044
rect 35018 61990 35020 62042
rect 35082 61990 35094 62042
rect 35156 61990 35158 62042
rect 34996 61988 35020 61990
rect 35076 61988 35100 61990
rect 35156 61988 35180 61990
rect 34940 61968 35236 61988
rect 34940 60956 35236 60976
rect 34996 60954 35020 60956
rect 35076 60954 35100 60956
rect 35156 60954 35180 60956
rect 35018 60902 35020 60954
rect 35082 60902 35094 60954
rect 35156 60902 35158 60954
rect 34996 60900 35020 60902
rect 35076 60900 35100 60902
rect 35156 60900 35180 60902
rect 34940 60880 35236 60900
rect 35268 60042 35296 67186
rect 35452 65550 35480 75822
rect 35440 65544 35492 65550
rect 35440 65486 35492 65492
rect 35452 64874 35480 65486
rect 35360 64846 35480 64874
rect 35256 60036 35308 60042
rect 35256 59978 35308 59984
rect 34940 59868 35236 59888
rect 34996 59866 35020 59868
rect 35076 59866 35100 59868
rect 35156 59866 35180 59868
rect 35018 59814 35020 59866
rect 35082 59814 35094 59866
rect 35156 59814 35158 59866
rect 34996 59812 35020 59814
rect 35076 59812 35100 59814
rect 35156 59812 35180 59814
rect 34940 59792 35236 59812
rect 34796 59220 34848 59226
rect 34796 59162 34848 59168
rect 34940 58780 35236 58800
rect 34996 58778 35020 58780
rect 35076 58778 35100 58780
rect 35156 58778 35180 58780
rect 35018 58726 35020 58778
rect 35082 58726 35094 58778
rect 35156 58726 35158 58778
rect 34996 58724 35020 58726
rect 35076 58724 35100 58726
rect 35156 58724 35180 58726
rect 34940 58704 35236 58724
rect 34940 57692 35236 57712
rect 34996 57690 35020 57692
rect 35076 57690 35100 57692
rect 35156 57690 35180 57692
rect 35018 57638 35020 57690
rect 35082 57638 35094 57690
rect 35156 57638 35158 57690
rect 34996 57636 35020 57638
rect 35076 57636 35100 57638
rect 35156 57636 35180 57638
rect 34940 57616 35236 57636
rect 34940 56604 35236 56624
rect 34996 56602 35020 56604
rect 35076 56602 35100 56604
rect 35156 56602 35180 56604
rect 35018 56550 35020 56602
rect 35082 56550 35094 56602
rect 35156 56550 35158 56602
rect 34996 56548 35020 56550
rect 35076 56548 35100 56550
rect 35156 56548 35180 56550
rect 34940 56528 35236 56548
rect 35256 55820 35308 55826
rect 35256 55762 35308 55768
rect 34940 55516 35236 55536
rect 34996 55514 35020 55516
rect 35076 55514 35100 55516
rect 35156 55514 35180 55516
rect 35018 55462 35020 55514
rect 35082 55462 35094 55514
rect 35156 55462 35158 55514
rect 34996 55460 35020 55462
rect 35076 55460 35100 55462
rect 35156 55460 35180 55462
rect 34940 55440 35236 55460
rect 34940 54428 35236 54448
rect 34996 54426 35020 54428
rect 35076 54426 35100 54428
rect 35156 54426 35180 54428
rect 35018 54374 35020 54426
rect 35082 54374 35094 54426
rect 35156 54374 35158 54426
rect 34996 54372 35020 54374
rect 35076 54372 35100 54374
rect 35156 54372 35180 54374
rect 34940 54352 35236 54372
rect 34940 53340 35236 53360
rect 34996 53338 35020 53340
rect 35076 53338 35100 53340
rect 35156 53338 35180 53340
rect 35018 53286 35020 53338
rect 35082 53286 35094 53338
rect 35156 53286 35158 53338
rect 34996 53284 35020 53286
rect 35076 53284 35100 53286
rect 35156 53284 35180 53286
rect 34940 53264 35236 53284
rect 34940 52252 35236 52272
rect 34996 52250 35020 52252
rect 35076 52250 35100 52252
rect 35156 52250 35180 52252
rect 35018 52198 35020 52250
rect 35082 52198 35094 52250
rect 35156 52198 35158 52250
rect 34996 52196 35020 52198
rect 35076 52196 35100 52198
rect 35156 52196 35180 52198
rect 34940 52176 35236 52196
rect 34940 51164 35236 51184
rect 34996 51162 35020 51164
rect 35076 51162 35100 51164
rect 35156 51162 35180 51164
rect 35018 51110 35020 51162
rect 35082 51110 35094 51162
rect 35156 51110 35158 51162
rect 34996 51108 35020 51110
rect 35076 51108 35100 51110
rect 35156 51108 35180 51110
rect 34940 51088 35236 51108
rect 34940 50076 35236 50096
rect 34996 50074 35020 50076
rect 35076 50074 35100 50076
rect 35156 50074 35180 50076
rect 35018 50022 35020 50074
rect 35082 50022 35094 50074
rect 35156 50022 35158 50074
rect 34996 50020 35020 50022
rect 35076 50020 35100 50022
rect 35156 50020 35180 50022
rect 34940 50000 35236 50020
rect 34940 48988 35236 49008
rect 34996 48986 35020 48988
rect 35076 48986 35100 48988
rect 35156 48986 35180 48988
rect 35018 48934 35020 48986
rect 35082 48934 35094 48986
rect 35156 48934 35158 48986
rect 34996 48932 35020 48934
rect 35076 48932 35100 48934
rect 35156 48932 35180 48934
rect 34940 48912 35236 48932
rect 34940 47900 35236 47920
rect 34996 47898 35020 47900
rect 35076 47898 35100 47900
rect 35156 47898 35180 47900
rect 35018 47846 35020 47898
rect 35082 47846 35094 47898
rect 35156 47846 35158 47898
rect 34996 47844 35020 47846
rect 35076 47844 35100 47846
rect 35156 47844 35180 47846
rect 34940 47824 35236 47844
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 35268 43450 35296 55762
rect 35256 43444 35308 43450
rect 35256 43386 35308 43392
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 34612 39976 34664 39982
rect 34612 39918 34664 39924
rect 35256 39976 35308 39982
rect 35256 39918 35308 39924
rect 34704 39908 34756 39914
rect 34704 39850 34756 39856
rect 34716 39506 34744 39850
rect 34796 39840 34848 39846
rect 34796 39782 34848 39788
rect 34704 39500 34756 39506
rect 34704 39442 34756 39448
rect 34520 39092 34572 39098
rect 34520 39034 34572 39040
rect 34520 33856 34572 33862
rect 34520 33798 34572 33804
rect 34532 30326 34560 33798
rect 34808 31210 34836 39782
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 35268 34406 35296 39918
rect 35256 34400 35308 34406
rect 35256 34342 35308 34348
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34796 31204 34848 31210
rect 34796 31146 34848 31152
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34520 30320 34572 30326
rect 34520 30262 34572 30268
rect 34532 26246 34560 30262
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 34796 29640 34848 29646
rect 34796 29582 34848 29588
rect 34716 26450 34744 29582
rect 34808 29034 34836 29582
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34796 29028 34848 29034
rect 34796 28970 34848 28976
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34704 26444 34756 26450
rect 34704 26386 34756 26392
rect 34520 26240 34572 26246
rect 34520 26182 34572 26188
rect 34532 24750 34560 26182
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34520 24744 34572 24750
rect 34520 24686 34572 24692
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 34336 21956 34388 21962
rect 34336 21898 34388 21904
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 34520 18692 34572 18698
rect 34520 18634 34572 18640
rect 34532 18290 34560 18634
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34520 18284 34572 18290
rect 34520 18226 34572 18232
rect 34244 17536 34296 17542
rect 34244 17478 34296 17484
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35268 14958 35296 34342
rect 35360 29170 35388 64846
rect 35808 62824 35860 62830
rect 35808 62766 35860 62772
rect 35440 61192 35492 61198
rect 35440 61134 35492 61140
rect 35452 57050 35480 61134
rect 35440 57044 35492 57050
rect 35440 56986 35492 56992
rect 35348 29164 35400 29170
rect 35348 29106 35400 29112
rect 35452 27554 35480 56986
rect 35820 45554 35848 62766
rect 35900 60240 35952 60246
rect 35900 60182 35952 60188
rect 35912 60042 35940 60182
rect 35900 60036 35952 60042
rect 35900 59978 35952 59984
rect 36096 49162 36124 96426
rect 36360 92200 36412 92206
rect 36360 92142 36412 92148
rect 36372 77178 36400 92142
rect 36360 77172 36412 77178
rect 36360 77114 36412 77120
rect 36372 71126 36400 77114
rect 36360 71120 36412 71126
rect 36360 71062 36412 71068
rect 36544 65748 36596 65754
rect 36544 65690 36596 65696
rect 36556 54738 36584 65690
rect 36636 62144 36688 62150
rect 36636 62086 36688 62092
rect 36544 54732 36596 54738
rect 36544 54674 36596 54680
rect 36648 52562 36676 62086
rect 36268 52556 36320 52562
rect 36268 52498 36320 52504
rect 36636 52556 36688 52562
rect 36636 52498 36688 52504
rect 37004 52556 37056 52562
rect 37004 52498 37056 52504
rect 36084 49156 36136 49162
rect 36084 49098 36136 49104
rect 35728 45526 35848 45554
rect 35728 39302 35756 45526
rect 35808 40112 35860 40118
rect 35808 40054 35860 40060
rect 35716 39296 35768 39302
rect 35716 39238 35768 39244
rect 35532 39092 35584 39098
rect 35532 39034 35584 39040
rect 35360 27526 35480 27554
rect 35360 26858 35388 27526
rect 35348 26852 35400 26858
rect 35348 26794 35400 26800
rect 35360 24274 35388 26794
rect 35544 25430 35572 39034
rect 35728 31754 35756 39238
rect 35820 36242 35848 40054
rect 36176 37392 36228 37398
rect 36176 37334 36228 37340
rect 35808 36236 35860 36242
rect 35808 36178 35860 36184
rect 35636 31726 35756 31754
rect 35532 25424 35584 25430
rect 35532 25366 35584 25372
rect 35440 24608 35492 24614
rect 35440 24550 35492 24556
rect 35348 24268 35400 24274
rect 35348 24210 35400 24216
rect 35452 23050 35480 24550
rect 35440 23044 35492 23050
rect 35440 22986 35492 22992
rect 35636 21894 35664 31726
rect 36084 24812 36136 24818
rect 36084 24754 36136 24760
rect 35808 24744 35860 24750
rect 35808 24686 35860 24692
rect 35716 24608 35768 24614
rect 35716 24550 35768 24556
rect 35624 21888 35676 21894
rect 35624 21830 35676 21836
rect 35728 21690 35756 24550
rect 35348 21684 35400 21690
rect 35348 21626 35400 21632
rect 35716 21684 35768 21690
rect 35716 21626 35768 21632
rect 35256 14952 35308 14958
rect 35256 14894 35308 14900
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 35360 11762 35388 21626
rect 35624 21344 35676 21350
rect 35624 21286 35676 21292
rect 35636 16574 35664 21286
rect 35820 18698 35848 24686
rect 36096 24614 36124 24754
rect 36084 24608 36136 24614
rect 36084 24550 36136 24556
rect 36188 22166 36216 37334
rect 36280 35562 36308 52498
rect 36452 52488 36504 52494
rect 36452 52430 36504 52436
rect 36360 40520 36412 40526
rect 36360 40462 36412 40468
rect 36268 35556 36320 35562
rect 36268 35498 36320 35504
rect 36176 22160 36228 22166
rect 36176 22102 36228 22108
rect 36084 22024 36136 22030
rect 36084 21966 36136 21972
rect 35808 18692 35860 18698
rect 35808 18634 35860 18640
rect 35452 16546 35664 16574
rect 36096 16574 36124 21966
rect 36096 16546 36216 16574
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 35452 5234 35480 16546
rect 35532 10192 35584 10198
rect 35532 10134 35584 10140
rect 35440 5228 35492 5234
rect 35440 5170 35492 5176
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34244 4072 34296 4078
rect 34244 4014 34296 4020
rect 34796 4072 34848 4078
rect 34796 4014 34848 4020
rect 35440 4072 35492 4078
rect 35440 4014 35492 4020
rect 34152 2644 34204 2650
rect 34152 2586 34204 2592
rect 33968 2372 34020 2378
rect 33968 2314 34020 2320
rect 33980 800 34008 2314
rect 34256 800 34284 4014
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34440 800 34468 3538
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 34624 800 34652 2382
rect 34808 800 34836 4014
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35256 2916 35308 2922
rect 35256 2858 35308 2864
rect 35348 2916 35400 2922
rect 35348 2858 35400 2864
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35072 1556 35124 1562
rect 35072 1498 35124 1504
rect 35084 800 35112 1498
rect 35268 800 35296 2858
rect 35360 1562 35388 2858
rect 35348 1556 35400 1562
rect 35348 1498 35400 1504
rect 35452 800 35480 4014
rect 35544 2990 35572 10134
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 35624 3596 35676 3602
rect 35624 3538 35676 3544
rect 35532 2984 35584 2990
rect 35532 2926 35584 2932
rect 35636 800 35664 3538
rect 35808 3120 35860 3126
rect 35808 3062 35860 3068
rect 35820 800 35848 3062
rect 35992 2644 36044 2650
rect 35992 2586 36044 2592
rect 36004 2106 36032 2586
rect 35992 2100 36044 2106
rect 35992 2042 36044 2048
rect 36096 800 36124 4014
rect 36188 2650 36216 16546
rect 36372 10606 36400 40462
rect 36464 13530 36492 52430
rect 37016 51950 37044 52498
rect 37004 51944 37056 51950
rect 37004 51886 37056 51892
rect 36636 51876 36688 51882
rect 36636 51818 36688 51824
rect 36648 48142 36676 51818
rect 36820 50176 36872 50182
rect 36820 50118 36872 50124
rect 36728 49224 36780 49230
rect 36728 49166 36780 49172
rect 36636 48136 36688 48142
rect 36636 48078 36688 48084
rect 36648 45554 36676 48078
rect 36740 47530 36768 49166
rect 36728 47524 36780 47530
rect 36728 47466 36780 47472
rect 36648 45526 36768 45554
rect 36544 41064 36596 41070
rect 36544 41006 36596 41012
rect 36556 40526 36584 41006
rect 36544 40520 36596 40526
rect 36544 40462 36596 40468
rect 36544 30048 36596 30054
rect 36544 29990 36596 29996
rect 36556 29306 36584 29990
rect 36544 29300 36596 29306
rect 36544 29242 36596 29248
rect 36636 24336 36688 24342
rect 36636 24278 36688 24284
rect 36648 24206 36676 24278
rect 36636 24200 36688 24206
rect 36636 24142 36688 24148
rect 36452 13524 36504 13530
rect 36452 13466 36504 13472
rect 36648 10606 36676 24142
rect 36740 10606 36768 45526
rect 36832 16574 36860 50118
rect 36912 47524 36964 47530
rect 36912 47466 36964 47472
rect 36924 22098 36952 47466
rect 37108 47122 37136 96902
rect 37556 76288 37608 76294
rect 37556 76230 37608 76236
rect 37568 57458 37596 76230
rect 37844 63034 37872 97106
rect 38580 96626 38608 99200
rect 39500 97238 39528 99200
rect 40328 97306 40356 99200
rect 40316 97300 40368 97306
rect 40316 97242 40368 97248
rect 39488 97232 39540 97238
rect 39488 97174 39540 97180
rect 40500 97164 40552 97170
rect 40500 97106 40552 97112
rect 39672 96960 39724 96966
rect 39672 96902 39724 96908
rect 38568 96620 38620 96626
rect 38568 96562 38620 96568
rect 38752 96552 38804 96558
rect 38752 96494 38804 96500
rect 38660 96484 38712 96490
rect 38660 96426 38712 96432
rect 38672 75886 38700 96426
rect 38764 94926 38792 96494
rect 38752 94920 38804 94926
rect 38752 94862 38804 94868
rect 38016 75880 38068 75886
rect 38016 75822 38068 75828
rect 38660 75880 38712 75886
rect 38660 75822 38712 75828
rect 37924 69828 37976 69834
rect 37924 69770 37976 69776
rect 37832 63028 37884 63034
rect 37832 62970 37884 62976
rect 37740 59424 37792 59430
rect 37740 59366 37792 59372
rect 37752 59090 37780 59366
rect 37740 59084 37792 59090
rect 37740 59026 37792 59032
rect 37556 57452 37608 57458
rect 37556 57394 37608 57400
rect 37464 56908 37516 56914
rect 37464 56850 37516 56856
rect 37476 56370 37504 56850
rect 37464 56364 37516 56370
rect 37464 56306 37516 56312
rect 37832 54528 37884 54534
rect 37832 54470 37884 54476
rect 37372 52488 37424 52494
rect 37372 52430 37424 52436
rect 37096 47116 37148 47122
rect 37096 47058 37148 47064
rect 36912 22092 36964 22098
rect 36912 22034 36964 22040
rect 36832 16546 36952 16574
rect 36360 10600 36412 10606
rect 36360 10542 36412 10548
rect 36636 10600 36688 10606
rect 36636 10542 36688 10548
rect 36728 10600 36780 10606
rect 36728 10542 36780 10548
rect 36636 4072 36688 4078
rect 36636 4014 36688 4020
rect 36268 2984 36320 2990
rect 36268 2926 36320 2932
rect 36176 2644 36228 2650
rect 36176 2586 36228 2592
rect 36280 800 36308 2926
rect 36452 2304 36504 2310
rect 36452 2246 36504 2252
rect 36464 800 36492 2246
rect 36648 800 36676 4014
rect 36820 3596 36872 3602
rect 36820 3538 36872 3544
rect 36832 800 36860 3538
rect 36924 2650 36952 16546
rect 37188 13524 37240 13530
rect 37188 13466 37240 13472
rect 37200 12986 37228 13466
rect 37188 12980 37240 12986
rect 37188 12922 37240 12928
rect 37384 11218 37412 52430
rect 37844 52426 37872 54470
rect 37832 52420 37884 52426
rect 37832 52362 37884 52368
rect 37844 51814 37872 52362
rect 37832 51808 37884 51814
rect 37832 51750 37884 51756
rect 37832 48000 37884 48006
rect 37832 47942 37884 47948
rect 37556 43784 37608 43790
rect 37556 43726 37608 43732
rect 37568 11626 37596 43726
rect 37844 16182 37872 47942
rect 37832 16176 37884 16182
rect 37832 16118 37884 16124
rect 37740 14272 37792 14278
rect 37740 14214 37792 14220
rect 37752 14074 37780 14214
rect 37740 14068 37792 14074
rect 37740 14010 37792 14016
rect 37556 11620 37608 11626
rect 37556 11562 37608 11568
rect 37372 11212 37424 11218
rect 37372 11154 37424 11160
rect 37280 4684 37332 4690
rect 37280 4626 37332 4632
rect 37096 2848 37148 2854
rect 37096 2790 37148 2796
rect 36912 2644 36964 2650
rect 36912 2586 36964 2592
rect 37108 800 37136 2790
rect 37292 800 37320 4626
rect 37832 4072 37884 4078
rect 37832 4014 37884 4020
rect 37464 3596 37516 3602
rect 37464 3538 37516 3544
rect 37476 800 37504 3538
rect 37648 2916 37700 2922
rect 37648 2858 37700 2864
rect 37660 800 37688 2858
rect 37844 800 37872 4014
rect 37936 2582 37964 69770
rect 38028 52562 38056 75822
rect 38200 65680 38252 65686
rect 38200 65622 38252 65628
rect 38108 56364 38160 56370
rect 38108 56306 38160 56312
rect 38016 52556 38068 52562
rect 38016 52498 38068 52504
rect 38028 47190 38056 52498
rect 38016 47184 38068 47190
rect 38016 47126 38068 47132
rect 38028 11082 38056 47126
rect 38120 38418 38148 56306
rect 38212 49230 38240 65622
rect 38292 59696 38344 59702
rect 38292 59638 38344 59644
rect 38304 59566 38332 59638
rect 38292 59560 38344 59566
rect 38292 59502 38344 59508
rect 38304 53106 38332 59502
rect 38292 53100 38344 53106
rect 38292 53042 38344 53048
rect 38200 49224 38252 49230
rect 38200 49166 38252 49172
rect 38660 43376 38712 43382
rect 38660 43318 38712 43324
rect 38672 42906 38700 43318
rect 38660 42900 38712 42906
rect 38660 42842 38712 42848
rect 38108 38412 38160 38418
rect 38108 38354 38160 38360
rect 38108 18692 38160 18698
rect 38108 18634 38160 18640
rect 38120 18086 38148 18634
rect 38108 18080 38160 18086
rect 38108 18022 38160 18028
rect 38120 12306 38148 18022
rect 38108 12300 38160 12306
rect 38108 12242 38160 12248
rect 38016 11076 38068 11082
rect 38016 11018 38068 11024
rect 38200 10464 38252 10470
rect 38200 10406 38252 10412
rect 38108 3596 38160 3602
rect 38108 3538 38160 3544
rect 37924 2576 37976 2582
rect 37924 2518 37976 2524
rect 38120 800 38148 3538
rect 38212 3194 38240 10406
rect 38764 6730 38792 94862
rect 39396 90432 39448 90438
rect 39396 90374 39448 90380
rect 38844 73840 38896 73846
rect 38844 73782 38896 73788
rect 38856 59566 38884 73782
rect 38844 59560 38896 59566
rect 38844 59502 38896 59508
rect 39028 59492 39080 59498
rect 39028 59434 39080 59440
rect 39040 59226 39068 59434
rect 39028 59220 39080 59226
rect 39028 59162 39080 59168
rect 39304 52352 39356 52358
rect 39304 52294 39356 52300
rect 38844 43716 38896 43722
rect 38844 43658 38896 43664
rect 38856 43450 38884 43658
rect 38844 43444 38896 43450
rect 38844 43386 38896 43392
rect 39316 16574 39344 52294
rect 39408 25498 39436 90374
rect 39488 82340 39540 82346
rect 39488 82282 39540 82288
rect 39396 25492 39448 25498
rect 39396 25434 39448 25440
rect 39500 18834 39528 82282
rect 39580 73908 39632 73914
rect 39580 73850 39632 73856
rect 39488 18828 39540 18834
rect 39488 18770 39540 18776
rect 39316 16546 39436 16574
rect 38752 6724 38804 6730
rect 38752 6666 38804 6672
rect 38764 6322 38792 6666
rect 38752 6316 38804 6322
rect 38752 6258 38804 6264
rect 39120 4684 39172 4690
rect 39120 4626 39172 4632
rect 38476 4072 38528 4078
rect 38476 4014 38528 4020
rect 38200 3188 38252 3194
rect 38200 3130 38252 3136
rect 38212 2990 38240 3130
rect 38200 2984 38252 2990
rect 38200 2926 38252 2932
rect 38292 2440 38344 2446
rect 38292 2382 38344 2388
rect 38304 800 38332 2382
rect 38488 800 38516 4014
rect 38936 3120 38988 3126
rect 38936 3062 38988 3068
rect 38660 2984 38712 2990
rect 38660 2926 38712 2932
rect 38672 800 38700 2926
rect 38752 2848 38804 2854
rect 38752 2790 38804 2796
rect 38764 2514 38792 2790
rect 38948 2582 38976 3062
rect 38936 2576 38988 2582
rect 38936 2518 38988 2524
rect 38752 2508 38804 2514
rect 38752 2450 38804 2456
rect 38844 2372 38896 2378
rect 38844 2314 38896 2320
rect 38856 800 38884 2314
rect 39132 800 39160 4626
rect 39304 3596 39356 3602
rect 39304 3538 39356 3544
rect 39316 800 39344 3538
rect 39408 2650 39436 16546
rect 39592 13258 39620 73850
rect 39684 64870 39712 96902
rect 40512 93770 40540 97106
rect 40684 96688 40736 96694
rect 40684 96630 40736 96636
rect 40500 93764 40552 93770
rect 40500 93706 40552 93712
rect 40512 93158 40540 93706
rect 40500 93152 40552 93158
rect 40500 93094 40552 93100
rect 39856 84720 39908 84726
rect 39856 84662 39908 84668
rect 39764 68128 39816 68134
rect 39764 68070 39816 68076
rect 39672 64864 39724 64870
rect 39672 64806 39724 64812
rect 39672 51264 39724 51270
rect 39672 51206 39724 51212
rect 39580 13252 39632 13258
rect 39580 13194 39632 13200
rect 39684 9178 39712 51206
rect 39776 43994 39804 68070
rect 39764 43988 39816 43994
rect 39764 43930 39816 43936
rect 39764 42220 39816 42226
rect 39764 42162 39816 42168
rect 39776 40118 39804 42162
rect 39764 40112 39816 40118
rect 39764 40054 39816 40060
rect 39764 36168 39816 36174
rect 39764 36110 39816 36116
rect 39776 13870 39804 36110
rect 39868 35154 39896 84662
rect 39948 73840 40000 73846
rect 39948 73782 40000 73788
rect 39960 73302 39988 73782
rect 39948 73296 40000 73302
rect 39948 73238 40000 73244
rect 39948 62212 40000 62218
rect 39948 62154 40000 62160
rect 39856 35148 39908 35154
rect 39856 35090 39908 35096
rect 39960 34134 39988 62154
rect 40316 45348 40368 45354
rect 40316 45290 40368 45296
rect 40328 44470 40356 45290
rect 40316 44464 40368 44470
rect 40316 44406 40368 44412
rect 40040 43716 40092 43722
rect 40040 43658 40092 43664
rect 40052 43382 40080 43658
rect 40040 43376 40092 43382
rect 40040 43318 40092 43324
rect 40224 43240 40276 43246
rect 40224 43182 40276 43188
rect 40040 39092 40092 39098
rect 40040 39034 40092 39040
rect 40052 35290 40080 39034
rect 40040 35284 40092 35290
rect 40040 35226 40092 35232
rect 39948 34128 40000 34134
rect 39948 34070 40000 34076
rect 39948 31816 40000 31822
rect 39948 31758 40000 31764
rect 39856 17672 39908 17678
rect 39856 17614 39908 17620
rect 39764 13864 39816 13870
rect 39764 13806 39816 13812
rect 39672 9172 39724 9178
rect 39672 9114 39724 9120
rect 39776 7750 39804 13806
rect 39764 7744 39816 7750
rect 39764 7686 39816 7692
rect 39672 4684 39724 4690
rect 39672 4626 39724 4632
rect 39396 2644 39448 2650
rect 39396 2586 39448 2592
rect 39488 1216 39540 1222
rect 39488 1158 39540 1164
rect 39500 800 39528 1158
rect 39684 800 39712 4626
rect 39776 3670 39804 7686
rect 39764 3664 39816 3670
rect 39764 3606 39816 3612
rect 39868 2582 39896 17614
rect 39960 10198 39988 31758
rect 40236 31754 40264 43182
rect 40144 31726 40264 31754
rect 40040 29844 40092 29850
rect 40040 29786 40092 29792
rect 40052 28966 40080 29786
rect 40144 29238 40172 31726
rect 40132 29232 40184 29238
rect 40132 29174 40184 29180
rect 40040 28960 40092 28966
rect 40040 28902 40092 28908
rect 40144 28694 40172 29174
rect 40132 28688 40184 28694
rect 40132 28630 40184 28636
rect 40040 26580 40092 26586
rect 40040 26522 40092 26528
rect 40052 23662 40080 26522
rect 40328 23730 40356 44406
rect 40500 43172 40552 43178
rect 40500 43114 40552 43120
rect 40512 29850 40540 43114
rect 40592 39840 40644 39846
rect 40592 39782 40644 39788
rect 40604 39030 40632 39782
rect 40592 39024 40644 39030
rect 40592 38966 40644 38972
rect 40500 29844 40552 29850
rect 40500 29786 40552 29792
rect 40316 23724 40368 23730
rect 40316 23666 40368 23672
rect 40040 23656 40092 23662
rect 40040 23598 40092 23604
rect 40040 16108 40092 16114
rect 40040 16050 40092 16056
rect 39948 10192 40000 10198
rect 39948 10134 40000 10140
rect 39948 4072 40000 4078
rect 39948 4014 40000 4020
rect 39856 2576 39908 2582
rect 39856 2518 39908 2524
rect 39960 800 39988 4014
rect 40052 2650 40080 16050
rect 40696 10538 40724 96630
rect 41248 96626 41276 99200
rect 42076 97238 42104 99200
rect 42996 97306 43024 99200
rect 42984 97300 43036 97306
rect 42984 97242 43036 97248
rect 42064 97232 42116 97238
rect 42064 97174 42116 97180
rect 43076 97164 43128 97170
rect 43076 97106 43128 97112
rect 42064 97096 42116 97102
rect 42064 97038 42116 97044
rect 41236 96620 41288 96626
rect 41236 96562 41288 96568
rect 41328 96484 41380 96490
rect 41328 96426 41380 96432
rect 41052 90228 41104 90234
rect 41052 90170 41104 90176
rect 41064 88058 41092 90170
rect 41052 88052 41104 88058
rect 41052 87994 41104 88000
rect 40776 80096 40828 80102
rect 40776 80038 40828 80044
rect 40788 63986 40816 80038
rect 40776 63980 40828 63986
rect 40776 63922 40828 63928
rect 40776 39976 40828 39982
rect 40776 39918 40828 39924
rect 40788 39642 40816 39918
rect 41064 39914 41092 87994
rect 41340 80102 41368 96426
rect 41880 94376 41932 94382
rect 41880 94318 41932 94324
rect 41892 82346 41920 94318
rect 42076 84794 42104 97038
rect 42248 96960 42300 96966
rect 42248 96902 42300 96908
rect 42260 95062 42288 96902
rect 42248 95056 42300 95062
rect 42248 94998 42300 95004
rect 42064 84788 42116 84794
rect 42064 84730 42116 84736
rect 41880 82340 41932 82346
rect 41880 82282 41932 82288
rect 41328 80096 41380 80102
rect 41328 80038 41380 80044
rect 42892 79824 42944 79830
rect 42892 79766 42944 79772
rect 42616 79756 42668 79762
rect 42616 79698 42668 79704
rect 42628 79665 42656 79698
rect 42614 79656 42670 79665
rect 42614 79591 42670 79600
rect 42708 61600 42760 61606
rect 42708 61542 42760 61548
rect 42720 61402 42748 61542
rect 41604 61396 41656 61402
rect 41604 61338 41656 61344
rect 42708 61396 42760 61402
rect 42708 61338 42760 61344
rect 41144 61260 41196 61266
rect 41144 61202 41196 61208
rect 41420 61260 41472 61266
rect 41420 61202 41472 61208
rect 41052 39908 41104 39914
rect 41052 39850 41104 39856
rect 40776 39636 40828 39642
rect 40776 39578 40828 39584
rect 40868 36304 40920 36310
rect 40868 36246 40920 36252
rect 40776 33108 40828 33114
rect 40776 33050 40828 33056
rect 40788 31890 40816 33050
rect 40776 31884 40828 31890
rect 40776 31826 40828 31832
rect 40788 12714 40816 31826
rect 40776 12708 40828 12714
rect 40776 12650 40828 12656
rect 40684 10532 40736 10538
rect 40684 10474 40736 10480
rect 40224 10260 40276 10266
rect 40224 10202 40276 10208
rect 40236 2990 40264 10202
rect 40788 9042 40816 12650
rect 40880 9382 40908 36246
rect 40960 33856 41012 33862
rect 40960 33798 41012 33804
rect 40972 24138 41000 33798
rect 41064 30054 41092 39850
rect 41156 39098 41184 61202
rect 41236 39908 41288 39914
rect 41236 39850 41288 39856
rect 41248 39302 41276 39850
rect 41236 39296 41288 39302
rect 41236 39238 41288 39244
rect 41144 39092 41196 39098
rect 41144 39034 41196 39040
rect 41328 38344 41380 38350
rect 41328 38286 41380 38292
rect 41340 36310 41368 38286
rect 41328 36304 41380 36310
rect 41328 36246 41380 36252
rect 41236 30184 41288 30190
rect 41236 30126 41288 30132
rect 41052 30048 41104 30054
rect 41052 29990 41104 29996
rect 41248 29170 41276 30126
rect 41236 29164 41288 29170
rect 41236 29106 41288 29112
rect 40960 24132 41012 24138
rect 40960 24074 41012 24080
rect 41052 12912 41104 12918
rect 41052 12854 41104 12860
rect 41064 12646 41092 12854
rect 41144 12844 41196 12850
rect 41144 12786 41196 12792
rect 41052 12640 41104 12646
rect 41052 12582 41104 12588
rect 40868 9376 40920 9382
rect 40868 9318 40920 9324
rect 40776 9036 40828 9042
rect 40776 8978 40828 8984
rect 41064 7478 41092 12582
rect 41052 7472 41104 7478
rect 41052 7414 41104 7420
rect 41156 4758 41184 12786
rect 41248 11762 41276 29106
rect 41432 26994 41460 61202
rect 41616 39982 41644 61338
rect 42904 61266 42932 79766
rect 41696 61260 41748 61266
rect 41696 61202 41748 61208
rect 42892 61260 42944 61266
rect 42892 61202 42944 61208
rect 41708 51270 41736 61202
rect 41880 61192 41932 61198
rect 41880 61134 41932 61140
rect 41892 56234 41920 61134
rect 43088 59090 43116 97106
rect 43444 97096 43496 97102
rect 43444 97038 43496 97044
rect 43456 96694 43484 97038
rect 43444 96688 43496 96694
rect 43444 96630 43496 96636
rect 43824 96626 43852 99200
rect 44744 97238 44772 99200
rect 44732 97232 44784 97238
rect 44732 97174 44784 97180
rect 45468 97164 45520 97170
rect 45468 97106 45520 97112
rect 44916 96960 44968 96966
rect 44916 96902 44968 96908
rect 43812 96620 43864 96626
rect 43812 96562 43864 96568
rect 44824 93900 44876 93906
rect 44824 93842 44876 93848
rect 44456 90024 44508 90030
rect 44456 89966 44508 89972
rect 44180 89956 44232 89962
rect 44180 89898 44232 89904
rect 43812 88528 43864 88534
rect 43812 88470 43864 88476
rect 43536 86284 43588 86290
rect 43536 86226 43588 86232
rect 43168 79756 43220 79762
rect 43168 79698 43220 79704
rect 43076 59084 43128 59090
rect 43076 59026 43128 59032
rect 41880 56228 41932 56234
rect 41880 56170 41932 56176
rect 42708 55344 42760 55350
rect 42708 55286 42760 55292
rect 42720 52630 42748 55286
rect 42708 52624 42760 52630
rect 42708 52566 42760 52572
rect 42156 52556 42208 52562
rect 42156 52498 42208 52504
rect 41880 51944 41932 51950
rect 41880 51886 41932 51892
rect 41696 51264 41748 51270
rect 41696 51206 41748 51212
rect 41604 39976 41656 39982
rect 41604 39918 41656 39924
rect 41616 34474 41644 39918
rect 41604 34468 41656 34474
rect 41604 34410 41656 34416
rect 41420 26988 41472 26994
rect 41420 26930 41472 26936
rect 41432 24410 41460 26930
rect 41708 26790 41736 51206
rect 41892 45490 41920 51886
rect 42168 51882 42196 52498
rect 42156 51876 42208 51882
rect 42156 51818 42208 51824
rect 43076 51808 43128 51814
rect 43076 51750 43128 51756
rect 42340 50720 42392 50726
rect 42340 50662 42392 50668
rect 42352 49230 42380 50662
rect 42340 49224 42392 49230
rect 42340 49166 42392 49172
rect 42352 48210 42380 49166
rect 42340 48204 42392 48210
rect 42340 48146 42392 48152
rect 41880 45484 41932 45490
rect 41880 45426 41932 45432
rect 41892 44470 41920 45426
rect 41880 44464 41932 44470
rect 41880 44406 41932 44412
rect 42892 42900 42944 42906
rect 42892 42842 42944 42848
rect 42800 42152 42852 42158
rect 42800 42094 42852 42100
rect 42812 41750 42840 42094
rect 42800 41744 42852 41750
rect 42800 41686 42852 41692
rect 42524 40996 42576 41002
rect 42524 40938 42576 40944
rect 42064 39636 42116 39642
rect 42064 39578 42116 39584
rect 42076 36242 42104 39578
rect 42536 38418 42564 40938
rect 42904 38418 42932 42842
rect 42984 41744 43036 41750
rect 42984 41686 43036 41692
rect 42524 38412 42576 38418
rect 42524 38354 42576 38360
rect 42892 38412 42944 38418
rect 42892 38354 42944 38360
rect 42536 38282 42564 38354
rect 42996 38350 43024 41686
rect 43088 38418 43116 51750
rect 43076 38412 43128 38418
rect 43076 38354 43128 38360
rect 42984 38344 43036 38350
rect 42984 38286 43036 38292
rect 42524 38276 42576 38282
rect 42524 38218 42576 38224
rect 42892 37936 42944 37942
rect 42892 37878 42944 37884
rect 42064 36236 42116 36242
rect 42064 36178 42116 36184
rect 41788 32224 41840 32230
rect 41788 32166 41840 32172
rect 41696 26784 41748 26790
rect 41696 26726 41748 26732
rect 41420 24404 41472 24410
rect 41420 24346 41472 24352
rect 41708 23798 41736 26726
rect 41696 23792 41748 23798
rect 41696 23734 41748 23740
rect 41420 13252 41472 13258
rect 41420 13194 41472 13200
rect 41236 11756 41288 11762
rect 41236 11698 41288 11704
rect 41144 4752 41196 4758
rect 41144 4694 41196 4700
rect 40316 4072 40368 4078
rect 40316 4014 40368 4020
rect 40960 4072 41012 4078
rect 40960 4014 41012 4020
rect 40224 2984 40276 2990
rect 40224 2926 40276 2932
rect 40132 2848 40184 2854
rect 40132 2790 40184 2796
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 40144 800 40172 2790
rect 40328 800 40356 4014
rect 40500 3596 40552 3602
rect 40500 3538 40552 3544
rect 40512 800 40540 3538
rect 40684 2372 40736 2378
rect 40684 2314 40736 2320
rect 40696 800 40724 2314
rect 40972 800 41000 4014
rect 41328 2916 41380 2922
rect 41328 2858 41380 2864
rect 41144 2848 41196 2854
rect 41144 2790 41196 2796
rect 41156 800 41184 2790
rect 41340 800 41368 2858
rect 41432 2650 41460 13194
rect 41604 12912 41656 12918
rect 41604 12854 41656 12860
rect 41616 12782 41644 12854
rect 41604 12776 41656 12782
rect 41604 12718 41656 12724
rect 41800 6914 41828 32166
rect 42076 27538 42104 36178
rect 42800 35216 42852 35222
rect 42800 35158 42852 35164
rect 42812 27538 42840 35158
rect 42904 27538 42932 37878
rect 43076 31816 43128 31822
rect 43076 31758 43128 31764
rect 43088 30326 43116 31758
rect 43076 30320 43128 30326
rect 43076 30262 43128 30268
rect 42064 27532 42116 27538
rect 42064 27474 42116 27480
rect 42800 27532 42852 27538
rect 42800 27474 42852 27480
rect 42892 27532 42944 27538
rect 42892 27474 42944 27480
rect 42708 27464 42760 27470
rect 42984 27464 43036 27470
rect 42760 27412 42840 27418
rect 42708 27406 42840 27412
rect 42984 27406 43036 27412
rect 42720 27390 42840 27406
rect 42616 27328 42668 27334
rect 42616 27270 42668 27276
rect 42628 27062 42656 27270
rect 42616 27056 42668 27062
rect 42616 26998 42668 27004
rect 42812 26314 42840 27390
rect 42800 26308 42852 26314
rect 42800 26250 42852 26256
rect 42248 25832 42300 25838
rect 42248 25774 42300 25780
rect 42260 23798 42288 25774
rect 42248 23792 42300 23798
rect 42248 23734 42300 23740
rect 42800 18760 42852 18766
rect 42800 18702 42852 18708
rect 42812 18086 42840 18702
rect 42800 18080 42852 18086
rect 42800 18022 42852 18028
rect 42432 16244 42484 16250
rect 42432 16186 42484 16192
rect 41616 6886 41828 6914
rect 41512 4072 41564 4078
rect 41512 4014 41564 4020
rect 41420 2644 41472 2650
rect 41420 2586 41472 2592
rect 41524 800 41552 4014
rect 41616 2990 41644 6886
rect 41696 3596 41748 3602
rect 41696 3538 41748 3544
rect 42340 3596 42392 3602
rect 42340 3538 42392 3544
rect 41604 2984 41656 2990
rect 41604 2926 41656 2932
rect 41708 800 41736 3538
rect 42156 3528 42208 3534
rect 42156 3470 42208 3476
rect 41972 2304 42024 2310
rect 41972 2246 42024 2252
rect 41984 800 42012 2246
rect 42168 800 42196 3470
rect 42352 800 42380 3538
rect 42444 2582 42472 16186
rect 42812 11218 42840 18022
rect 42996 14482 43024 27406
rect 43076 22024 43128 22030
rect 43074 21992 43076 22001
rect 43128 21992 43130 22001
rect 43074 21927 43130 21936
rect 43076 19712 43128 19718
rect 43076 19654 43128 19660
rect 43088 19514 43116 19654
rect 43076 19508 43128 19514
rect 43076 19450 43128 19456
rect 43180 19310 43208 79698
rect 43442 79656 43498 79665
rect 43442 79591 43498 79600
rect 43456 79558 43484 79591
rect 43444 79552 43496 79558
rect 43444 79494 43496 79500
rect 43444 75404 43496 75410
rect 43444 75346 43496 75352
rect 43456 54670 43484 75346
rect 43548 69970 43576 86226
rect 43824 76974 43852 88470
rect 43812 76968 43864 76974
rect 43812 76910 43864 76916
rect 43824 73166 43852 76910
rect 44088 75880 44140 75886
rect 44088 75822 44140 75828
rect 44100 74458 44128 75822
rect 44192 74662 44220 89898
rect 44468 87446 44496 89966
rect 44456 87440 44508 87446
rect 44456 87382 44508 87388
rect 44180 74656 44232 74662
rect 44180 74598 44232 74604
rect 44088 74452 44140 74458
rect 44088 74394 44140 74400
rect 44100 73642 44128 74394
rect 44088 73636 44140 73642
rect 44088 73578 44140 73584
rect 43812 73160 43864 73166
rect 43812 73102 43864 73108
rect 43536 69964 43588 69970
rect 43536 69906 43588 69912
rect 43548 55146 43576 69906
rect 44272 65408 44324 65414
rect 44272 65350 44324 65356
rect 44284 60314 44312 65350
rect 44548 61668 44600 61674
rect 44548 61610 44600 61616
rect 44560 61334 44588 61610
rect 44548 61328 44600 61334
rect 44548 61270 44600 61276
rect 44272 60308 44324 60314
rect 44272 60250 44324 60256
rect 44272 55276 44324 55282
rect 44272 55218 44324 55224
rect 43628 55208 43680 55214
rect 43628 55150 43680 55156
rect 44180 55208 44232 55214
rect 44180 55150 44232 55156
rect 43536 55140 43588 55146
rect 43536 55082 43588 55088
rect 43444 54664 43496 54670
rect 43444 54606 43496 54612
rect 43352 49700 43404 49706
rect 43352 49642 43404 49648
rect 43364 49162 43392 49642
rect 43352 49156 43404 49162
rect 43352 49098 43404 49104
rect 43260 46572 43312 46578
rect 43260 46514 43312 46520
rect 43272 38554 43300 46514
rect 43548 38826 43576 55082
rect 43536 38820 43588 38826
rect 43536 38762 43588 38768
rect 43260 38548 43312 38554
rect 43260 38490 43312 38496
rect 43352 38548 43404 38554
rect 43352 38490 43404 38496
rect 43364 37942 43392 38490
rect 43352 37936 43404 37942
rect 43352 37878 43404 37884
rect 43548 34610 43576 38762
rect 43536 34604 43588 34610
rect 43536 34546 43588 34552
rect 43536 32428 43588 32434
rect 43536 32370 43588 32376
rect 43352 31816 43404 31822
rect 43352 31758 43404 31764
rect 43260 26308 43312 26314
rect 43260 26250 43312 26256
rect 43168 19304 43220 19310
rect 43168 19246 43220 19252
rect 42984 14476 43036 14482
rect 42984 14418 43036 14424
rect 43272 13326 43300 26250
rect 43364 24886 43392 31758
rect 43548 27470 43576 32370
rect 43536 27464 43588 27470
rect 43536 27406 43588 27412
rect 43352 24880 43404 24886
rect 43352 24822 43404 24828
rect 43640 20262 43668 55150
rect 43720 49088 43772 49094
rect 43720 49030 43772 49036
rect 43732 30410 43760 49030
rect 43812 40112 43864 40118
rect 43812 40054 43864 40060
rect 43824 37738 43852 40054
rect 43812 37732 43864 37738
rect 43812 37674 43864 37680
rect 43824 30546 43852 37674
rect 44192 34202 44220 55150
rect 44284 45554 44312 55218
rect 44456 55208 44508 55214
rect 44456 55150 44508 55156
rect 44468 54874 44496 55150
rect 44456 54868 44508 54874
rect 44456 54810 44508 54816
rect 44284 45526 44404 45554
rect 44272 45280 44324 45286
rect 44272 45222 44324 45228
rect 44284 44266 44312 45222
rect 44272 44260 44324 44266
rect 44272 44202 44324 44208
rect 44376 44146 44404 45526
rect 44284 44118 44404 44146
rect 44284 41274 44312 44118
rect 44364 42016 44416 42022
rect 44364 41958 44416 41964
rect 44272 41268 44324 41274
rect 44272 41210 44324 41216
rect 44284 39574 44312 41210
rect 44272 39568 44324 39574
rect 44272 39510 44324 39516
rect 44180 34196 44232 34202
rect 44180 34138 44232 34144
rect 44376 31754 44404 41958
rect 44560 33998 44588 61270
rect 44640 56228 44692 56234
rect 44640 56170 44692 56176
rect 44652 41206 44680 56170
rect 44732 43240 44784 43246
rect 44732 43182 44784 43188
rect 44640 41200 44692 41206
rect 44640 41142 44692 41148
rect 44548 33992 44600 33998
rect 44548 33934 44600 33940
rect 44560 31754 44588 33934
rect 44376 31726 44496 31754
rect 44560 31726 44680 31754
rect 43824 30518 44036 30546
rect 43732 30382 43852 30410
rect 43720 30320 43772 30326
rect 43720 30262 43772 30268
rect 43732 29102 43760 30262
rect 43720 29096 43772 29102
rect 43720 29038 43772 29044
rect 43720 28008 43772 28014
rect 43720 27950 43772 27956
rect 43732 27674 43760 27950
rect 43720 27668 43772 27674
rect 43720 27610 43772 27616
rect 43732 23050 43760 27610
rect 43824 26042 43852 30382
rect 44008 28014 44036 30518
rect 44180 28212 44232 28218
rect 44180 28154 44232 28160
rect 44192 28014 44220 28154
rect 43996 28008 44048 28014
rect 43996 27950 44048 27956
rect 44180 28008 44232 28014
rect 44180 27950 44232 27956
rect 44272 27940 44324 27946
rect 44272 27882 44324 27888
rect 43812 26036 43864 26042
rect 43812 25978 43864 25984
rect 44088 26036 44140 26042
rect 44088 25978 44140 25984
rect 44100 25498 44128 25978
rect 44284 25974 44312 27882
rect 44468 26042 44496 31726
rect 44652 28422 44680 31726
rect 44640 28416 44692 28422
rect 44640 28358 44692 28364
rect 44548 28008 44600 28014
rect 44548 27950 44600 27956
rect 44560 27878 44588 27950
rect 44548 27872 44600 27878
rect 44548 27814 44600 27820
rect 44456 26036 44508 26042
rect 44456 25978 44508 25984
rect 44272 25968 44324 25974
rect 44272 25910 44324 25916
rect 44088 25492 44140 25498
rect 44088 25434 44140 25440
rect 44364 25288 44416 25294
rect 44364 25230 44416 25236
rect 43720 23044 43772 23050
rect 43720 22986 43772 22992
rect 43720 21684 43772 21690
rect 43720 21626 43772 21632
rect 43628 20256 43680 20262
rect 43628 20198 43680 20204
rect 43260 13320 43312 13326
rect 43260 13262 43312 13268
rect 42800 11212 42852 11218
rect 42800 11154 42852 11160
rect 43352 7268 43404 7274
rect 43352 7210 43404 7216
rect 43364 4826 43392 7210
rect 43640 6914 43668 20198
rect 43456 6886 43668 6914
rect 43456 5098 43484 6886
rect 43444 5092 43496 5098
rect 43444 5034 43496 5040
rect 43352 4820 43404 4826
rect 43352 4762 43404 4768
rect 42708 4072 42760 4078
rect 42708 4014 42760 4020
rect 42432 2576 42484 2582
rect 42432 2518 42484 2524
rect 42524 2440 42576 2446
rect 42524 2382 42576 2388
rect 42536 800 42564 2382
rect 42720 800 42748 4014
rect 43352 4004 43404 4010
rect 43352 3946 43404 3952
rect 42984 3596 43036 3602
rect 42984 3538 43036 3544
rect 42996 800 43024 3538
rect 43168 2916 43220 2922
rect 43168 2858 43220 2864
rect 43076 2440 43128 2446
rect 43076 2382 43128 2388
rect 43088 1222 43116 2382
rect 43076 1216 43128 1222
rect 43076 1158 43128 1164
rect 43180 800 43208 2858
rect 43364 800 43392 3946
rect 43536 3052 43588 3058
rect 43536 2994 43588 3000
rect 43548 800 43576 2994
rect 43732 2990 43760 21626
rect 43812 17536 43864 17542
rect 43812 17478 43864 17484
rect 43720 2984 43772 2990
rect 43720 2926 43772 2932
rect 43824 2582 43852 17478
rect 44376 14482 44404 25230
rect 44560 23254 44588 27814
rect 44548 23248 44600 23254
rect 44548 23190 44600 23196
rect 44454 19544 44510 19553
rect 44454 19479 44510 19488
rect 44468 19378 44496 19479
rect 44548 19440 44600 19446
rect 44546 19408 44548 19417
rect 44600 19408 44602 19417
rect 44456 19372 44508 19378
rect 44546 19343 44602 19352
rect 44456 19314 44508 19320
rect 44652 19310 44680 28358
rect 44640 19304 44692 19310
rect 44640 19246 44692 19252
rect 44456 17672 44508 17678
rect 44456 17614 44508 17620
rect 44468 16726 44496 17614
rect 44640 17196 44692 17202
rect 44640 17138 44692 17144
rect 44652 16726 44680 17138
rect 44744 16794 44772 43182
rect 44836 40118 44864 93842
rect 44928 89894 44956 96902
rect 45480 93906 45508 97106
rect 45572 96966 45600 99200
rect 45560 96960 45612 96966
rect 45560 96902 45612 96908
rect 46112 96552 46164 96558
rect 46112 96494 46164 96500
rect 45468 93900 45520 93906
rect 45468 93842 45520 93848
rect 44916 89888 44968 89894
rect 44916 89830 44968 89836
rect 45100 87440 45152 87446
rect 45100 87382 45152 87388
rect 44916 86216 44968 86222
rect 44916 86158 44968 86164
rect 44928 54058 44956 86158
rect 45008 85604 45060 85610
rect 45008 85546 45060 85552
rect 44916 54052 44968 54058
rect 44916 53994 44968 54000
rect 44824 40112 44876 40118
rect 44824 40054 44876 40060
rect 44824 39976 44876 39982
rect 44824 39918 44876 39924
rect 44836 39846 44864 39918
rect 44824 39840 44876 39846
rect 44824 39782 44876 39788
rect 44732 16788 44784 16794
rect 44732 16730 44784 16736
rect 44456 16720 44508 16726
rect 44456 16662 44508 16668
rect 44640 16720 44692 16726
rect 44640 16662 44692 16668
rect 44836 14958 44864 39782
rect 44916 39500 44968 39506
rect 44916 39442 44968 39448
rect 44824 14952 44876 14958
rect 44824 14894 44876 14900
rect 44364 14476 44416 14482
rect 44364 14418 44416 14424
rect 44732 14476 44784 14482
rect 44732 14418 44784 14424
rect 44824 14476 44876 14482
rect 44928 14464 44956 39442
rect 45020 32230 45048 85546
rect 45112 45554 45140 87382
rect 45468 85332 45520 85338
rect 45468 85274 45520 85280
rect 45192 85128 45244 85134
rect 45192 85070 45244 85076
rect 45204 53990 45232 85070
rect 45284 73840 45336 73846
rect 45284 73782 45336 73788
rect 45192 53984 45244 53990
rect 45192 53926 45244 53932
rect 45296 48346 45324 73782
rect 45480 65414 45508 85274
rect 45560 68400 45612 68406
rect 45560 68342 45612 68348
rect 45468 65408 45520 65414
rect 45468 65350 45520 65356
rect 45480 64938 45508 65350
rect 45468 64932 45520 64938
rect 45468 64874 45520 64880
rect 45572 64818 45600 68342
rect 45480 64790 45600 64818
rect 45376 63776 45428 63782
rect 45376 63718 45428 63724
rect 45284 48340 45336 48346
rect 45284 48282 45336 48288
rect 45388 46918 45416 63718
rect 45480 63578 45508 64790
rect 45468 63572 45520 63578
rect 45468 63514 45520 63520
rect 45480 62150 45508 63514
rect 45468 62144 45520 62150
rect 45468 62086 45520 62092
rect 45560 56772 45612 56778
rect 45560 56714 45612 56720
rect 45572 52698 45600 56714
rect 45744 56432 45796 56438
rect 45744 56374 45796 56380
rect 45560 52692 45612 52698
rect 45560 52634 45612 52640
rect 45376 46912 45428 46918
rect 45376 46854 45428 46860
rect 45112 45526 45232 45554
rect 45100 44260 45152 44266
rect 45100 44202 45152 44208
rect 45112 43314 45140 44202
rect 45100 43308 45152 43314
rect 45100 43250 45152 43256
rect 45204 39982 45232 45526
rect 45192 39976 45244 39982
rect 45192 39918 45244 39924
rect 45008 32224 45060 32230
rect 45008 32166 45060 32172
rect 45008 29572 45060 29578
rect 45008 29514 45060 29520
rect 45020 29306 45048 29514
rect 45008 29300 45060 29306
rect 45008 29242 45060 29248
rect 45100 29300 45152 29306
rect 45100 29242 45152 29248
rect 45008 26920 45060 26926
rect 45008 26862 45060 26868
rect 45020 19310 45048 26862
rect 45112 25770 45140 29242
rect 45100 25764 45152 25770
rect 45100 25706 45152 25712
rect 45284 20324 45336 20330
rect 45284 20266 45336 20272
rect 45296 19854 45324 20266
rect 45284 19848 45336 19854
rect 45284 19790 45336 19796
rect 45098 19544 45154 19553
rect 45098 19479 45154 19488
rect 45112 19378 45140 19479
rect 45100 19372 45152 19378
rect 45100 19314 45152 19320
rect 45008 19304 45060 19310
rect 45008 19246 45060 19252
rect 45192 19304 45244 19310
rect 45192 19246 45244 19252
rect 45204 18902 45232 19246
rect 45192 18896 45244 18902
rect 45192 18838 45244 18844
rect 44876 14436 44956 14464
rect 45008 14476 45060 14482
rect 44824 14418 44876 14424
rect 45008 14418 45060 14424
rect 44546 14376 44602 14385
rect 44546 14311 44548 14320
rect 44600 14311 44602 14320
rect 44548 14282 44600 14288
rect 44744 14226 44772 14418
rect 45020 14226 45048 14418
rect 44744 14198 45048 14226
rect 44744 13734 44772 14198
rect 44732 13728 44784 13734
rect 44732 13670 44784 13676
rect 44180 11620 44232 11626
rect 44180 11562 44232 11568
rect 44192 11218 44220 11562
rect 44456 11280 44508 11286
rect 44456 11222 44508 11228
rect 44088 11212 44140 11218
rect 44088 11154 44140 11160
rect 44180 11212 44232 11218
rect 44180 11154 44232 11160
rect 44100 7206 44128 11154
rect 44468 11082 44496 11222
rect 44456 11076 44508 11082
rect 44456 11018 44508 11024
rect 44364 9512 44416 9518
rect 44364 9454 44416 9460
rect 44088 7200 44140 7206
rect 44088 7142 44140 7148
rect 44100 4690 44128 7142
rect 44088 4684 44140 4690
rect 44088 4626 44140 4632
rect 43996 3936 44048 3942
rect 43996 3878 44048 3884
rect 43812 2576 43864 2582
rect 43812 2518 43864 2524
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 44008 800 44036 3878
rect 44180 2916 44232 2922
rect 44180 2858 44232 2864
rect 44192 800 44220 2858
rect 44376 2582 44404 9454
rect 44468 9450 44496 11018
rect 44456 9444 44508 9450
rect 44456 9386 44508 9392
rect 45100 7812 45152 7818
rect 45100 7754 45152 7760
rect 44548 4684 44600 4690
rect 44548 4626 44600 4632
rect 44364 2576 44416 2582
rect 44364 2518 44416 2524
rect 44364 1420 44416 1426
rect 44364 1362 44416 1368
rect 44376 800 44404 1362
rect 44560 800 44588 4626
rect 44824 3596 44876 3602
rect 44824 3538 44876 3544
rect 44836 800 44864 3538
rect 45008 2644 45060 2650
rect 45008 2586 45060 2592
rect 45020 800 45048 2586
rect 45112 2582 45140 7754
rect 45204 6798 45232 18838
rect 45296 9518 45324 19790
rect 45374 19408 45430 19417
rect 45374 19343 45376 19352
rect 45428 19343 45430 19352
rect 45376 19314 45428 19320
rect 45374 14376 45430 14385
rect 45374 14311 45376 14320
rect 45428 14311 45430 14320
rect 45376 14282 45428 14288
rect 45284 9512 45336 9518
rect 45284 9454 45336 9460
rect 45652 9512 45704 9518
rect 45652 9454 45704 9460
rect 45192 6792 45244 6798
rect 45192 6734 45244 6740
rect 45192 4004 45244 4010
rect 45192 3946 45244 3952
rect 45100 2576 45152 2582
rect 45100 2518 45152 2524
rect 45204 800 45232 3946
rect 45560 2916 45612 2922
rect 45560 2858 45612 2864
rect 45376 2848 45428 2854
rect 45376 2790 45428 2796
rect 45388 800 45416 2790
rect 45572 800 45600 2858
rect 45664 2106 45692 9454
rect 45756 2990 45784 56374
rect 46020 48000 46072 48006
rect 46020 47942 46072 47948
rect 45928 44736 45980 44742
rect 45928 44678 45980 44684
rect 45836 4684 45888 4690
rect 45836 4626 45888 4632
rect 45744 2984 45796 2990
rect 45744 2926 45796 2932
rect 45652 2100 45704 2106
rect 45652 2042 45704 2048
rect 45848 800 45876 4626
rect 45940 2582 45968 44678
rect 46032 23118 46060 47942
rect 46124 42770 46152 96494
rect 46400 96218 46428 99200
rect 47320 97238 47348 99200
rect 48148 97238 48176 99200
rect 47308 97232 47360 97238
rect 47308 97174 47360 97180
rect 48136 97232 48188 97238
rect 48136 97174 48188 97180
rect 48320 97164 48372 97170
rect 48320 97106 48372 97112
rect 47584 97028 47636 97034
rect 47584 96970 47636 96976
rect 46480 96552 46532 96558
rect 46480 96494 46532 96500
rect 46756 96552 46808 96558
rect 46756 96494 46808 96500
rect 47032 96552 47084 96558
rect 47032 96494 47084 96500
rect 47216 96552 47268 96558
rect 47216 96494 47268 96500
rect 46388 96212 46440 96218
rect 46388 96154 46440 96160
rect 46492 91798 46520 96494
rect 46768 95674 46796 96494
rect 46848 96076 46900 96082
rect 46848 96018 46900 96024
rect 46756 95668 46808 95674
rect 46756 95610 46808 95616
rect 46480 91792 46532 91798
rect 46480 91734 46532 91740
rect 46860 89962 46888 96018
rect 46848 89956 46900 89962
rect 46848 89898 46900 89904
rect 46860 86698 46888 89898
rect 46848 86692 46900 86698
rect 46848 86634 46900 86640
rect 46296 86352 46348 86358
rect 46296 86294 46348 86300
rect 46308 85202 46336 86294
rect 46492 85202 46796 85218
rect 46296 85196 46348 85202
rect 46296 85138 46348 85144
rect 46492 85196 46808 85202
rect 46492 85190 46756 85196
rect 46308 79626 46336 85138
rect 46492 84998 46520 85190
rect 46756 85138 46808 85144
rect 46572 85128 46624 85134
rect 46572 85070 46624 85076
rect 46940 85128 46992 85134
rect 46940 85070 46992 85076
rect 46480 84992 46532 84998
rect 46480 84934 46532 84940
rect 46584 84194 46612 85070
rect 46584 84166 46704 84194
rect 46676 80054 46704 84166
rect 46676 80026 46796 80054
rect 46296 79620 46348 79626
rect 46296 79562 46348 79568
rect 46204 68468 46256 68474
rect 46204 68410 46256 68416
rect 46216 68134 46244 68410
rect 46388 68332 46440 68338
rect 46388 68274 46440 68280
rect 46204 68128 46256 68134
rect 46204 68070 46256 68076
rect 46400 60734 46428 68274
rect 46768 65686 46796 80026
rect 46848 68264 46900 68270
rect 46848 68206 46900 68212
rect 46756 65680 46808 65686
rect 46756 65622 46808 65628
rect 46768 65074 46796 65622
rect 46756 65068 46808 65074
rect 46756 65010 46808 65016
rect 46400 60706 46520 60734
rect 46296 53032 46348 53038
rect 46296 52974 46348 52980
rect 46204 49224 46256 49230
rect 46204 49166 46256 49172
rect 46112 42764 46164 42770
rect 46112 42706 46164 42712
rect 46112 27464 46164 27470
rect 46112 27406 46164 27412
rect 46124 27062 46152 27406
rect 46112 27056 46164 27062
rect 46112 26998 46164 27004
rect 46020 23112 46072 23118
rect 46020 23054 46072 23060
rect 46112 19712 46164 19718
rect 46112 19654 46164 19660
rect 46124 19378 46152 19654
rect 46112 19372 46164 19378
rect 46112 19314 46164 19320
rect 46216 16454 46244 49166
rect 46308 37806 46336 52974
rect 46492 52562 46520 60706
rect 46860 56778 46888 68206
rect 46952 66638 46980 85070
rect 46940 66632 46992 66638
rect 46940 66574 46992 66580
rect 46940 57384 46992 57390
rect 46940 57326 46992 57332
rect 46848 56772 46900 56778
rect 46848 56714 46900 56720
rect 46952 54874 46980 57326
rect 46940 54868 46992 54874
rect 46940 54810 46992 54816
rect 46756 54052 46808 54058
rect 46756 53994 46808 54000
rect 46768 52970 46796 53994
rect 46848 53984 46900 53990
rect 46848 53926 46900 53932
rect 46860 53038 46888 53926
rect 46848 53032 46900 53038
rect 46848 52974 46900 52980
rect 46756 52964 46808 52970
rect 46756 52906 46808 52912
rect 46480 52556 46532 52562
rect 46480 52498 46532 52504
rect 46768 45554 46796 52906
rect 47044 49162 47072 96494
rect 47032 49156 47084 49162
rect 47032 49098 47084 49104
rect 46676 45526 46796 45554
rect 46676 37874 46704 45526
rect 46848 44192 46900 44198
rect 46848 44134 46900 44140
rect 46756 38412 46808 38418
rect 46756 38354 46808 38360
rect 46664 37868 46716 37874
rect 46664 37810 46716 37816
rect 46296 37800 46348 37806
rect 46296 37742 46348 37748
rect 46572 37800 46624 37806
rect 46572 37742 46624 37748
rect 46308 29850 46336 37742
rect 46296 29844 46348 29850
rect 46296 29786 46348 29792
rect 46308 29578 46336 29786
rect 46296 29572 46348 29578
rect 46296 29514 46348 29520
rect 46584 29510 46612 37742
rect 46676 29646 46704 37810
rect 46664 29640 46716 29646
rect 46664 29582 46716 29588
rect 46572 29504 46624 29510
rect 46572 29446 46624 29452
rect 46296 26988 46348 26994
rect 46296 26930 46348 26936
rect 46308 26790 46336 26930
rect 46296 26784 46348 26790
rect 46296 26726 46348 26732
rect 46480 17128 46532 17134
rect 46480 17070 46532 17076
rect 46204 16448 46256 16454
rect 46204 16390 46256 16396
rect 46296 5296 46348 5302
rect 46296 5238 46348 5244
rect 46020 4072 46072 4078
rect 46020 4014 46072 4020
rect 45928 2576 45980 2582
rect 45928 2518 45980 2524
rect 46032 800 46060 4014
rect 46308 3602 46336 5238
rect 46388 3936 46440 3942
rect 46388 3878 46440 3884
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 46204 2372 46256 2378
rect 46204 2314 46256 2320
rect 46112 2304 46164 2310
rect 46112 2246 46164 2252
rect 46124 1426 46152 2246
rect 46112 1420 46164 1426
rect 46112 1362 46164 1368
rect 46216 800 46244 2314
rect 46400 800 46428 3878
rect 46492 2514 46520 17070
rect 46664 14272 46716 14278
rect 46664 14214 46716 14220
rect 46676 13938 46704 14214
rect 46664 13932 46716 13938
rect 46664 13874 46716 13880
rect 46768 3670 46796 38354
rect 46860 37806 46888 44134
rect 47032 40112 47084 40118
rect 47032 40054 47084 40060
rect 47044 37942 47072 40054
rect 47032 37936 47084 37942
rect 47032 37878 47084 37884
rect 46848 37800 46900 37806
rect 46848 37742 46900 37748
rect 46848 29300 46900 29306
rect 46848 29242 46900 29248
rect 46860 29102 46888 29242
rect 46848 29096 46900 29102
rect 46848 29038 46900 29044
rect 46848 25152 46900 25158
rect 46848 25094 46900 25100
rect 46860 18630 46888 25094
rect 46848 18624 46900 18630
rect 46848 18566 46900 18572
rect 47228 11286 47256 96494
rect 47492 96416 47544 96422
rect 47492 96358 47544 96364
rect 47308 32428 47360 32434
rect 47308 32370 47360 32376
rect 47216 11280 47268 11286
rect 47216 11222 47268 11228
rect 47032 4684 47084 4690
rect 47032 4626 47084 4632
rect 46756 3664 46808 3670
rect 46756 3606 46808 3612
rect 46572 3596 46624 3602
rect 46572 3538 46624 3544
rect 46480 2508 46532 2514
rect 46480 2450 46532 2456
rect 46584 800 46612 3538
rect 46848 1420 46900 1426
rect 46848 1362 46900 1368
rect 46860 800 46888 1362
rect 47044 800 47072 4626
rect 47216 3528 47268 3534
rect 47216 3470 47268 3476
rect 47228 800 47256 3470
rect 47320 3194 47348 32370
rect 47400 22024 47452 22030
rect 47400 21966 47452 21972
rect 47412 18766 47440 21966
rect 47400 18760 47452 18766
rect 47400 18702 47452 18708
rect 47504 11150 47532 96358
rect 47596 84114 47624 96970
rect 47952 91520 48004 91526
rect 47952 91462 48004 91468
rect 47584 84108 47636 84114
rect 47584 84050 47636 84056
rect 47676 76492 47728 76498
rect 47676 76434 47728 76440
rect 47584 69216 47636 69222
rect 47584 69158 47636 69164
rect 47596 56438 47624 69158
rect 47584 56432 47636 56438
rect 47584 56374 47636 56380
rect 47584 50856 47636 50862
rect 47584 50798 47636 50804
rect 47596 50726 47624 50798
rect 47584 50720 47636 50726
rect 47584 50662 47636 50668
rect 47596 45422 47624 50662
rect 47584 45416 47636 45422
rect 47584 45358 47636 45364
rect 47584 22500 47636 22506
rect 47584 22442 47636 22448
rect 47492 11144 47544 11150
rect 47492 11086 47544 11092
rect 47596 9382 47624 22442
rect 47688 16794 47716 76434
rect 47964 63782 47992 91462
rect 47952 63776 48004 63782
rect 47952 63718 48004 63724
rect 47768 56160 47820 56166
rect 47768 56102 47820 56108
rect 47780 55622 47808 56102
rect 47768 55616 47820 55622
rect 47768 55558 47820 55564
rect 48044 50924 48096 50930
rect 48044 50866 48096 50872
rect 48056 50454 48084 50866
rect 48044 50448 48096 50454
rect 48044 50390 48096 50396
rect 48228 49700 48280 49706
rect 48228 49642 48280 49648
rect 48240 49162 48268 49642
rect 48228 49156 48280 49162
rect 48228 49098 48280 49104
rect 48136 41200 48188 41206
rect 48136 41142 48188 41148
rect 48148 38418 48176 41142
rect 48136 38412 48188 38418
rect 48136 38354 48188 38360
rect 48044 34604 48096 34610
rect 48044 34546 48096 34552
rect 47952 22092 48004 22098
rect 47952 22034 48004 22040
rect 47964 22001 47992 22034
rect 47950 21992 48006 22001
rect 47950 21927 48006 21936
rect 48056 16794 48084 34546
rect 48148 31278 48176 38354
rect 48136 31272 48188 31278
rect 48136 31214 48188 31220
rect 48332 29782 48360 97106
rect 49068 96626 49096 99200
rect 49896 97170 49924 99200
rect 50300 97404 50596 97424
rect 50356 97402 50380 97404
rect 50436 97402 50460 97404
rect 50516 97402 50540 97404
rect 50378 97350 50380 97402
rect 50442 97350 50454 97402
rect 50516 97350 50518 97402
rect 50356 97348 50380 97350
rect 50436 97348 50460 97350
rect 50516 97348 50540 97350
rect 50300 97328 50596 97348
rect 50816 97238 50844 99200
rect 50804 97232 50856 97238
rect 50804 97174 50856 97180
rect 49884 97164 49936 97170
rect 49884 97106 49936 97112
rect 50896 97164 50948 97170
rect 50896 97106 50948 97112
rect 49056 96620 49108 96626
rect 49056 96562 49108 96568
rect 49148 96484 49200 96490
rect 49148 96426 49200 96432
rect 49160 96218 49188 96426
rect 50300 96316 50596 96336
rect 50356 96314 50380 96316
rect 50436 96314 50460 96316
rect 50516 96314 50540 96316
rect 50378 96262 50380 96314
rect 50442 96262 50454 96314
rect 50516 96262 50518 96314
rect 50356 96260 50380 96262
rect 50436 96260 50460 96262
rect 50516 96260 50540 96262
rect 50300 96240 50596 96260
rect 49148 96212 49200 96218
rect 49148 96154 49200 96160
rect 50300 95228 50596 95248
rect 50356 95226 50380 95228
rect 50436 95226 50460 95228
rect 50516 95226 50540 95228
rect 50378 95174 50380 95226
rect 50442 95174 50454 95226
rect 50516 95174 50518 95226
rect 50356 95172 50380 95174
rect 50436 95172 50460 95174
rect 50516 95172 50540 95174
rect 50300 95152 50596 95172
rect 50300 94140 50596 94160
rect 50356 94138 50380 94140
rect 50436 94138 50460 94140
rect 50516 94138 50540 94140
rect 50378 94086 50380 94138
rect 50442 94086 50454 94138
rect 50516 94086 50518 94138
rect 50356 94084 50380 94086
rect 50436 94084 50460 94086
rect 50516 94084 50540 94086
rect 50300 94064 50596 94084
rect 49884 93968 49936 93974
rect 49884 93910 49936 93916
rect 49056 91860 49108 91866
rect 49056 91802 49108 91808
rect 48964 91792 49016 91798
rect 48964 91734 49016 91740
rect 48976 89622 49004 91734
rect 48964 89616 49016 89622
rect 48964 89558 49016 89564
rect 48976 78130 49004 89558
rect 49068 86290 49096 91802
rect 49700 88596 49752 88602
rect 49700 88538 49752 88544
rect 49056 86284 49108 86290
rect 49056 86226 49108 86232
rect 49068 78538 49096 86226
rect 49608 80232 49660 80238
rect 49608 80174 49660 80180
rect 49056 78532 49108 78538
rect 49056 78474 49108 78480
rect 48964 78124 49016 78130
rect 48964 78066 49016 78072
rect 48780 73160 48832 73166
rect 48780 73102 48832 73108
rect 48792 72214 48820 73102
rect 48780 72208 48832 72214
rect 48780 72150 48832 72156
rect 48792 61742 48820 72150
rect 48976 63510 49004 78066
rect 48964 63504 49016 63510
rect 48964 63446 49016 63452
rect 48780 61736 48832 61742
rect 48780 61678 48832 61684
rect 48780 56228 48832 56234
rect 48780 56170 48832 56176
rect 48792 55690 48820 56170
rect 49068 55690 49096 78474
rect 49516 66088 49568 66094
rect 49516 66030 49568 66036
rect 49422 64560 49478 64569
rect 49422 64495 49424 64504
rect 49476 64495 49478 64504
rect 49424 64466 49476 64472
rect 49436 64054 49464 64466
rect 49528 64462 49556 66030
rect 49516 64456 49568 64462
rect 49516 64398 49568 64404
rect 49424 64048 49476 64054
rect 49424 63990 49476 63996
rect 49516 63504 49568 63510
rect 49516 63446 49568 63452
rect 49528 62286 49556 63446
rect 49620 62354 49648 80174
rect 49712 80170 49740 88538
rect 49792 80232 49844 80238
rect 49792 80174 49844 80180
rect 49700 80164 49752 80170
rect 49700 80106 49752 80112
rect 49700 64660 49752 64666
rect 49700 64602 49752 64608
rect 49712 64122 49740 64602
rect 49700 64116 49752 64122
rect 49700 64058 49752 64064
rect 49712 63850 49740 64058
rect 49700 63844 49752 63850
rect 49700 63786 49752 63792
rect 49608 62348 49660 62354
rect 49608 62290 49660 62296
rect 49516 62280 49568 62286
rect 49516 62222 49568 62228
rect 49528 55826 49556 62222
rect 49608 61668 49660 61674
rect 49608 61610 49660 61616
rect 49148 55820 49200 55826
rect 49148 55762 49200 55768
rect 49516 55820 49568 55826
rect 49516 55762 49568 55768
rect 48780 55684 48832 55690
rect 48780 55626 48832 55632
rect 49056 55684 49108 55690
rect 49056 55626 49108 55632
rect 49160 55214 49188 55762
rect 49160 55186 49280 55214
rect 48412 49768 48464 49774
rect 48412 49710 48464 49716
rect 48424 38282 48452 49710
rect 48964 48884 49016 48890
rect 48964 48826 49016 48832
rect 48976 40118 49004 48826
rect 48964 40112 49016 40118
rect 48964 40054 49016 40060
rect 48504 38412 48556 38418
rect 48504 38354 48556 38360
rect 48412 38276 48464 38282
rect 48412 38218 48464 38224
rect 48516 38162 48544 38354
rect 48424 38134 48544 38162
rect 48424 37874 48452 38134
rect 48412 37868 48464 37874
rect 48412 37810 48464 37816
rect 48424 36650 48452 37810
rect 48412 36644 48464 36650
rect 48412 36586 48464 36592
rect 48320 29776 48372 29782
rect 48320 29718 48372 29724
rect 48332 22506 48360 29718
rect 48320 22500 48372 22506
rect 48320 22442 48372 22448
rect 48424 17954 48452 36586
rect 49252 23594 49280 55186
rect 49516 51060 49568 51066
rect 49516 51002 49568 51008
rect 49528 49910 49556 51002
rect 49516 49904 49568 49910
rect 49516 49846 49568 49852
rect 49528 49774 49556 49846
rect 49516 49768 49568 49774
rect 49516 49710 49568 49716
rect 49424 42764 49476 42770
rect 49424 42706 49476 42712
rect 49436 41614 49464 42706
rect 49424 41608 49476 41614
rect 49424 41550 49476 41556
rect 49436 28014 49464 41550
rect 49620 38418 49648 61610
rect 49700 55820 49752 55826
rect 49700 55762 49752 55768
rect 49712 55622 49740 55762
rect 49700 55616 49752 55622
rect 49700 55558 49752 55564
rect 49712 55282 49740 55558
rect 49700 55276 49752 55282
rect 49700 55218 49752 55224
rect 49700 40044 49752 40050
rect 49700 39986 49752 39992
rect 49712 39642 49740 39986
rect 49700 39636 49752 39642
rect 49700 39578 49752 39584
rect 49608 38412 49660 38418
rect 49608 38354 49660 38360
rect 49516 37800 49568 37806
rect 49516 37742 49568 37748
rect 49424 28008 49476 28014
rect 49424 27950 49476 27956
rect 49424 23792 49476 23798
rect 49424 23734 49476 23740
rect 49240 23588 49292 23594
rect 49240 23530 49292 23536
rect 48964 23520 49016 23526
rect 48964 23462 49016 23468
rect 48872 22568 48924 22574
rect 48872 22510 48924 22516
rect 48884 21622 48912 22510
rect 48872 21616 48924 21622
rect 48872 21558 48924 21564
rect 48424 17926 48544 17954
rect 48320 17672 48372 17678
rect 48320 17614 48372 17620
rect 48332 16794 48360 17614
rect 47676 16788 47728 16794
rect 47676 16730 47728 16736
rect 48044 16788 48096 16794
rect 48044 16730 48096 16736
rect 48320 16788 48372 16794
rect 48320 16730 48372 16736
rect 48516 16658 48544 17926
rect 48504 16652 48556 16658
rect 48504 16594 48556 16600
rect 48228 11824 48280 11830
rect 48228 11766 48280 11772
rect 48240 11286 48268 11766
rect 48228 11280 48280 11286
rect 48228 11222 48280 11228
rect 48976 9654 49004 23462
rect 49056 17060 49108 17066
rect 49056 17002 49108 17008
rect 48964 9648 49016 9654
rect 48964 9590 49016 9596
rect 47584 9376 47636 9382
rect 47584 9318 47636 9324
rect 49068 9178 49096 17002
rect 49056 9172 49108 9178
rect 49056 9114 49108 9120
rect 48688 6656 48740 6662
rect 48688 6598 48740 6604
rect 48700 6458 48728 6598
rect 48688 6452 48740 6458
rect 48688 6394 48740 6400
rect 47584 4684 47636 4690
rect 47584 4626 47636 4632
rect 48228 4684 48280 4690
rect 48228 4626 48280 4632
rect 47308 3188 47360 3194
rect 47308 3130 47360 3136
rect 47320 2990 47348 3130
rect 47308 2984 47360 2990
rect 47308 2926 47360 2932
rect 47400 2916 47452 2922
rect 47400 2858 47452 2864
rect 47412 800 47440 2858
rect 47596 800 47624 4626
rect 48136 4276 48188 4282
rect 48136 4218 48188 4224
rect 47860 3528 47912 3534
rect 47860 3470 47912 3476
rect 47872 800 47900 3470
rect 48148 2582 48176 4218
rect 48136 2576 48188 2582
rect 48136 2518 48188 2524
rect 48044 2440 48096 2446
rect 48044 2382 48096 2388
rect 47952 2304 48004 2310
rect 47952 2246 48004 2252
rect 47964 1426 47992 2246
rect 47952 1420 48004 1426
rect 47952 1362 48004 1368
rect 48056 800 48084 2382
rect 48240 800 48268 4626
rect 48504 4480 48556 4486
rect 48504 4422 48556 4428
rect 48412 4072 48464 4078
rect 48412 4014 48464 4020
rect 48424 800 48452 4014
rect 48516 2582 48544 4422
rect 48872 4072 48924 4078
rect 48872 4014 48924 4020
rect 48504 2576 48556 2582
rect 48504 2518 48556 2524
rect 48688 2100 48740 2106
rect 48688 2042 48740 2048
rect 48700 800 48728 2042
rect 48884 800 48912 4014
rect 49056 3596 49108 3602
rect 49056 3538 49108 3544
rect 49068 800 49096 3538
rect 49240 2916 49292 2922
rect 49240 2858 49292 2864
rect 49252 800 49280 2858
rect 49436 2650 49464 23734
rect 49528 23526 49556 37742
rect 49608 36916 49660 36922
rect 49608 36858 49660 36864
rect 49620 36718 49648 36858
rect 49608 36712 49660 36718
rect 49608 36654 49660 36660
rect 49620 25838 49648 36654
rect 49608 25832 49660 25838
rect 49608 25774 49660 25780
rect 49700 25764 49752 25770
rect 49700 25706 49752 25712
rect 49516 23520 49568 23526
rect 49516 23462 49568 23468
rect 49516 22704 49568 22710
rect 49516 22646 49568 22652
rect 49528 2990 49556 22646
rect 49712 16658 49740 25706
rect 49700 16652 49752 16658
rect 49700 16594 49752 16600
rect 49700 14272 49752 14278
rect 49700 14214 49752 14220
rect 49608 14000 49660 14006
rect 49608 13942 49660 13948
rect 49620 9042 49648 13942
rect 49712 13938 49740 14214
rect 49700 13932 49752 13938
rect 49700 13874 49752 13880
rect 49608 9036 49660 9042
rect 49608 8978 49660 8984
rect 49608 4072 49660 4078
rect 49608 4014 49660 4020
rect 49516 2984 49568 2990
rect 49516 2926 49568 2932
rect 49620 2774 49648 4014
rect 49700 3596 49752 3602
rect 49700 3538 49752 3544
rect 49528 2746 49648 2774
rect 49424 2644 49476 2650
rect 49424 2586 49476 2592
rect 49528 898 49556 2746
rect 49436 870 49556 898
rect 49436 800 49464 870
rect 49712 800 49740 3538
rect 49804 1358 49832 80174
rect 49896 66094 49924 93910
rect 50300 93052 50596 93072
rect 50356 93050 50380 93052
rect 50436 93050 50460 93052
rect 50516 93050 50540 93052
rect 50378 92998 50380 93050
rect 50442 92998 50454 93050
rect 50516 92998 50518 93050
rect 50356 92996 50380 92998
rect 50436 92996 50460 92998
rect 50516 92996 50540 92998
rect 50300 92976 50596 92996
rect 50300 91964 50596 91984
rect 50356 91962 50380 91964
rect 50436 91962 50460 91964
rect 50516 91962 50540 91964
rect 50378 91910 50380 91962
rect 50442 91910 50454 91962
rect 50516 91910 50518 91962
rect 50356 91908 50380 91910
rect 50436 91908 50460 91910
rect 50516 91908 50540 91910
rect 50300 91888 50596 91908
rect 50300 90876 50596 90896
rect 50356 90874 50380 90876
rect 50436 90874 50460 90876
rect 50516 90874 50540 90876
rect 50378 90822 50380 90874
rect 50442 90822 50454 90874
rect 50516 90822 50518 90874
rect 50356 90820 50380 90822
rect 50436 90820 50460 90822
rect 50516 90820 50540 90822
rect 50300 90800 50596 90820
rect 49976 90160 50028 90166
rect 49976 90102 50028 90108
rect 49988 67634 50016 90102
rect 50300 89788 50596 89808
rect 50356 89786 50380 89788
rect 50436 89786 50460 89788
rect 50516 89786 50540 89788
rect 50378 89734 50380 89786
rect 50442 89734 50454 89786
rect 50516 89734 50518 89786
rect 50356 89732 50380 89734
rect 50436 89732 50460 89734
rect 50516 89732 50540 89734
rect 50300 89712 50596 89732
rect 50068 88800 50120 88806
rect 50068 88742 50120 88748
rect 50080 84194 50108 88742
rect 50300 88700 50596 88720
rect 50356 88698 50380 88700
rect 50436 88698 50460 88700
rect 50516 88698 50540 88700
rect 50378 88646 50380 88698
rect 50442 88646 50454 88698
rect 50516 88646 50518 88698
rect 50356 88644 50380 88646
rect 50436 88644 50460 88646
rect 50516 88644 50540 88646
rect 50300 88624 50596 88644
rect 50300 87612 50596 87632
rect 50356 87610 50380 87612
rect 50436 87610 50460 87612
rect 50516 87610 50540 87612
rect 50378 87558 50380 87610
rect 50442 87558 50454 87610
rect 50516 87558 50518 87610
rect 50356 87556 50380 87558
rect 50436 87556 50460 87558
rect 50516 87556 50540 87558
rect 50300 87536 50596 87556
rect 50300 86524 50596 86544
rect 50356 86522 50380 86524
rect 50436 86522 50460 86524
rect 50516 86522 50540 86524
rect 50378 86470 50380 86522
rect 50442 86470 50454 86522
rect 50516 86470 50518 86522
rect 50356 86468 50380 86470
rect 50436 86468 50460 86470
rect 50516 86468 50540 86470
rect 50300 86448 50596 86468
rect 50300 85436 50596 85456
rect 50356 85434 50380 85436
rect 50436 85434 50460 85436
rect 50516 85434 50540 85436
rect 50378 85382 50380 85434
rect 50442 85382 50454 85434
rect 50516 85382 50518 85434
rect 50356 85380 50380 85382
rect 50436 85380 50460 85382
rect 50516 85380 50540 85382
rect 50300 85360 50596 85380
rect 50160 85332 50212 85338
rect 50160 85274 50212 85280
rect 50172 84726 50200 85274
rect 50160 84720 50212 84726
rect 50160 84662 50212 84668
rect 50300 84348 50596 84368
rect 50356 84346 50380 84348
rect 50436 84346 50460 84348
rect 50516 84346 50540 84348
rect 50378 84294 50380 84346
rect 50442 84294 50454 84346
rect 50516 84294 50518 84346
rect 50356 84292 50380 84294
rect 50436 84292 50460 84294
rect 50516 84292 50540 84294
rect 50300 84272 50596 84292
rect 50080 84166 50200 84194
rect 50172 80238 50200 84166
rect 50300 83260 50596 83280
rect 50356 83258 50380 83260
rect 50436 83258 50460 83260
rect 50516 83258 50540 83260
rect 50378 83206 50380 83258
rect 50442 83206 50454 83258
rect 50516 83206 50518 83258
rect 50356 83204 50380 83206
rect 50436 83204 50460 83206
rect 50516 83204 50540 83206
rect 50300 83184 50596 83204
rect 50300 82172 50596 82192
rect 50356 82170 50380 82172
rect 50436 82170 50460 82172
rect 50516 82170 50540 82172
rect 50378 82118 50380 82170
rect 50442 82118 50454 82170
rect 50516 82118 50518 82170
rect 50356 82116 50380 82118
rect 50436 82116 50460 82118
rect 50516 82116 50540 82118
rect 50300 82096 50596 82116
rect 50300 81084 50596 81104
rect 50356 81082 50380 81084
rect 50436 81082 50460 81084
rect 50516 81082 50540 81084
rect 50378 81030 50380 81082
rect 50442 81030 50454 81082
rect 50516 81030 50518 81082
rect 50356 81028 50380 81030
rect 50436 81028 50460 81030
rect 50516 81028 50540 81030
rect 50300 81008 50596 81028
rect 50068 80232 50120 80238
rect 50068 80174 50120 80180
rect 50160 80232 50212 80238
rect 50160 80174 50212 80180
rect 50080 72554 50108 80174
rect 50712 80164 50764 80170
rect 50712 80106 50764 80112
rect 50300 79996 50596 80016
rect 50356 79994 50380 79996
rect 50436 79994 50460 79996
rect 50516 79994 50540 79996
rect 50378 79942 50380 79994
rect 50442 79942 50454 79994
rect 50516 79942 50518 79994
rect 50356 79940 50380 79942
rect 50436 79940 50460 79942
rect 50516 79940 50540 79942
rect 50300 79920 50596 79940
rect 50300 78908 50596 78928
rect 50356 78906 50380 78908
rect 50436 78906 50460 78908
rect 50516 78906 50540 78908
rect 50378 78854 50380 78906
rect 50442 78854 50454 78906
rect 50516 78854 50518 78906
rect 50356 78852 50380 78854
rect 50436 78852 50460 78854
rect 50516 78852 50540 78854
rect 50300 78832 50596 78852
rect 50300 77820 50596 77840
rect 50356 77818 50380 77820
rect 50436 77818 50460 77820
rect 50516 77818 50540 77820
rect 50378 77766 50380 77818
rect 50442 77766 50454 77818
rect 50516 77766 50518 77818
rect 50356 77764 50380 77766
rect 50436 77764 50460 77766
rect 50516 77764 50540 77766
rect 50300 77744 50596 77764
rect 50300 76732 50596 76752
rect 50356 76730 50380 76732
rect 50436 76730 50460 76732
rect 50516 76730 50540 76732
rect 50378 76678 50380 76730
rect 50442 76678 50454 76730
rect 50516 76678 50518 76730
rect 50356 76676 50380 76678
rect 50436 76676 50460 76678
rect 50516 76676 50540 76678
rect 50300 76656 50596 76676
rect 50300 75644 50596 75664
rect 50356 75642 50380 75644
rect 50436 75642 50460 75644
rect 50516 75642 50540 75644
rect 50378 75590 50380 75642
rect 50442 75590 50454 75642
rect 50516 75590 50518 75642
rect 50356 75588 50380 75590
rect 50436 75588 50460 75590
rect 50516 75588 50540 75590
rect 50300 75568 50596 75588
rect 50300 74556 50596 74576
rect 50356 74554 50380 74556
rect 50436 74554 50460 74556
rect 50516 74554 50540 74556
rect 50378 74502 50380 74554
rect 50442 74502 50454 74554
rect 50516 74502 50518 74554
rect 50356 74500 50380 74502
rect 50436 74500 50460 74502
rect 50516 74500 50540 74502
rect 50300 74480 50596 74500
rect 50300 73468 50596 73488
rect 50356 73466 50380 73468
rect 50436 73466 50460 73468
rect 50516 73466 50540 73468
rect 50378 73414 50380 73466
rect 50442 73414 50454 73466
rect 50516 73414 50518 73466
rect 50356 73412 50380 73414
rect 50436 73412 50460 73414
rect 50516 73412 50540 73414
rect 50300 73392 50596 73412
rect 50068 72548 50120 72554
rect 50068 72490 50120 72496
rect 50620 72548 50672 72554
rect 50620 72490 50672 72496
rect 50300 72380 50596 72400
rect 50356 72378 50380 72380
rect 50436 72378 50460 72380
rect 50516 72378 50540 72380
rect 50378 72326 50380 72378
rect 50442 72326 50454 72378
rect 50516 72326 50518 72378
rect 50356 72324 50380 72326
rect 50436 72324 50460 72326
rect 50516 72324 50540 72326
rect 50300 72304 50596 72324
rect 50300 71292 50596 71312
rect 50356 71290 50380 71292
rect 50436 71290 50460 71292
rect 50516 71290 50540 71292
rect 50378 71238 50380 71290
rect 50442 71238 50454 71290
rect 50516 71238 50518 71290
rect 50356 71236 50380 71238
rect 50436 71236 50460 71238
rect 50516 71236 50540 71238
rect 50300 71216 50596 71236
rect 50300 70204 50596 70224
rect 50356 70202 50380 70204
rect 50436 70202 50460 70204
rect 50516 70202 50540 70204
rect 50378 70150 50380 70202
rect 50442 70150 50454 70202
rect 50516 70150 50518 70202
rect 50356 70148 50380 70150
rect 50436 70148 50460 70150
rect 50516 70148 50540 70150
rect 50300 70128 50596 70148
rect 50160 69964 50212 69970
rect 50160 69906 50212 69912
rect 49988 67606 50108 67634
rect 49884 66088 49936 66094
rect 49884 66030 49936 66036
rect 50080 64598 50108 67606
rect 50068 64592 50120 64598
rect 50068 64534 50120 64540
rect 49882 64424 49938 64433
rect 49882 64359 49884 64368
rect 49936 64359 49938 64368
rect 49884 64330 49936 64336
rect 50172 64326 50200 69906
rect 50300 69116 50596 69136
rect 50356 69114 50380 69116
rect 50436 69114 50460 69116
rect 50516 69114 50540 69116
rect 50378 69062 50380 69114
rect 50442 69062 50454 69114
rect 50516 69062 50518 69114
rect 50356 69060 50380 69062
rect 50436 69060 50460 69062
rect 50516 69060 50540 69062
rect 50300 69040 50596 69060
rect 50300 68028 50596 68048
rect 50356 68026 50380 68028
rect 50436 68026 50460 68028
rect 50516 68026 50540 68028
rect 50378 67974 50380 68026
rect 50442 67974 50454 68026
rect 50516 67974 50518 68026
rect 50356 67972 50380 67974
rect 50436 67972 50460 67974
rect 50516 67972 50540 67974
rect 50300 67952 50596 67972
rect 50300 66940 50596 66960
rect 50356 66938 50380 66940
rect 50436 66938 50460 66940
rect 50516 66938 50540 66940
rect 50378 66886 50380 66938
rect 50442 66886 50454 66938
rect 50516 66886 50518 66938
rect 50356 66884 50380 66886
rect 50436 66884 50460 66886
rect 50516 66884 50540 66886
rect 50300 66864 50596 66884
rect 50300 65852 50596 65872
rect 50356 65850 50380 65852
rect 50436 65850 50460 65852
rect 50516 65850 50540 65852
rect 50378 65798 50380 65850
rect 50442 65798 50454 65850
rect 50516 65798 50518 65850
rect 50356 65796 50380 65798
rect 50436 65796 50460 65798
rect 50516 65796 50540 65798
rect 50300 65776 50596 65796
rect 50300 64764 50596 64784
rect 50356 64762 50380 64764
rect 50436 64762 50460 64764
rect 50516 64762 50540 64764
rect 50378 64710 50380 64762
rect 50442 64710 50454 64762
rect 50516 64710 50518 64762
rect 50356 64708 50380 64710
rect 50436 64708 50460 64710
rect 50516 64708 50540 64710
rect 50300 64688 50596 64708
rect 50344 64592 50396 64598
rect 50342 64560 50344 64569
rect 50396 64560 50398 64569
rect 50342 64495 50398 64504
rect 50250 64424 50306 64433
rect 50250 64359 50252 64368
rect 50304 64359 50306 64368
rect 50252 64330 50304 64336
rect 49976 64320 50028 64326
rect 49976 64262 50028 64268
rect 50160 64320 50212 64326
rect 50160 64262 50212 64268
rect 49988 64054 50016 64262
rect 49976 64048 50028 64054
rect 49976 63990 50028 63996
rect 50300 63676 50596 63696
rect 50356 63674 50380 63676
rect 50436 63674 50460 63676
rect 50516 63674 50540 63676
rect 50378 63622 50380 63674
rect 50442 63622 50454 63674
rect 50516 63622 50518 63674
rect 50356 63620 50380 63622
rect 50436 63620 50460 63622
rect 50516 63620 50540 63622
rect 50300 63600 50596 63620
rect 50300 62588 50596 62608
rect 50356 62586 50380 62588
rect 50436 62586 50460 62588
rect 50516 62586 50540 62588
rect 50378 62534 50380 62586
rect 50442 62534 50454 62586
rect 50516 62534 50518 62586
rect 50356 62532 50380 62534
rect 50436 62532 50460 62534
rect 50516 62532 50540 62534
rect 50300 62512 50596 62532
rect 50300 61500 50596 61520
rect 50356 61498 50380 61500
rect 50436 61498 50460 61500
rect 50516 61498 50540 61500
rect 50378 61446 50380 61498
rect 50442 61446 50454 61498
rect 50516 61446 50518 61498
rect 50356 61444 50380 61446
rect 50436 61444 50460 61446
rect 50516 61444 50540 61446
rect 50300 61424 50596 61444
rect 50300 60412 50596 60432
rect 50356 60410 50380 60412
rect 50436 60410 50460 60412
rect 50516 60410 50540 60412
rect 50378 60358 50380 60410
rect 50442 60358 50454 60410
rect 50516 60358 50518 60410
rect 50356 60356 50380 60358
rect 50436 60356 50460 60358
rect 50516 60356 50540 60358
rect 50300 60336 50596 60356
rect 50300 59324 50596 59344
rect 50356 59322 50380 59324
rect 50436 59322 50460 59324
rect 50516 59322 50540 59324
rect 50378 59270 50380 59322
rect 50442 59270 50454 59322
rect 50516 59270 50518 59322
rect 50356 59268 50380 59270
rect 50436 59268 50460 59270
rect 50516 59268 50540 59270
rect 50300 59248 50596 59268
rect 50300 58236 50596 58256
rect 50356 58234 50380 58236
rect 50436 58234 50460 58236
rect 50516 58234 50540 58236
rect 50378 58182 50380 58234
rect 50442 58182 50454 58234
rect 50516 58182 50518 58234
rect 50356 58180 50380 58182
rect 50436 58180 50460 58182
rect 50516 58180 50540 58182
rect 50300 58160 50596 58180
rect 50300 57148 50596 57168
rect 50356 57146 50380 57148
rect 50436 57146 50460 57148
rect 50516 57146 50540 57148
rect 50378 57094 50380 57146
rect 50442 57094 50454 57146
rect 50516 57094 50518 57146
rect 50356 57092 50380 57094
rect 50436 57092 50460 57094
rect 50516 57092 50540 57094
rect 50300 57072 50596 57092
rect 50436 56840 50488 56846
rect 50436 56782 50488 56788
rect 50448 56302 50476 56782
rect 49976 56296 50028 56302
rect 49976 56238 50028 56244
rect 50436 56296 50488 56302
rect 50436 56238 50488 56244
rect 49988 18630 50016 56238
rect 50068 56160 50120 56166
rect 50068 56102 50120 56108
rect 50080 40050 50108 56102
rect 50300 56060 50596 56080
rect 50356 56058 50380 56060
rect 50436 56058 50460 56060
rect 50516 56058 50540 56060
rect 50378 56006 50380 56058
rect 50442 56006 50454 56058
rect 50516 56006 50518 56058
rect 50356 56004 50380 56006
rect 50436 56004 50460 56006
rect 50516 56004 50540 56006
rect 50300 55984 50596 56004
rect 50300 54972 50596 54992
rect 50356 54970 50380 54972
rect 50436 54970 50460 54972
rect 50516 54970 50540 54972
rect 50378 54918 50380 54970
rect 50442 54918 50454 54970
rect 50516 54918 50518 54970
rect 50356 54916 50380 54918
rect 50436 54916 50460 54918
rect 50516 54916 50540 54918
rect 50300 54896 50596 54916
rect 50300 53884 50596 53904
rect 50356 53882 50380 53884
rect 50436 53882 50460 53884
rect 50516 53882 50540 53884
rect 50378 53830 50380 53882
rect 50442 53830 50454 53882
rect 50516 53830 50518 53882
rect 50356 53828 50380 53830
rect 50436 53828 50460 53830
rect 50516 53828 50540 53830
rect 50300 53808 50596 53828
rect 50300 52796 50596 52816
rect 50356 52794 50380 52796
rect 50436 52794 50460 52796
rect 50516 52794 50540 52796
rect 50378 52742 50380 52794
rect 50442 52742 50454 52794
rect 50516 52742 50518 52794
rect 50356 52740 50380 52742
rect 50436 52740 50460 52742
rect 50516 52740 50540 52742
rect 50300 52720 50596 52740
rect 50300 51708 50596 51728
rect 50356 51706 50380 51708
rect 50436 51706 50460 51708
rect 50516 51706 50540 51708
rect 50378 51654 50380 51706
rect 50442 51654 50454 51706
rect 50516 51654 50518 51706
rect 50356 51652 50380 51654
rect 50436 51652 50460 51654
rect 50516 51652 50540 51654
rect 50300 51632 50596 51652
rect 50300 50620 50596 50640
rect 50356 50618 50380 50620
rect 50436 50618 50460 50620
rect 50516 50618 50540 50620
rect 50378 50566 50380 50618
rect 50442 50566 50454 50618
rect 50516 50566 50518 50618
rect 50356 50564 50380 50566
rect 50436 50564 50460 50566
rect 50516 50564 50540 50566
rect 50300 50544 50596 50564
rect 50300 49532 50596 49552
rect 50356 49530 50380 49532
rect 50436 49530 50460 49532
rect 50516 49530 50540 49532
rect 50378 49478 50380 49530
rect 50442 49478 50454 49530
rect 50516 49478 50518 49530
rect 50356 49476 50380 49478
rect 50436 49476 50460 49478
rect 50516 49476 50540 49478
rect 50300 49456 50596 49476
rect 50300 48444 50596 48464
rect 50356 48442 50380 48444
rect 50436 48442 50460 48444
rect 50516 48442 50540 48444
rect 50378 48390 50380 48442
rect 50442 48390 50454 48442
rect 50516 48390 50518 48442
rect 50356 48388 50380 48390
rect 50436 48388 50460 48390
rect 50516 48388 50540 48390
rect 50300 48368 50596 48388
rect 50300 47356 50596 47376
rect 50356 47354 50380 47356
rect 50436 47354 50460 47356
rect 50516 47354 50540 47356
rect 50378 47302 50380 47354
rect 50442 47302 50454 47354
rect 50516 47302 50518 47354
rect 50356 47300 50380 47302
rect 50436 47300 50460 47302
rect 50516 47300 50540 47302
rect 50300 47280 50596 47300
rect 50300 46268 50596 46288
rect 50356 46266 50380 46268
rect 50436 46266 50460 46268
rect 50516 46266 50540 46268
rect 50378 46214 50380 46266
rect 50442 46214 50454 46266
rect 50516 46214 50518 46266
rect 50356 46212 50380 46214
rect 50436 46212 50460 46214
rect 50516 46212 50540 46214
rect 50300 46192 50596 46212
rect 50300 45180 50596 45200
rect 50356 45178 50380 45180
rect 50436 45178 50460 45180
rect 50516 45178 50540 45180
rect 50378 45126 50380 45178
rect 50442 45126 50454 45178
rect 50516 45126 50518 45178
rect 50356 45124 50380 45126
rect 50436 45124 50460 45126
rect 50516 45124 50540 45126
rect 50300 45104 50596 45124
rect 50300 44092 50596 44112
rect 50356 44090 50380 44092
rect 50436 44090 50460 44092
rect 50516 44090 50540 44092
rect 50378 44038 50380 44090
rect 50442 44038 50454 44090
rect 50516 44038 50518 44090
rect 50356 44036 50380 44038
rect 50436 44036 50460 44038
rect 50516 44036 50540 44038
rect 50300 44016 50596 44036
rect 50300 43004 50596 43024
rect 50356 43002 50380 43004
rect 50436 43002 50460 43004
rect 50516 43002 50540 43004
rect 50378 42950 50380 43002
rect 50442 42950 50454 43002
rect 50516 42950 50518 43002
rect 50356 42948 50380 42950
rect 50436 42948 50460 42950
rect 50516 42948 50540 42950
rect 50300 42928 50596 42948
rect 50300 41916 50596 41936
rect 50356 41914 50380 41916
rect 50436 41914 50460 41916
rect 50516 41914 50540 41916
rect 50378 41862 50380 41914
rect 50442 41862 50454 41914
rect 50516 41862 50518 41914
rect 50356 41860 50380 41862
rect 50436 41860 50460 41862
rect 50516 41860 50540 41862
rect 50300 41840 50596 41860
rect 50300 40828 50596 40848
rect 50356 40826 50380 40828
rect 50436 40826 50460 40828
rect 50516 40826 50540 40828
rect 50378 40774 50380 40826
rect 50442 40774 50454 40826
rect 50516 40774 50518 40826
rect 50356 40772 50380 40774
rect 50436 40772 50460 40774
rect 50516 40772 50540 40774
rect 50300 40752 50596 40772
rect 50068 40044 50120 40050
rect 50068 39986 50120 39992
rect 50300 39740 50596 39760
rect 50356 39738 50380 39740
rect 50436 39738 50460 39740
rect 50516 39738 50540 39740
rect 50378 39686 50380 39738
rect 50442 39686 50454 39738
rect 50516 39686 50518 39738
rect 50356 39684 50380 39686
rect 50436 39684 50460 39686
rect 50516 39684 50540 39686
rect 50300 39664 50596 39684
rect 50300 38652 50596 38672
rect 50356 38650 50380 38652
rect 50436 38650 50460 38652
rect 50516 38650 50540 38652
rect 50378 38598 50380 38650
rect 50442 38598 50454 38650
rect 50516 38598 50518 38650
rect 50356 38596 50380 38598
rect 50436 38596 50460 38598
rect 50516 38596 50540 38598
rect 50300 38576 50596 38596
rect 50160 37664 50212 37670
rect 50160 37606 50212 37612
rect 50068 21956 50120 21962
rect 50068 21898 50120 21904
rect 50080 20806 50108 21898
rect 50068 20800 50120 20806
rect 50068 20742 50120 20748
rect 49976 18624 50028 18630
rect 49976 18566 50028 18572
rect 50080 5846 50108 20742
rect 50172 19174 50200 37606
rect 50300 37564 50596 37584
rect 50356 37562 50380 37564
rect 50436 37562 50460 37564
rect 50516 37562 50540 37564
rect 50378 37510 50380 37562
rect 50442 37510 50454 37562
rect 50516 37510 50518 37562
rect 50356 37508 50380 37510
rect 50436 37508 50460 37510
rect 50516 37508 50540 37510
rect 50300 37488 50596 37508
rect 50300 36476 50596 36496
rect 50356 36474 50380 36476
rect 50436 36474 50460 36476
rect 50516 36474 50540 36476
rect 50378 36422 50380 36474
rect 50442 36422 50454 36474
rect 50516 36422 50518 36474
rect 50356 36420 50380 36422
rect 50436 36420 50460 36422
rect 50516 36420 50540 36422
rect 50300 36400 50596 36420
rect 50300 35388 50596 35408
rect 50356 35386 50380 35388
rect 50436 35386 50460 35388
rect 50516 35386 50540 35388
rect 50378 35334 50380 35386
rect 50442 35334 50454 35386
rect 50516 35334 50518 35386
rect 50356 35332 50380 35334
rect 50436 35332 50460 35334
rect 50516 35332 50540 35334
rect 50300 35312 50596 35332
rect 50300 34300 50596 34320
rect 50356 34298 50380 34300
rect 50436 34298 50460 34300
rect 50516 34298 50540 34300
rect 50378 34246 50380 34298
rect 50442 34246 50454 34298
rect 50516 34246 50518 34298
rect 50356 34244 50380 34246
rect 50436 34244 50460 34246
rect 50516 34244 50540 34246
rect 50300 34224 50596 34244
rect 50300 33212 50596 33232
rect 50356 33210 50380 33212
rect 50436 33210 50460 33212
rect 50516 33210 50540 33212
rect 50378 33158 50380 33210
rect 50442 33158 50454 33210
rect 50516 33158 50518 33210
rect 50356 33156 50380 33158
rect 50436 33156 50460 33158
rect 50516 33156 50540 33158
rect 50300 33136 50596 33156
rect 50300 32124 50596 32144
rect 50356 32122 50380 32124
rect 50436 32122 50460 32124
rect 50516 32122 50540 32124
rect 50378 32070 50380 32122
rect 50442 32070 50454 32122
rect 50516 32070 50518 32122
rect 50356 32068 50380 32070
rect 50436 32068 50460 32070
rect 50516 32068 50540 32070
rect 50300 32048 50596 32068
rect 50300 31036 50596 31056
rect 50356 31034 50380 31036
rect 50436 31034 50460 31036
rect 50516 31034 50540 31036
rect 50378 30982 50380 31034
rect 50442 30982 50454 31034
rect 50516 30982 50518 31034
rect 50356 30980 50380 30982
rect 50436 30980 50460 30982
rect 50516 30980 50540 30982
rect 50300 30960 50596 30980
rect 50300 29948 50596 29968
rect 50356 29946 50380 29948
rect 50436 29946 50460 29948
rect 50516 29946 50540 29948
rect 50378 29894 50380 29946
rect 50442 29894 50454 29946
rect 50516 29894 50518 29946
rect 50356 29892 50380 29894
rect 50436 29892 50460 29894
rect 50516 29892 50540 29894
rect 50300 29872 50596 29892
rect 50300 28860 50596 28880
rect 50356 28858 50380 28860
rect 50436 28858 50460 28860
rect 50516 28858 50540 28860
rect 50378 28806 50380 28858
rect 50442 28806 50454 28858
rect 50516 28806 50518 28858
rect 50356 28804 50380 28806
rect 50436 28804 50460 28806
rect 50516 28804 50540 28806
rect 50300 28784 50596 28804
rect 50300 27772 50596 27792
rect 50356 27770 50380 27772
rect 50436 27770 50460 27772
rect 50516 27770 50540 27772
rect 50378 27718 50380 27770
rect 50442 27718 50454 27770
rect 50516 27718 50518 27770
rect 50356 27716 50380 27718
rect 50436 27716 50460 27718
rect 50516 27716 50540 27718
rect 50300 27696 50596 27716
rect 50300 26684 50596 26704
rect 50356 26682 50380 26684
rect 50436 26682 50460 26684
rect 50516 26682 50540 26684
rect 50378 26630 50380 26682
rect 50442 26630 50454 26682
rect 50516 26630 50518 26682
rect 50356 26628 50380 26630
rect 50436 26628 50460 26630
rect 50516 26628 50540 26630
rect 50300 26608 50596 26628
rect 50300 25596 50596 25616
rect 50356 25594 50380 25596
rect 50436 25594 50460 25596
rect 50516 25594 50540 25596
rect 50378 25542 50380 25594
rect 50442 25542 50454 25594
rect 50516 25542 50518 25594
rect 50356 25540 50380 25542
rect 50436 25540 50460 25542
rect 50516 25540 50540 25542
rect 50300 25520 50596 25540
rect 50300 24508 50596 24528
rect 50356 24506 50380 24508
rect 50436 24506 50460 24508
rect 50516 24506 50540 24508
rect 50378 24454 50380 24506
rect 50442 24454 50454 24506
rect 50516 24454 50518 24506
rect 50356 24452 50380 24454
rect 50436 24452 50460 24454
rect 50516 24452 50540 24454
rect 50300 24432 50596 24452
rect 50300 23420 50596 23440
rect 50356 23418 50380 23420
rect 50436 23418 50460 23420
rect 50516 23418 50540 23420
rect 50378 23366 50380 23418
rect 50442 23366 50454 23418
rect 50516 23366 50518 23418
rect 50356 23364 50380 23366
rect 50436 23364 50460 23366
rect 50516 23364 50540 23366
rect 50300 23344 50596 23364
rect 50300 22332 50596 22352
rect 50356 22330 50380 22332
rect 50436 22330 50460 22332
rect 50516 22330 50540 22332
rect 50378 22278 50380 22330
rect 50442 22278 50454 22330
rect 50516 22278 50518 22330
rect 50356 22276 50380 22278
rect 50436 22276 50460 22278
rect 50516 22276 50540 22278
rect 50300 22256 50596 22276
rect 50300 21244 50596 21264
rect 50356 21242 50380 21244
rect 50436 21242 50460 21244
rect 50516 21242 50540 21244
rect 50378 21190 50380 21242
rect 50442 21190 50454 21242
rect 50516 21190 50518 21242
rect 50356 21188 50380 21190
rect 50436 21188 50460 21190
rect 50516 21188 50540 21190
rect 50300 21168 50596 21188
rect 50300 20156 50596 20176
rect 50356 20154 50380 20156
rect 50436 20154 50460 20156
rect 50516 20154 50540 20156
rect 50378 20102 50380 20154
rect 50442 20102 50454 20154
rect 50516 20102 50518 20154
rect 50356 20100 50380 20102
rect 50436 20100 50460 20102
rect 50516 20100 50540 20102
rect 50300 20080 50596 20100
rect 50632 19310 50660 72490
rect 50724 72282 50752 80106
rect 50804 80096 50856 80102
rect 50804 80038 50856 80044
rect 50712 72276 50764 72282
rect 50712 72218 50764 72224
rect 50724 56302 50752 72218
rect 50712 56296 50764 56302
rect 50712 56238 50764 56244
rect 50816 47054 50844 80038
rect 50908 77926 50936 97106
rect 51644 96626 51672 99200
rect 52564 97170 52592 99200
rect 53392 97238 53420 99200
rect 53380 97232 53432 97238
rect 53380 97174 53432 97180
rect 52552 97164 52604 97170
rect 52552 97106 52604 97112
rect 53472 97164 53524 97170
rect 53472 97106 53524 97112
rect 52736 96960 52788 96966
rect 52736 96902 52788 96908
rect 51632 96620 51684 96626
rect 51632 96562 51684 96568
rect 51724 96484 51776 96490
rect 51724 96426 51776 96432
rect 50896 77920 50948 77926
rect 50896 77862 50948 77868
rect 51448 74316 51500 74322
rect 51448 74258 51500 74264
rect 50988 64660 51040 64666
rect 50988 64602 51040 64608
rect 50896 64320 50948 64326
rect 50896 64262 50948 64268
rect 50908 64122 50936 64262
rect 50896 64116 50948 64122
rect 50896 64058 50948 64064
rect 51000 63578 51028 64602
rect 51460 64326 51488 74258
rect 51448 64320 51500 64326
rect 51448 64262 51500 64268
rect 50988 63572 51040 63578
rect 50988 63514 51040 63520
rect 50988 61736 51040 61742
rect 50988 61678 51040 61684
rect 50804 47048 50856 47054
rect 50804 46990 50856 46996
rect 50804 43444 50856 43450
rect 50804 43386 50856 43392
rect 50816 37670 50844 43386
rect 51000 39642 51028 61678
rect 51460 58954 51488 64262
rect 51448 58948 51500 58954
rect 51448 58890 51500 58896
rect 51736 52494 51764 96426
rect 52460 91180 52512 91186
rect 52460 91122 52512 91128
rect 52472 89350 52500 91122
rect 52460 89344 52512 89350
rect 52460 89286 52512 89292
rect 52000 74316 52052 74322
rect 52000 74258 52052 74264
rect 51908 57316 51960 57322
rect 51908 57258 51960 57264
rect 51724 52488 51776 52494
rect 51724 52430 51776 52436
rect 50988 39636 51040 39642
rect 50988 39578 51040 39584
rect 50896 37800 50948 37806
rect 50896 37742 50948 37748
rect 50804 37664 50856 37670
rect 50804 37606 50856 37612
rect 50620 19304 50672 19310
rect 50620 19246 50672 19252
rect 50160 19168 50212 19174
rect 50160 19110 50212 19116
rect 50620 19168 50672 19174
rect 50620 19110 50672 19116
rect 50300 19068 50596 19088
rect 50356 19066 50380 19068
rect 50436 19066 50460 19068
rect 50516 19066 50540 19068
rect 50378 19014 50380 19066
rect 50442 19014 50454 19066
rect 50516 19014 50518 19066
rect 50356 19012 50380 19014
rect 50436 19012 50460 19014
rect 50516 19012 50540 19014
rect 50300 18992 50596 19012
rect 50632 18698 50660 19110
rect 50620 18692 50672 18698
rect 50620 18634 50672 18640
rect 50300 17980 50596 18000
rect 50356 17978 50380 17980
rect 50436 17978 50460 17980
rect 50516 17978 50540 17980
rect 50378 17926 50380 17978
rect 50442 17926 50454 17978
rect 50516 17926 50518 17978
rect 50356 17924 50380 17926
rect 50436 17924 50460 17926
rect 50516 17924 50540 17926
rect 50300 17904 50596 17924
rect 50300 16892 50596 16912
rect 50356 16890 50380 16892
rect 50436 16890 50460 16892
rect 50516 16890 50540 16892
rect 50378 16838 50380 16890
rect 50442 16838 50454 16890
rect 50516 16838 50518 16890
rect 50356 16836 50380 16838
rect 50436 16836 50460 16838
rect 50516 16836 50540 16838
rect 50300 16816 50596 16836
rect 50160 16652 50212 16658
rect 50160 16594 50212 16600
rect 50172 5914 50200 16594
rect 50300 15804 50596 15824
rect 50356 15802 50380 15804
rect 50436 15802 50460 15804
rect 50516 15802 50540 15804
rect 50378 15750 50380 15802
rect 50442 15750 50454 15802
rect 50516 15750 50518 15802
rect 50356 15748 50380 15750
rect 50436 15748 50460 15750
rect 50516 15748 50540 15750
rect 50300 15728 50596 15748
rect 50300 14716 50596 14736
rect 50356 14714 50380 14716
rect 50436 14714 50460 14716
rect 50516 14714 50540 14716
rect 50378 14662 50380 14714
rect 50442 14662 50454 14714
rect 50516 14662 50518 14714
rect 50356 14660 50380 14662
rect 50436 14660 50460 14662
rect 50516 14660 50540 14662
rect 50300 14640 50596 14660
rect 50300 13628 50596 13648
rect 50356 13626 50380 13628
rect 50436 13626 50460 13628
rect 50516 13626 50540 13628
rect 50378 13574 50380 13626
rect 50442 13574 50454 13626
rect 50516 13574 50518 13626
rect 50356 13572 50380 13574
rect 50436 13572 50460 13574
rect 50516 13572 50540 13574
rect 50300 13552 50596 13572
rect 50300 12540 50596 12560
rect 50356 12538 50380 12540
rect 50436 12538 50460 12540
rect 50516 12538 50540 12540
rect 50378 12486 50380 12538
rect 50442 12486 50454 12538
rect 50516 12486 50518 12538
rect 50356 12484 50380 12486
rect 50436 12484 50460 12486
rect 50516 12484 50540 12486
rect 50300 12464 50596 12484
rect 50300 11452 50596 11472
rect 50356 11450 50380 11452
rect 50436 11450 50460 11452
rect 50516 11450 50540 11452
rect 50378 11398 50380 11450
rect 50442 11398 50454 11450
rect 50516 11398 50518 11450
rect 50356 11396 50380 11398
rect 50436 11396 50460 11398
rect 50516 11396 50540 11398
rect 50300 11376 50596 11396
rect 50816 11286 50844 37606
rect 50908 19854 50936 37742
rect 51356 36372 51408 36378
rect 51356 36314 51408 36320
rect 51448 36372 51500 36378
rect 51448 36314 51500 36320
rect 51368 36122 51396 36314
rect 51460 36242 51488 36314
rect 51448 36236 51500 36242
rect 51448 36178 51500 36184
rect 51632 36236 51684 36242
rect 51632 36178 51684 36184
rect 51816 36236 51868 36242
rect 51816 36178 51868 36184
rect 51644 36122 51672 36178
rect 51368 36094 51672 36122
rect 51724 36168 51776 36174
rect 51724 36110 51776 36116
rect 51736 35222 51764 36110
rect 51724 35216 51776 35222
rect 51724 35158 51776 35164
rect 51736 34610 51764 35158
rect 51828 34678 51856 36178
rect 51920 36174 51948 57258
rect 52012 48142 52040 74258
rect 52460 74248 52512 74254
rect 52460 74190 52512 74196
rect 52092 74112 52144 74118
rect 52092 74054 52144 74060
rect 52104 73846 52132 74054
rect 52092 73840 52144 73846
rect 52092 73782 52144 73788
rect 52368 67176 52420 67182
rect 52368 67118 52420 67124
rect 52276 52488 52328 52494
rect 52276 52430 52328 52436
rect 52000 48136 52052 48142
rect 52000 48078 52052 48084
rect 51908 36168 51960 36174
rect 51908 36110 51960 36116
rect 51816 34672 51868 34678
rect 51816 34614 51868 34620
rect 51724 34604 51776 34610
rect 51724 34546 51776 34552
rect 51828 28994 51856 34614
rect 51828 28966 51948 28994
rect 51920 27538 51948 28966
rect 51908 27532 51960 27538
rect 51908 27474 51960 27480
rect 50896 19848 50948 19854
rect 50896 19790 50948 19796
rect 51264 18080 51316 18086
rect 51264 18022 51316 18028
rect 51080 11620 51132 11626
rect 51080 11562 51132 11568
rect 50804 11280 50856 11286
rect 50804 11222 50856 11228
rect 51092 11014 51120 11562
rect 51080 11008 51132 11014
rect 51080 10950 51132 10956
rect 50300 10364 50596 10384
rect 50356 10362 50380 10364
rect 50436 10362 50460 10364
rect 50516 10362 50540 10364
rect 50378 10310 50380 10362
rect 50442 10310 50454 10362
rect 50516 10310 50518 10362
rect 50356 10308 50380 10310
rect 50436 10308 50460 10310
rect 50516 10308 50540 10310
rect 50300 10288 50596 10308
rect 50300 9276 50596 9296
rect 50356 9274 50380 9276
rect 50436 9274 50460 9276
rect 50516 9274 50540 9276
rect 50378 9222 50380 9274
rect 50442 9222 50454 9274
rect 50516 9222 50518 9274
rect 50356 9220 50380 9222
rect 50436 9220 50460 9222
rect 50516 9220 50540 9222
rect 50300 9200 50596 9220
rect 50712 8356 50764 8362
rect 50712 8298 50764 8304
rect 50300 8188 50596 8208
rect 50356 8186 50380 8188
rect 50436 8186 50460 8188
rect 50516 8186 50540 8188
rect 50378 8134 50380 8186
rect 50442 8134 50454 8186
rect 50516 8134 50518 8186
rect 50356 8132 50380 8134
rect 50436 8132 50460 8134
rect 50516 8132 50540 8134
rect 50300 8112 50596 8132
rect 50300 7100 50596 7120
rect 50356 7098 50380 7100
rect 50436 7098 50460 7100
rect 50516 7098 50540 7100
rect 50378 7046 50380 7098
rect 50442 7046 50454 7098
rect 50516 7046 50518 7098
rect 50356 7044 50380 7046
rect 50436 7044 50460 7046
rect 50516 7044 50540 7046
rect 50300 7024 50596 7044
rect 50300 6012 50596 6032
rect 50356 6010 50380 6012
rect 50436 6010 50460 6012
rect 50516 6010 50540 6012
rect 50378 5958 50380 6010
rect 50442 5958 50454 6010
rect 50516 5958 50518 6010
rect 50356 5956 50380 5958
rect 50436 5956 50460 5958
rect 50516 5956 50540 5958
rect 50300 5936 50596 5956
rect 50160 5908 50212 5914
rect 50160 5850 50212 5856
rect 50068 5840 50120 5846
rect 50068 5782 50120 5788
rect 50300 4924 50596 4944
rect 50356 4922 50380 4924
rect 50436 4922 50460 4924
rect 50516 4922 50540 4924
rect 50378 4870 50380 4922
rect 50442 4870 50454 4922
rect 50516 4870 50518 4922
rect 50356 4868 50380 4870
rect 50436 4868 50460 4870
rect 50516 4868 50540 4870
rect 50300 4848 50596 4868
rect 50160 4072 50212 4078
rect 50080 4032 50160 4060
rect 49884 2508 49936 2514
rect 49884 2450 49936 2456
rect 49792 1352 49844 1358
rect 49792 1294 49844 1300
rect 49896 800 49924 2450
rect 50080 800 50108 4032
rect 50160 4014 50212 4020
rect 50300 3836 50596 3856
rect 50356 3834 50380 3836
rect 50436 3834 50460 3836
rect 50516 3834 50540 3836
rect 50378 3782 50380 3834
rect 50442 3782 50454 3834
rect 50516 3782 50518 3834
rect 50356 3780 50380 3782
rect 50436 3780 50460 3782
rect 50516 3780 50540 3782
rect 50300 3760 50596 3780
rect 50160 2848 50212 2854
rect 50160 2790 50212 2796
rect 50172 1442 50200 2790
rect 50300 2748 50596 2768
rect 50356 2746 50380 2748
rect 50436 2746 50460 2748
rect 50516 2746 50540 2748
rect 50378 2694 50380 2746
rect 50442 2694 50454 2746
rect 50516 2694 50518 2746
rect 50356 2692 50380 2694
rect 50436 2692 50460 2694
rect 50516 2692 50540 2694
rect 50300 2672 50596 2692
rect 50724 2650 50752 8298
rect 50988 7880 51040 7886
rect 50988 7822 51040 7828
rect 50804 4072 50856 4078
rect 50804 4014 50856 4020
rect 50712 2644 50764 2650
rect 50712 2586 50764 2592
rect 50528 2304 50580 2310
rect 50528 2246 50580 2252
rect 50172 1414 50292 1442
rect 50264 800 50292 1414
rect 50540 1170 50568 2246
rect 50816 1442 50844 4014
rect 50896 3596 50948 3602
rect 50896 3538 50948 3544
rect 50448 1142 50568 1170
rect 50724 1414 50844 1442
rect 50448 800 50476 1142
rect 50724 800 50752 1414
rect 50908 800 50936 3538
rect 51000 2582 51028 7822
rect 51276 2990 51304 18022
rect 52012 11626 52040 48078
rect 52184 43444 52236 43450
rect 52184 43386 52236 43392
rect 52196 36242 52224 43386
rect 52184 36236 52236 36242
rect 52184 36178 52236 36184
rect 52288 24206 52316 52430
rect 52380 37466 52408 67118
rect 52472 64054 52500 74190
rect 52644 67108 52696 67114
rect 52644 67050 52696 67056
rect 52552 67040 52604 67046
rect 52552 66982 52604 66988
rect 52564 65618 52592 66982
rect 52552 65612 52604 65618
rect 52552 65554 52604 65560
rect 52460 64048 52512 64054
rect 52460 63990 52512 63996
rect 52552 61260 52604 61266
rect 52552 61202 52604 61208
rect 52564 60858 52592 61202
rect 52552 60852 52604 60858
rect 52552 60794 52604 60800
rect 52656 52086 52684 67050
rect 52748 60654 52776 96902
rect 53196 89344 53248 89350
rect 53196 89286 53248 89292
rect 53012 64048 53064 64054
rect 53012 63990 53064 63996
rect 52920 61396 52972 61402
rect 52920 61338 52972 61344
rect 52932 61266 52960 61338
rect 52920 61260 52972 61266
rect 52920 61202 52972 61208
rect 52736 60648 52788 60654
rect 52736 60590 52788 60596
rect 53024 54602 53052 63990
rect 53104 63232 53156 63238
rect 53104 63174 53156 63180
rect 53012 54596 53064 54602
rect 53012 54538 53064 54544
rect 52644 52080 52696 52086
rect 52644 52022 52696 52028
rect 52460 48612 52512 48618
rect 52460 48554 52512 48560
rect 52472 48210 52500 48554
rect 52460 48204 52512 48210
rect 52460 48146 52512 48152
rect 52368 37460 52420 37466
rect 52368 37402 52420 37408
rect 52380 36786 52408 37402
rect 52368 36780 52420 36786
rect 52368 36722 52420 36728
rect 52276 24200 52328 24206
rect 52276 24142 52328 24148
rect 52000 11620 52052 11626
rect 52000 11562 52052 11568
rect 53116 9586 53144 63174
rect 53208 48210 53236 89286
rect 53288 74452 53340 74458
rect 53288 74394 53340 74400
rect 53300 71126 53328 74394
rect 53380 74384 53432 74390
rect 53380 74326 53432 74332
rect 53288 71120 53340 71126
rect 53288 71062 53340 71068
rect 53392 71058 53420 74326
rect 53380 71052 53432 71058
rect 53380 70994 53432 71000
rect 53288 66496 53340 66502
rect 53288 66438 53340 66444
rect 53196 48204 53248 48210
rect 53196 48146 53248 48152
rect 53300 18086 53328 66438
rect 53380 56228 53432 56234
rect 53380 56170 53432 56176
rect 53392 53718 53420 56170
rect 53380 53712 53432 53718
rect 53380 53654 53432 53660
rect 53380 50448 53432 50454
rect 53380 50390 53432 50396
rect 53392 18902 53420 50390
rect 53484 28762 53512 97106
rect 54312 96626 54340 99200
rect 55140 97170 55168 99200
rect 55968 97238 55996 99200
rect 56508 97572 56560 97578
rect 56508 97514 56560 97520
rect 55956 97232 56008 97238
rect 55956 97174 56008 97180
rect 55128 97164 55180 97170
rect 55128 97106 55180 97112
rect 56416 97164 56468 97170
rect 56416 97106 56468 97112
rect 54300 96620 54352 96626
rect 54300 96562 54352 96568
rect 54392 96484 54444 96490
rect 54392 96426 54444 96432
rect 53840 95600 53892 95606
rect 53840 95542 53892 95548
rect 53748 89140 53800 89146
rect 53748 89082 53800 89088
rect 53656 77920 53708 77926
rect 53656 77862 53708 77868
rect 53564 65612 53616 65618
rect 53564 65554 53616 65560
rect 53576 62422 53604 65554
rect 53564 62416 53616 62422
rect 53564 62358 53616 62364
rect 53564 59084 53616 59090
rect 53564 59026 53616 59032
rect 53576 46170 53604 59026
rect 53668 52698 53696 77862
rect 53760 56846 53788 89082
rect 53852 82482 53880 95542
rect 53932 94852 53984 94858
rect 53932 94794 53984 94800
rect 53944 85270 53972 94794
rect 53932 85264 53984 85270
rect 53932 85206 53984 85212
rect 53840 82476 53892 82482
rect 53840 82418 53892 82424
rect 54300 81864 54352 81870
rect 54300 81806 54352 81812
rect 54208 61804 54260 61810
rect 54208 61746 54260 61752
rect 53748 56840 53800 56846
rect 53748 56782 53800 56788
rect 53656 52692 53708 52698
rect 53656 52634 53708 52640
rect 53564 46164 53616 46170
rect 53564 46106 53616 46112
rect 53668 43178 53696 52634
rect 53760 50454 53788 56782
rect 54220 56302 54248 61746
rect 54208 56296 54260 56302
rect 54208 56238 54260 56244
rect 53840 54664 53892 54670
rect 53840 54606 53892 54612
rect 53852 53718 53880 54606
rect 53840 53712 53892 53718
rect 53840 53654 53892 53660
rect 53748 50448 53800 50454
rect 53748 50390 53800 50396
rect 53748 49156 53800 49162
rect 53748 49098 53800 49104
rect 53760 44198 53788 49098
rect 53748 44192 53800 44198
rect 53748 44134 53800 44140
rect 53656 43172 53708 43178
rect 53656 43114 53708 43120
rect 53748 40928 53800 40934
rect 53748 40870 53800 40876
rect 53656 40180 53708 40186
rect 53656 40122 53708 40128
rect 53564 34740 53616 34746
rect 53564 34682 53616 34688
rect 53472 28756 53524 28762
rect 53472 28698 53524 28704
rect 53380 18896 53432 18902
rect 53380 18838 53432 18844
rect 53288 18080 53340 18086
rect 53288 18022 53340 18028
rect 53196 11076 53248 11082
rect 53196 11018 53248 11024
rect 53104 9580 53156 9586
rect 53104 9522 53156 9528
rect 53208 9110 53236 11018
rect 53196 9104 53248 9110
rect 53196 9046 53248 9052
rect 53576 6730 53604 34682
rect 53564 6724 53616 6730
rect 53564 6666 53616 6672
rect 52460 6248 52512 6254
rect 52460 6190 52512 6196
rect 52472 5030 52500 6190
rect 53576 6186 53604 6666
rect 53564 6180 53616 6186
rect 53564 6122 53616 6128
rect 52460 5024 52512 5030
rect 52460 4966 52512 4972
rect 52552 4684 52604 4690
rect 52552 4626 52604 4632
rect 53104 4684 53156 4690
rect 53104 4626 53156 4632
rect 51448 4072 51500 4078
rect 51368 4032 51448 4060
rect 51264 2984 51316 2990
rect 51264 2926 51316 2932
rect 51080 2916 51132 2922
rect 51080 2858 51132 2864
rect 50988 2576 51040 2582
rect 50988 2518 51040 2524
rect 51092 800 51120 2858
rect 51368 2122 51396 4032
rect 51448 4014 51500 4020
rect 51908 4004 51960 4010
rect 51908 3946 51960 3952
rect 51448 2916 51500 2922
rect 51448 2858 51500 2864
rect 51276 2094 51396 2122
rect 51276 800 51304 2094
rect 51460 800 51488 2858
rect 51724 2440 51776 2446
rect 51724 2382 51776 2388
rect 51540 2304 51592 2310
rect 51540 2246 51592 2252
rect 51552 2106 51580 2246
rect 51540 2100 51592 2106
rect 51540 2042 51592 2048
rect 51736 800 51764 2382
rect 51920 800 51948 3946
rect 52092 3596 52144 3602
rect 52092 3538 52144 3544
rect 52104 800 52132 3538
rect 52368 3052 52420 3058
rect 52368 2994 52420 3000
rect 52380 2582 52408 2994
rect 52368 2576 52420 2582
rect 52368 2518 52420 2524
rect 52276 2100 52328 2106
rect 52276 2042 52328 2048
rect 52288 800 52316 2042
rect 52564 800 52592 4626
rect 52736 3596 52788 3602
rect 52736 3538 52788 3544
rect 52748 800 52776 3538
rect 52920 2372 52972 2378
rect 52920 2314 52972 2320
rect 52932 800 52960 2314
rect 53116 800 53144 4626
rect 53288 3596 53340 3602
rect 53288 3538 53340 3544
rect 53300 800 53328 3538
rect 53564 2848 53616 2854
rect 53564 2790 53616 2796
rect 53576 800 53604 2790
rect 53668 2582 53696 40122
rect 53760 39574 53788 40870
rect 53748 39568 53800 39574
rect 53748 39510 53800 39516
rect 53852 31346 53880 53654
rect 54024 53644 54076 53650
rect 54024 53586 54076 53592
rect 54036 53514 54064 53586
rect 54024 53508 54076 53514
rect 54024 53450 54076 53456
rect 54036 53174 54064 53450
rect 54208 53440 54260 53446
rect 54208 53382 54260 53388
rect 54024 53168 54076 53174
rect 54024 53110 54076 53116
rect 53840 31340 53892 31346
rect 53840 31282 53892 31288
rect 54220 24818 54248 53382
rect 54208 24812 54260 24818
rect 54208 24754 54260 24760
rect 54116 19168 54168 19174
rect 54116 19110 54168 19116
rect 53840 11756 53892 11762
rect 53840 11698 53892 11704
rect 53852 11218 53880 11698
rect 53840 11212 53892 11218
rect 53840 11154 53892 11160
rect 53840 6452 53892 6458
rect 53840 6394 53892 6400
rect 53748 4072 53800 4078
rect 53748 4014 53800 4020
rect 53656 2576 53708 2582
rect 53656 2518 53708 2524
rect 53760 800 53788 4014
rect 53852 2582 53880 6394
rect 53932 3596 53984 3602
rect 53932 3538 53984 3544
rect 53840 2576 53892 2582
rect 53840 2518 53892 2524
rect 53944 800 53972 3538
rect 54128 2990 54156 19110
rect 54312 11218 54340 81806
rect 54404 60314 54432 96426
rect 56428 94994 56456 97106
rect 56520 95946 56548 97514
rect 56888 96626 56916 99200
rect 57716 97238 57744 99200
rect 58636 97238 58664 99200
rect 57704 97232 57756 97238
rect 57704 97174 57756 97180
rect 58624 97232 58676 97238
rect 58624 97174 58676 97180
rect 57980 97028 58032 97034
rect 57980 96970 58032 96976
rect 56876 96620 56928 96626
rect 56876 96562 56928 96568
rect 56968 96484 57020 96490
rect 56968 96426 57020 96432
rect 56508 95940 56560 95946
rect 56508 95882 56560 95888
rect 55404 94988 55456 94994
rect 55404 94930 55456 94936
rect 56416 94988 56468 94994
rect 56416 94930 56468 94936
rect 54576 94920 54628 94926
rect 54576 94862 54628 94868
rect 54484 87712 54536 87718
rect 54484 87654 54536 87660
rect 54496 81870 54524 87654
rect 54484 81864 54536 81870
rect 54484 81806 54536 81812
rect 54484 76968 54536 76974
rect 54484 76910 54536 76916
rect 54496 75410 54524 76910
rect 54484 75404 54536 75410
rect 54484 75346 54536 75352
rect 54392 60308 54444 60314
rect 54392 60250 54444 60256
rect 54484 60104 54536 60110
rect 54484 60046 54536 60052
rect 54496 59498 54524 60046
rect 54484 59492 54536 59498
rect 54484 59434 54536 59440
rect 54484 56296 54536 56302
rect 54484 56238 54536 56244
rect 54392 53508 54444 53514
rect 54392 53450 54444 53456
rect 54404 52562 54432 53450
rect 54392 52556 54444 52562
rect 54392 52498 54444 52504
rect 54496 14278 54524 56238
rect 54588 52154 54616 94862
rect 55036 91112 55088 91118
rect 55036 91054 55088 91060
rect 55048 88942 55076 91054
rect 55036 88936 55088 88942
rect 55036 88878 55088 88884
rect 54668 86352 54720 86358
rect 54668 86294 54720 86300
rect 54576 52148 54628 52154
rect 54576 52090 54628 52096
rect 54588 51950 54616 52090
rect 54576 51944 54628 51950
rect 54576 51886 54628 51892
rect 54680 34746 54708 86294
rect 55312 72140 55364 72146
rect 55312 72082 55364 72088
rect 55220 72004 55272 72010
rect 55220 71946 55272 71952
rect 54852 71936 54904 71942
rect 54852 71878 54904 71884
rect 54864 63918 54892 71878
rect 55232 70378 55260 71946
rect 55220 70372 55272 70378
rect 55220 70314 55272 70320
rect 55232 69902 55260 70314
rect 55220 69896 55272 69902
rect 55220 69838 55272 69844
rect 55324 64530 55352 72082
rect 55312 64524 55364 64530
rect 55312 64466 55364 64472
rect 54852 63912 54904 63918
rect 54852 63854 54904 63860
rect 54852 60580 54904 60586
rect 54852 60522 54904 60528
rect 54760 60308 54812 60314
rect 54760 60250 54812 60256
rect 54772 47666 54800 60250
rect 54864 59634 54892 60522
rect 54852 59628 54904 59634
rect 54852 59570 54904 59576
rect 55128 51876 55180 51882
rect 55128 51818 55180 51824
rect 54760 47660 54812 47666
rect 54760 47602 54812 47608
rect 54760 44872 54812 44878
rect 54760 44814 54812 44820
rect 54668 34740 54720 34746
rect 54668 34682 54720 34688
rect 54484 14272 54536 14278
rect 54484 14214 54536 14220
rect 54300 11212 54352 11218
rect 54300 11154 54352 11160
rect 54312 10606 54340 11154
rect 54300 10600 54352 10606
rect 54300 10542 54352 10548
rect 54300 4072 54352 4078
rect 54300 4014 54352 4020
rect 54116 2984 54168 2990
rect 54116 2926 54168 2932
rect 54116 2508 54168 2514
rect 54116 2450 54168 2456
rect 54128 800 54156 2450
rect 54312 800 54340 4014
rect 54576 3596 54628 3602
rect 54576 3538 54628 3544
rect 54588 800 54616 3538
rect 54772 2650 54800 44814
rect 55140 43110 55168 51818
rect 55416 49162 55444 94930
rect 55588 76628 55640 76634
rect 55588 76570 55640 76576
rect 56232 76628 56284 76634
rect 56232 76570 56284 76576
rect 55496 56160 55548 56166
rect 55496 56102 55548 56108
rect 55404 49156 55456 49162
rect 55404 49098 55456 49104
rect 55128 43104 55180 43110
rect 55128 43046 55180 43052
rect 55508 39506 55536 56102
rect 55496 39500 55548 39506
rect 55496 39442 55548 39448
rect 55036 20392 55088 20398
rect 55036 20334 55088 20340
rect 55048 18766 55076 20334
rect 55036 18760 55088 18766
rect 55036 18702 55088 18708
rect 55048 18222 55076 18702
rect 55036 18216 55088 18222
rect 55036 18158 55088 18164
rect 55312 18216 55364 18222
rect 55312 18158 55364 18164
rect 55324 17066 55352 18158
rect 55312 17060 55364 17066
rect 55312 17002 55364 17008
rect 55220 14884 55272 14890
rect 55220 14826 55272 14832
rect 55232 14278 55260 14826
rect 55220 14272 55272 14278
rect 55220 14214 55272 14220
rect 55036 11144 55088 11150
rect 55036 11086 55088 11092
rect 55048 10606 55076 11086
rect 55232 11082 55260 14214
rect 55220 11076 55272 11082
rect 55220 11018 55272 11024
rect 55232 10962 55260 11018
rect 55232 10934 55352 10962
rect 55220 10804 55272 10810
rect 55220 10746 55272 10752
rect 55036 10600 55088 10606
rect 55036 10542 55088 10548
rect 54944 4072 54996 4078
rect 54944 4014 54996 4020
rect 54852 3052 54904 3058
rect 54852 2994 54904 3000
rect 54760 2644 54812 2650
rect 54760 2586 54812 2592
rect 54864 1578 54892 2994
rect 54772 1550 54892 1578
rect 54772 800 54800 1550
rect 54956 800 54984 4014
rect 55128 3596 55180 3602
rect 55128 3538 55180 3544
rect 55036 2440 55088 2446
rect 55036 2382 55088 2388
rect 55048 2106 55076 2382
rect 55036 2100 55088 2106
rect 55036 2042 55088 2048
rect 55140 800 55168 3538
rect 55232 3194 55260 10746
rect 55324 10606 55352 10934
rect 55600 10606 55628 76570
rect 56244 76090 56272 76570
rect 56232 76084 56284 76090
rect 56232 76026 56284 76032
rect 56048 64524 56100 64530
rect 56048 64466 56100 64472
rect 55772 59424 55824 59430
rect 55772 59366 55824 59372
rect 55784 28014 55812 59366
rect 55864 57928 55916 57934
rect 55864 57870 55916 57876
rect 55772 28008 55824 28014
rect 55772 27950 55824 27956
rect 55772 15156 55824 15162
rect 55772 15098 55824 15104
rect 55312 10600 55364 10606
rect 55312 10542 55364 10548
rect 55588 10600 55640 10606
rect 55588 10542 55640 10548
rect 55600 9518 55628 10542
rect 55588 9512 55640 9518
rect 55588 9454 55640 9460
rect 55588 4072 55640 4078
rect 55588 4014 55640 4020
rect 55220 3188 55272 3194
rect 55220 3130 55272 3136
rect 55232 2990 55260 3130
rect 55220 2984 55272 2990
rect 55220 2926 55272 2932
rect 55312 2916 55364 2922
rect 55312 2858 55364 2864
rect 55324 800 55352 2858
rect 55600 800 55628 4014
rect 55784 2582 55812 15098
rect 55876 4554 55904 57870
rect 56060 50998 56088 64466
rect 56520 57934 56548 95882
rect 56980 85202 57008 96426
rect 57428 96076 57480 96082
rect 57428 96018 57480 96024
rect 57796 96076 57848 96082
rect 57796 96018 57848 96024
rect 56968 85196 57020 85202
rect 56968 85138 57020 85144
rect 56692 76424 56744 76430
rect 56692 76366 56744 76372
rect 56704 74322 56732 76366
rect 56692 74316 56744 74322
rect 56692 74258 56744 74264
rect 56968 74248 57020 74254
rect 56968 74190 57020 74196
rect 56980 73914 57008 74190
rect 56968 73908 57020 73914
rect 56968 73850 57020 73856
rect 57244 70440 57296 70446
rect 57440 70417 57468 96018
rect 57612 96008 57664 96014
rect 57612 95950 57664 95956
rect 57520 75472 57572 75478
rect 57520 75414 57572 75420
rect 57244 70382 57296 70388
rect 57426 70408 57482 70417
rect 56968 67040 57020 67046
rect 56968 66982 57020 66988
rect 56980 60110 57008 66982
rect 57060 63368 57112 63374
rect 57060 63310 57112 63316
rect 57072 60586 57100 63310
rect 57060 60580 57112 60586
rect 57060 60522 57112 60528
rect 56968 60104 57020 60110
rect 56968 60046 57020 60052
rect 57152 59628 57204 59634
rect 57152 59570 57204 59576
rect 57060 58540 57112 58546
rect 57060 58482 57112 58488
rect 56508 57928 56560 57934
rect 56508 57870 56560 57876
rect 56520 57322 56548 57870
rect 56508 57316 56560 57322
rect 56508 57258 56560 57264
rect 56600 55412 56652 55418
rect 56600 55354 56652 55360
rect 56048 50992 56100 50998
rect 56048 50934 56100 50940
rect 55956 49768 56008 49774
rect 55956 49710 56008 49716
rect 55968 42634 55996 49710
rect 56060 43178 56088 50934
rect 56048 43172 56100 43178
rect 56048 43114 56100 43120
rect 55956 42628 56008 42634
rect 55956 42570 56008 42576
rect 55968 28082 55996 42570
rect 56612 34202 56640 55354
rect 56600 34196 56652 34202
rect 56600 34138 56652 34144
rect 57072 34066 57100 58482
rect 57060 34060 57112 34066
rect 57060 34002 57112 34008
rect 56968 33992 57020 33998
rect 56968 33934 57020 33940
rect 56980 33522 57008 33934
rect 56968 33516 57020 33522
rect 56968 33458 57020 33464
rect 56048 32768 56100 32774
rect 56048 32710 56100 32716
rect 55956 28076 56008 28082
rect 55956 28018 56008 28024
rect 55956 18624 56008 18630
rect 55956 18566 56008 18572
rect 55968 18290 55996 18566
rect 55956 18284 56008 18290
rect 55956 18226 56008 18232
rect 55956 12980 56008 12986
rect 55956 12922 56008 12928
rect 55968 12850 55996 12922
rect 55956 12844 56008 12850
rect 55956 12786 56008 12792
rect 56060 9110 56088 32710
rect 56232 28008 56284 28014
rect 56152 27956 56232 27962
rect 56152 27950 56284 27956
rect 56152 27934 56272 27950
rect 56152 21418 56180 27934
rect 56232 27872 56284 27878
rect 56232 27814 56284 27820
rect 56244 27674 56272 27814
rect 56232 27668 56284 27674
rect 56232 27610 56284 27616
rect 56600 27328 56652 27334
rect 56600 27270 56652 27276
rect 56612 22094 56640 27270
rect 57072 26926 57100 34002
rect 57060 26920 57112 26926
rect 57060 26862 57112 26868
rect 56784 25764 56836 25770
rect 56784 25706 56836 25712
rect 56796 22094 56824 25706
rect 56612 22066 56732 22094
rect 56796 22066 56916 22094
rect 56140 21412 56192 21418
rect 56140 21354 56192 21360
rect 56152 19786 56180 21354
rect 56140 19780 56192 19786
rect 56140 19722 56192 19728
rect 56140 12912 56192 12918
rect 56140 12854 56192 12860
rect 56152 12782 56180 12854
rect 56140 12776 56192 12782
rect 56140 12718 56192 12724
rect 56048 9104 56100 9110
rect 56048 9046 56100 9052
rect 55864 4548 55916 4554
rect 55864 4490 55916 4496
rect 56140 4072 56192 4078
rect 56140 4014 56192 4020
rect 55864 2848 55916 2854
rect 55864 2790 55916 2796
rect 55772 2576 55824 2582
rect 55772 2518 55824 2524
rect 55876 1578 55904 2790
rect 55956 2304 56008 2310
rect 55956 2246 56008 2252
rect 55784 1550 55904 1578
rect 55784 800 55812 1550
rect 55968 800 55996 2246
rect 56152 800 56180 4014
rect 56324 3596 56376 3602
rect 56324 3538 56376 3544
rect 56336 800 56364 3538
rect 56600 2916 56652 2922
rect 56600 2858 56652 2864
rect 56612 800 56640 2858
rect 56704 2582 56732 22066
rect 56784 4072 56836 4078
rect 56784 4014 56836 4020
rect 56692 2576 56744 2582
rect 56692 2518 56744 2524
rect 56796 800 56824 4014
rect 56888 2990 56916 22066
rect 57164 21350 57192 59570
rect 57152 21344 57204 21350
rect 57152 21286 57204 21292
rect 57256 14346 57284 70382
rect 57426 70343 57482 70352
rect 57336 62960 57388 62966
rect 57336 62902 57388 62908
rect 57348 39982 57376 62902
rect 57532 61946 57560 75414
rect 57520 61940 57572 61946
rect 57520 61882 57572 61888
rect 57428 61804 57480 61810
rect 57428 61746 57480 61752
rect 57440 61606 57468 61746
rect 57428 61600 57480 61606
rect 57428 61542 57480 61548
rect 57440 61266 57468 61542
rect 57428 61260 57480 61266
rect 57428 61202 57480 61208
rect 57532 60734 57560 61882
rect 57440 60706 57560 60734
rect 57440 58546 57468 60706
rect 57428 58540 57480 58546
rect 57428 58482 57480 58488
rect 57520 53032 57572 53038
rect 57520 52974 57572 52980
rect 57532 52630 57560 52974
rect 57520 52624 57572 52630
rect 57520 52566 57572 52572
rect 57428 48000 57480 48006
rect 57428 47942 57480 47948
rect 57440 47802 57468 47942
rect 57428 47796 57480 47802
rect 57428 47738 57480 47744
rect 57336 39976 57388 39982
rect 57336 39918 57388 39924
rect 57336 37732 57388 37738
rect 57336 37674 57388 37680
rect 57348 36786 57376 37674
rect 57336 36780 57388 36786
rect 57336 36722 57388 36728
rect 57336 35828 57388 35834
rect 57336 35770 57388 35776
rect 57348 34746 57376 35770
rect 57336 34740 57388 34746
rect 57336 34682 57388 34688
rect 57348 25974 57376 34682
rect 57428 33856 57480 33862
rect 57428 33798 57480 33804
rect 57336 25968 57388 25974
rect 57336 25910 57388 25916
rect 57440 18834 57468 33798
rect 57532 22642 57560 52566
rect 57624 35834 57652 95950
rect 57808 63374 57836 96018
rect 57992 95538 58020 96970
rect 59464 96626 59492 99200
rect 60384 97238 60412 99200
rect 61212 97238 61240 99200
rect 60372 97232 60424 97238
rect 60372 97174 60424 97180
rect 61200 97232 61252 97238
rect 61200 97174 61252 97180
rect 61384 97164 61436 97170
rect 61384 97106 61436 97112
rect 60740 96960 60792 96966
rect 60740 96902 60792 96908
rect 59452 96620 59504 96626
rect 59452 96562 59504 96568
rect 59544 96484 59596 96490
rect 59544 96426 59596 96432
rect 58164 96076 58216 96082
rect 58164 96018 58216 96024
rect 57980 95532 58032 95538
rect 57980 95474 58032 95480
rect 58072 93288 58124 93294
rect 58072 93230 58124 93236
rect 58084 76634 58112 93230
rect 58072 76628 58124 76634
rect 58072 76570 58124 76576
rect 57886 70408 57942 70417
rect 57886 70343 57942 70352
rect 57900 67046 57928 70343
rect 57888 67040 57940 67046
rect 57888 66982 57940 66988
rect 57796 63368 57848 63374
rect 57796 63310 57848 63316
rect 57934 61192 57986 61198
rect 57934 61134 57986 61140
rect 57946 61010 57974 61134
rect 57808 60982 57974 61010
rect 57808 59634 57836 60982
rect 57796 59628 57848 59634
rect 57796 59570 57848 59576
rect 58176 59566 58204 96018
rect 58532 95940 58584 95946
rect 58532 95882 58584 95888
rect 58348 76628 58400 76634
rect 58348 76570 58400 76576
rect 58164 59560 58216 59566
rect 58164 59502 58216 59508
rect 58164 58472 58216 58478
rect 58164 58414 58216 58420
rect 57704 53032 57756 53038
rect 57704 52974 57756 52980
rect 57980 53032 58032 53038
rect 57980 52974 58032 52980
rect 57716 37738 57744 52974
rect 57992 52698 58020 52974
rect 57980 52692 58032 52698
rect 57980 52634 58032 52640
rect 57888 48204 57940 48210
rect 57888 48146 57940 48152
rect 58072 48204 58124 48210
rect 58072 48146 58124 48152
rect 57900 47734 57928 48146
rect 57888 47728 57940 47734
rect 57888 47670 57940 47676
rect 57900 45286 57928 47670
rect 58084 45554 58112 48146
rect 57992 45526 58112 45554
rect 57888 45280 57940 45286
rect 57888 45222 57940 45228
rect 57992 44946 58020 45526
rect 57980 44940 58032 44946
rect 57980 44882 58032 44888
rect 57704 37732 57756 37738
rect 57704 37674 57756 37680
rect 57612 35828 57664 35834
rect 57612 35770 57664 35776
rect 57796 33992 57848 33998
rect 57796 33934 57848 33940
rect 57520 22636 57572 22642
rect 57520 22578 57572 22584
rect 57428 18828 57480 18834
rect 57428 18770 57480 18776
rect 57244 14340 57296 14346
rect 57244 14282 57296 14288
rect 56968 6656 57020 6662
rect 56968 6598 57020 6604
rect 56980 5098 57008 6598
rect 56968 5092 57020 5098
rect 56968 5034 57020 5040
rect 57428 4072 57480 4078
rect 57428 4014 57480 4020
rect 56968 3596 57020 3602
rect 56968 3538 57020 3544
rect 56876 2984 56928 2990
rect 56876 2926 56928 2932
rect 56980 800 57008 3538
rect 57152 3120 57204 3126
rect 57152 3062 57204 3068
rect 57164 800 57192 3062
rect 57440 800 57468 4014
rect 57612 2984 57664 2990
rect 57612 2926 57664 2932
rect 57624 800 57652 2926
rect 57808 2582 57836 33934
rect 57992 15638 58020 44882
rect 58072 32972 58124 32978
rect 58072 32914 58124 32920
rect 58084 15706 58112 32914
rect 58176 30190 58204 58414
rect 58256 54664 58308 54670
rect 58256 54606 58308 54612
rect 58268 53174 58296 54606
rect 58256 53168 58308 53174
rect 58256 53110 58308 53116
rect 58256 48272 58308 48278
rect 58256 48214 58308 48220
rect 58268 48006 58296 48214
rect 58256 48000 58308 48006
rect 58256 47942 58308 47948
rect 58164 30184 58216 30190
rect 58164 30126 58216 30132
rect 58268 18358 58296 47942
rect 58360 43110 58388 76570
rect 58348 43104 58400 43110
rect 58348 43046 58400 43052
rect 58256 18352 58308 18358
rect 58256 18294 58308 18300
rect 58072 15700 58124 15706
rect 58072 15642 58124 15648
rect 57980 15632 58032 15638
rect 57980 15574 58032 15580
rect 58072 9580 58124 9586
rect 58072 9522 58124 9528
rect 57980 3528 58032 3534
rect 57980 3470 58032 3476
rect 57796 2576 57848 2582
rect 57796 2518 57848 2524
rect 57796 2372 57848 2378
rect 57796 2314 57848 2320
rect 57808 800 57836 2314
rect 57992 800 58020 3470
rect 58084 2650 58112 9522
rect 58544 4622 58572 95882
rect 59556 93226 59584 96426
rect 60096 96212 60148 96218
rect 60096 96154 60148 96160
rect 60108 93854 60136 96154
rect 60108 93826 60412 93854
rect 59544 93220 59596 93226
rect 59544 93162 59596 93168
rect 59556 92614 59584 93162
rect 59544 92608 59596 92614
rect 59544 92550 59596 92556
rect 59912 87372 59964 87378
rect 59912 87314 59964 87320
rect 59924 87174 59952 87314
rect 59912 87168 59964 87174
rect 59912 87110 59964 87116
rect 60384 84046 60412 93826
rect 60556 92608 60608 92614
rect 60556 92550 60608 92556
rect 60372 84040 60424 84046
rect 60372 83982 60424 83988
rect 58624 78192 58676 78198
rect 58624 78134 58676 78140
rect 58636 61946 58664 78134
rect 60384 74534 60412 83982
rect 60200 74506 60412 74534
rect 59912 72548 59964 72554
rect 59912 72490 59964 72496
rect 59924 72146 59952 72490
rect 60004 72208 60056 72214
rect 60004 72150 60056 72156
rect 59912 72140 59964 72146
rect 59912 72082 59964 72088
rect 59544 72004 59596 72010
rect 59544 71946 59596 71952
rect 58900 65000 58952 65006
rect 58900 64942 58952 64948
rect 59452 65000 59504 65006
rect 59452 64942 59504 64948
rect 58624 61940 58676 61946
rect 58624 61882 58676 61888
rect 58636 58478 58664 61882
rect 58716 59560 58768 59566
rect 58716 59502 58768 59508
rect 58624 58472 58676 58478
rect 58624 58414 58676 58420
rect 58728 53718 58756 59502
rect 58912 59158 58940 64942
rect 58992 61056 59044 61062
rect 58992 60998 59044 61004
rect 59004 60858 59032 60998
rect 58992 60852 59044 60858
rect 58992 60794 59044 60800
rect 58900 59152 58952 59158
rect 58900 59094 58952 59100
rect 58716 53712 58768 53718
rect 58716 53654 58768 53660
rect 58808 52080 58860 52086
rect 58808 52022 58860 52028
rect 58820 49230 58848 52022
rect 58808 49224 58860 49230
rect 58808 49166 58860 49172
rect 58912 46986 58940 59094
rect 58900 46980 58952 46986
rect 58900 46922 58952 46928
rect 58900 45076 58952 45082
rect 58900 45018 58952 45024
rect 58624 43104 58676 43110
rect 58624 43046 58676 43052
rect 58636 16794 58664 43046
rect 58912 33046 58940 45018
rect 58900 33040 58952 33046
rect 58900 32982 58952 32988
rect 59004 21418 59032 60794
rect 59268 57044 59320 57050
rect 59268 56986 59320 56992
rect 59280 55758 59308 56986
rect 59268 55752 59320 55758
rect 59268 55694 59320 55700
rect 59268 51944 59320 51950
rect 59268 51886 59320 51892
rect 59280 36582 59308 51886
rect 59268 36576 59320 36582
rect 59268 36518 59320 36524
rect 59360 24744 59412 24750
rect 59360 24686 59412 24692
rect 58992 21412 59044 21418
rect 58992 21354 59044 21360
rect 58624 16788 58676 16794
rect 58624 16730 58676 16736
rect 59268 16244 59320 16250
rect 59268 16186 59320 16192
rect 58532 4616 58584 4622
rect 58532 4558 58584 4564
rect 58624 4072 58676 4078
rect 58624 4014 58676 4020
rect 58164 3596 58216 3602
rect 58164 3538 58216 3544
rect 58072 2644 58124 2650
rect 58072 2586 58124 2592
rect 58176 800 58204 3538
rect 58348 3052 58400 3058
rect 58348 2994 58400 3000
rect 58440 3052 58492 3058
rect 58440 2994 58492 3000
rect 58360 2582 58388 2994
rect 58348 2576 58400 2582
rect 58348 2518 58400 2524
rect 58452 800 58480 2994
rect 58636 800 58664 4014
rect 59176 4004 59228 4010
rect 59176 3946 59228 3952
rect 58808 3596 58860 3602
rect 58808 3538 58860 3544
rect 58820 800 58848 3538
rect 58992 2916 59044 2922
rect 58992 2858 59044 2864
rect 59004 800 59032 2858
rect 59188 800 59216 3946
rect 59280 2582 59308 16186
rect 59372 7818 59400 24686
rect 59464 18698 59492 64942
rect 59556 43790 59584 71946
rect 60016 70446 60044 72150
rect 60096 72140 60148 72146
rect 60096 72082 60148 72088
rect 60004 70440 60056 70446
rect 60004 70382 60056 70388
rect 60108 50522 60136 72082
rect 60200 65006 60228 74506
rect 60280 65068 60332 65074
rect 60280 65010 60332 65016
rect 60188 65000 60240 65006
rect 60188 64942 60240 64948
rect 60096 50516 60148 50522
rect 60096 50458 60148 50464
rect 59544 43784 59596 43790
rect 59544 43726 59596 43732
rect 59556 43246 59584 43726
rect 59544 43240 59596 43246
rect 59544 43182 59596 43188
rect 60200 27470 60228 64942
rect 60188 27464 60240 27470
rect 60188 27406 60240 27412
rect 60292 27402 60320 65010
rect 60568 64938 60596 92550
rect 60556 64932 60608 64938
rect 60556 64874 60608 64880
rect 60648 56908 60700 56914
rect 60648 56850 60700 56856
rect 60464 55072 60516 55078
rect 60464 55014 60516 55020
rect 60476 53174 60504 55014
rect 60660 53650 60688 56850
rect 60648 53644 60700 53650
rect 60648 53586 60700 53592
rect 60464 53168 60516 53174
rect 60464 53110 60516 53116
rect 60660 53038 60688 53586
rect 60648 53032 60700 53038
rect 60648 52974 60700 52980
rect 60372 46164 60424 46170
rect 60372 46106 60424 46112
rect 60384 39030 60412 46106
rect 60752 42770 60780 96902
rect 61108 84992 61160 84998
rect 61108 84934 61160 84940
rect 60924 62892 60976 62898
rect 60924 62834 60976 62840
rect 60936 53038 60964 62834
rect 61016 53440 61068 53446
rect 61016 53382 61068 53388
rect 61028 53038 61056 53382
rect 60924 53032 60976 53038
rect 60924 52974 60976 52980
rect 61016 53032 61068 53038
rect 61016 52974 61068 52980
rect 60740 42764 60792 42770
rect 60740 42706 60792 42712
rect 60936 40050 60964 52974
rect 60924 40044 60976 40050
rect 60924 39986 60976 39992
rect 60372 39024 60424 39030
rect 60372 38966 60424 38972
rect 60280 27396 60332 27402
rect 60280 27338 60332 27344
rect 60384 23186 60412 38966
rect 60740 28620 60792 28626
rect 60740 28562 60792 28568
rect 60648 28552 60700 28558
rect 60648 28494 60700 28500
rect 60660 27946 60688 28494
rect 60648 27940 60700 27946
rect 60648 27882 60700 27888
rect 60752 23186 60780 28562
rect 59728 23180 59780 23186
rect 59728 23122 59780 23128
rect 60372 23180 60424 23186
rect 60372 23122 60424 23128
rect 60740 23180 60792 23186
rect 60740 23122 60792 23128
rect 59740 22982 59768 23122
rect 60096 23112 60148 23118
rect 60096 23054 60148 23060
rect 59728 22976 59780 22982
rect 59728 22918 59780 22924
rect 59452 18692 59504 18698
rect 59452 18634 59504 18640
rect 59464 15094 59492 18634
rect 59740 18154 59768 22918
rect 59728 18148 59780 18154
rect 59728 18090 59780 18096
rect 59452 15088 59504 15094
rect 59452 15030 59504 15036
rect 60108 12986 60136 23054
rect 61120 17882 61148 84934
rect 61200 82408 61252 82414
rect 61200 82350 61252 82356
rect 60280 17876 60332 17882
rect 60280 17818 60332 17824
rect 61108 17876 61160 17882
rect 61108 17818 61160 17824
rect 60096 12980 60148 12986
rect 60096 12922 60148 12928
rect 60188 9580 60240 9586
rect 60188 9522 60240 9528
rect 60200 8566 60228 9522
rect 60188 8560 60240 8566
rect 60188 8502 60240 8508
rect 59360 7812 59412 7818
rect 59360 7754 59412 7760
rect 59728 6860 59780 6866
rect 59728 6802 59780 6808
rect 59740 6662 59768 6802
rect 60200 6730 60228 8502
rect 60188 6724 60240 6730
rect 60188 6666 60240 6672
rect 59728 6656 59780 6662
rect 59728 6598 59780 6604
rect 59636 6180 59688 6186
rect 59636 6122 59688 6128
rect 59360 3120 59412 3126
rect 59360 3062 59412 3068
rect 59268 2576 59320 2582
rect 59268 2518 59320 2524
rect 59372 2514 59400 3062
rect 59544 2984 59596 2990
rect 59464 2944 59544 2972
rect 59360 2508 59412 2514
rect 59360 2450 59412 2456
rect 59464 800 59492 2944
rect 59544 2926 59596 2932
rect 59648 2922 59676 6122
rect 59740 6118 59768 6598
rect 59728 6112 59780 6118
rect 59728 6054 59780 6060
rect 59820 4004 59872 4010
rect 59820 3946 59872 3952
rect 59636 2916 59688 2922
rect 59636 2858 59688 2864
rect 59636 2440 59688 2446
rect 59636 2382 59688 2388
rect 59648 800 59676 2382
rect 59832 800 59860 3946
rect 60096 2984 60148 2990
rect 60016 2944 60096 2972
rect 60016 800 60044 2944
rect 60096 2926 60148 2932
rect 60188 2848 60240 2854
rect 60188 2790 60240 2796
rect 60200 800 60228 2790
rect 60292 2650 60320 17818
rect 61016 4004 61068 4010
rect 61016 3946 61068 3952
rect 60464 3936 60516 3942
rect 60464 3878 60516 3884
rect 60280 2644 60332 2650
rect 60280 2586 60332 2592
rect 60476 800 60504 3878
rect 60648 3596 60700 3602
rect 60648 3538 60700 3544
rect 60660 800 60688 3538
rect 60832 2304 60884 2310
rect 60832 2246 60884 2252
rect 60844 800 60872 2246
rect 61028 800 61056 3946
rect 61212 2582 61240 82350
rect 61396 77722 61424 97106
rect 62132 96626 62160 99200
rect 62960 97170 62988 99200
rect 63880 97238 63908 99200
rect 63868 97232 63920 97238
rect 63868 97174 63920 97180
rect 62948 97164 63000 97170
rect 62948 97106 63000 97112
rect 63960 97164 64012 97170
rect 63960 97106 64012 97112
rect 63132 96960 63184 96966
rect 63132 96902 63184 96908
rect 62120 96620 62172 96626
rect 62120 96562 62172 96568
rect 62212 96484 62264 96490
rect 62212 96426 62264 96432
rect 61660 95396 61712 95402
rect 61660 95338 61712 95344
rect 61672 93854 61700 95338
rect 61672 93826 62068 93854
rect 61568 91588 61620 91594
rect 61568 91530 61620 91536
rect 61476 91112 61528 91118
rect 61476 91054 61528 91060
rect 61384 77716 61436 77722
rect 61384 77658 61436 77664
rect 61384 68876 61436 68882
rect 61384 68818 61436 68824
rect 61292 55140 61344 55146
rect 61292 55082 61344 55088
rect 61304 28626 61332 55082
rect 61396 53174 61424 68818
rect 61384 53168 61436 53174
rect 61384 53110 61436 53116
rect 61384 51264 61436 51270
rect 61384 51206 61436 51212
rect 61292 28620 61344 28626
rect 61292 28562 61344 28568
rect 61396 7886 61424 51206
rect 61488 13258 61516 91054
rect 61580 69902 61608 91530
rect 62040 83978 62068 93826
rect 62028 83972 62080 83978
rect 62028 83914 62080 83920
rect 61936 74316 61988 74322
rect 61936 74258 61988 74264
rect 61568 69896 61620 69902
rect 61568 69838 61620 69844
rect 61948 68814 61976 74258
rect 61936 68808 61988 68814
rect 61936 68750 61988 68756
rect 61948 64122 61976 68750
rect 61936 64116 61988 64122
rect 61936 64058 61988 64064
rect 61948 61606 61976 64058
rect 61936 61600 61988 61606
rect 61936 61542 61988 61548
rect 62040 60314 62068 83914
rect 62120 79620 62172 79626
rect 62120 79562 62172 79568
rect 62132 79150 62160 79562
rect 62120 79144 62172 79150
rect 62120 79086 62172 79092
rect 62028 60308 62080 60314
rect 62028 60250 62080 60256
rect 62040 55350 62068 60250
rect 62028 55344 62080 55350
rect 62028 55286 62080 55292
rect 62028 52964 62080 52970
rect 62028 52906 62080 52912
rect 62040 51814 62068 52906
rect 62028 51808 62080 51814
rect 62028 51750 62080 51756
rect 62224 42566 62252 96426
rect 63040 94240 63092 94246
rect 63040 94182 63092 94188
rect 63052 90030 63080 94182
rect 63040 90024 63092 90030
rect 63040 89966 63092 89972
rect 62304 84584 62356 84590
rect 62304 84526 62356 84532
rect 62212 42560 62264 42566
rect 62212 42502 62264 42508
rect 61568 39976 61620 39982
rect 61568 39918 61620 39924
rect 61580 26790 61608 39918
rect 61568 26784 61620 26790
rect 61568 26726 61620 26732
rect 62028 26784 62080 26790
rect 62028 26726 62080 26732
rect 61568 23180 61620 23186
rect 61568 23122 61620 23128
rect 61580 13326 61608 23122
rect 61844 22228 61896 22234
rect 61844 22170 61896 22176
rect 61752 19916 61804 19922
rect 61752 19858 61804 19864
rect 61660 14340 61712 14346
rect 61660 14282 61712 14288
rect 61568 13320 61620 13326
rect 61568 13262 61620 13268
rect 61476 13252 61528 13258
rect 61476 13194 61528 13200
rect 61384 7880 61436 7886
rect 61384 7822 61436 7828
rect 61292 3596 61344 3602
rect 61292 3538 61344 3544
rect 61200 2576 61252 2582
rect 61200 2518 61252 2524
rect 61304 800 61332 3538
rect 61568 3052 61620 3058
rect 61568 2994 61620 3000
rect 61476 2916 61528 2922
rect 61476 2858 61528 2864
rect 61488 800 61516 2858
rect 61580 2582 61608 2994
rect 61672 2990 61700 14282
rect 61764 10266 61792 19858
rect 61856 15094 61884 22170
rect 62040 20040 62068 26726
rect 61948 20012 62068 20040
rect 61948 18766 61976 20012
rect 62212 19984 62264 19990
rect 62212 19926 62264 19932
rect 62120 19236 62172 19242
rect 62120 19178 62172 19184
rect 61936 18760 61988 18766
rect 61936 18702 61988 18708
rect 62132 18426 62160 19178
rect 62120 18420 62172 18426
rect 62120 18362 62172 18368
rect 61844 15088 61896 15094
rect 61844 15030 61896 15036
rect 62224 10266 62252 19926
rect 61752 10260 61804 10266
rect 61752 10202 61804 10208
rect 62212 10260 62264 10266
rect 62212 10202 62264 10208
rect 62316 7698 62344 84526
rect 62856 79144 62908 79150
rect 62856 79086 62908 79092
rect 62764 77716 62816 77722
rect 62764 77658 62816 77664
rect 62396 68808 62448 68814
rect 62396 68750 62448 68756
rect 62408 47530 62436 68750
rect 62672 63980 62724 63986
rect 62672 63922 62724 63928
rect 62684 63889 62712 63922
rect 62670 63880 62726 63889
rect 62670 63815 62726 63824
rect 62396 47524 62448 47530
rect 62396 47466 62448 47472
rect 62776 19242 62804 77658
rect 62868 53786 62896 79086
rect 62856 53780 62908 53786
rect 62856 53722 62908 53728
rect 62868 53582 62896 53722
rect 63040 53644 63092 53650
rect 63040 53586 63092 53592
rect 62856 53576 62908 53582
rect 62856 53518 62908 53524
rect 62856 44328 62908 44334
rect 62856 44270 62908 44276
rect 62868 20262 62896 44270
rect 63052 36242 63080 53586
rect 63144 45354 63172 96902
rect 63224 94376 63276 94382
rect 63224 94318 63276 94324
rect 63236 72010 63264 94318
rect 63408 94308 63460 94314
rect 63408 94250 63460 94256
rect 63224 72004 63276 72010
rect 63224 71946 63276 71952
rect 63420 47666 63448 94250
rect 63592 71120 63644 71126
rect 63592 71062 63644 71068
rect 63604 70394 63632 71062
rect 63512 70366 63632 70394
rect 63408 47660 63460 47666
rect 63408 47602 63460 47608
rect 63132 45348 63184 45354
rect 63132 45290 63184 45296
rect 63132 43648 63184 43654
rect 63132 43590 63184 43596
rect 63040 36236 63092 36242
rect 63040 36178 63092 36184
rect 62948 34060 63000 34066
rect 62948 34002 63000 34008
rect 62856 20256 62908 20262
rect 62856 20198 62908 20204
rect 62764 19236 62816 19242
rect 62764 19178 62816 19184
rect 62960 18902 62988 34002
rect 63052 21894 63080 36178
rect 63040 21888 63092 21894
rect 63040 21830 63092 21836
rect 62948 18896 63000 18902
rect 62948 18838 63000 18844
rect 62672 18760 62724 18766
rect 62724 18720 62804 18748
rect 62672 18702 62724 18708
rect 62396 17536 62448 17542
rect 62396 17478 62448 17484
rect 62224 7670 62344 7698
rect 61936 6248 61988 6254
rect 61936 6190 61988 6196
rect 61752 4004 61804 4010
rect 61752 3946 61804 3952
rect 61660 2984 61712 2990
rect 61660 2926 61712 2932
rect 61568 2576 61620 2582
rect 61568 2518 61620 2524
rect 61764 2122 61792 3946
rect 61844 3528 61896 3534
rect 61844 3470 61896 3476
rect 61672 2094 61792 2122
rect 61672 800 61700 2094
rect 61856 800 61884 3470
rect 61948 2582 61976 6190
rect 62224 3126 62252 7670
rect 62304 3936 62356 3942
rect 62304 3878 62356 3884
rect 62212 3120 62264 3126
rect 62212 3062 62264 3068
rect 62120 2848 62172 2854
rect 62120 2790 62172 2796
rect 62028 2644 62080 2650
rect 62028 2586 62080 2592
rect 61936 2576 61988 2582
rect 61936 2518 61988 2524
rect 62040 800 62068 2586
rect 62132 2514 62160 2790
rect 62120 2508 62172 2514
rect 62120 2450 62172 2456
rect 62316 800 62344 3878
rect 62408 3670 62436 17478
rect 62488 14068 62540 14074
rect 62488 14010 62540 14016
rect 62396 3664 62448 3670
rect 62396 3606 62448 3612
rect 62500 3194 62528 14010
rect 62776 9897 62804 18720
rect 62948 10056 63000 10062
rect 62946 10024 62948 10033
rect 63000 10024 63002 10033
rect 62946 9959 63002 9968
rect 62762 9888 62818 9897
rect 62762 9823 62818 9832
rect 62776 7886 62804 9823
rect 62764 7880 62816 7886
rect 62764 7822 62816 7828
rect 62776 6866 62804 7822
rect 62764 6860 62816 6866
rect 62764 6802 62816 6808
rect 62856 4684 62908 4690
rect 62856 4626 62908 4632
rect 62488 3188 62540 3194
rect 62488 3130 62540 3136
rect 62500 2990 62528 3130
rect 62488 2984 62540 2990
rect 62488 2926 62540 2932
rect 62672 2916 62724 2922
rect 62672 2858 62724 2864
rect 62488 2848 62540 2854
rect 62488 2790 62540 2796
rect 62500 800 62528 2790
rect 62684 800 62712 2858
rect 62868 800 62896 4626
rect 63040 3596 63092 3602
rect 63040 3538 63092 3544
rect 63052 800 63080 3538
rect 63144 2582 63172 43590
rect 63408 39432 63460 39438
rect 63408 39374 63460 39380
rect 63316 36848 63368 36854
rect 63316 36790 63368 36796
rect 63328 36174 63356 36790
rect 63420 36174 63448 39374
rect 63316 36168 63368 36174
rect 63316 36110 63368 36116
rect 63408 36168 63460 36174
rect 63408 36110 63460 36116
rect 63408 35148 63460 35154
rect 63408 35090 63460 35096
rect 63420 34066 63448 35090
rect 63408 34060 63460 34066
rect 63408 34002 63460 34008
rect 63512 28694 63540 70366
rect 63684 68672 63736 68678
rect 63684 68614 63736 68620
rect 63592 67176 63644 67182
rect 63592 67118 63644 67124
rect 63604 66842 63632 67118
rect 63592 66836 63644 66842
rect 63592 66778 63644 66784
rect 63696 60734 63724 68614
rect 63604 60706 63724 60734
rect 63604 48278 63632 60706
rect 63972 59430 64000 97106
rect 64708 96626 64736 99200
rect 65536 97238 65564 99200
rect 66456 97238 66484 99200
rect 65524 97232 65576 97238
rect 65524 97174 65576 97180
rect 66444 97232 66496 97238
rect 66444 97174 66496 97180
rect 66536 97164 66588 97170
rect 66536 97106 66588 97112
rect 65984 97028 66036 97034
rect 65984 96970 66036 96976
rect 65660 96860 65956 96880
rect 65716 96858 65740 96860
rect 65796 96858 65820 96860
rect 65876 96858 65900 96860
rect 65738 96806 65740 96858
rect 65802 96806 65814 96858
rect 65876 96806 65878 96858
rect 65716 96804 65740 96806
rect 65796 96804 65820 96806
rect 65876 96804 65900 96806
rect 65660 96784 65956 96804
rect 64696 96620 64748 96626
rect 64696 96562 64748 96568
rect 64788 96484 64840 96490
rect 64788 96426 64840 96432
rect 64144 86760 64196 86766
rect 64144 86702 64196 86708
rect 63684 59424 63736 59430
rect 63684 59366 63736 59372
rect 63960 59424 64012 59430
rect 63960 59366 64012 59372
rect 63696 52970 63724 59366
rect 64052 57520 64104 57526
rect 64052 57462 64104 57468
rect 64064 56982 64092 57462
rect 64052 56976 64104 56982
rect 64052 56918 64104 56924
rect 64052 55820 64104 55826
rect 64052 55762 64104 55768
rect 63684 52964 63736 52970
rect 63684 52906 63736 52912
rect 63776 50448 63828 50454
rect 63776 50390 63828 50396
rect 63788 49910 63816 50390
rect 63776 49904 63828 49910
rect 63776 49846 63828 49852
rect 63592 48272 63644 48278
rect 63592 48214 63644 48220
rect 64064 39846 64092 55762
rect 64052 39840 64104 39846
rect 64052 39782 64104 39788
rect 63592 36236 63644 36242
rect 63592 36178 63644 36184
rect 63500 28688 63552 28694
rect 63500 28630 63552 28636
rect 63408 18896 63460 18902
rect 63408 18838 63460 18844
rect 63420 15026 63448 18838
rect 63408 15020 63460 15026
rect 63408 14962 63460 14968
rect 63604 12102 63632 36178
rect 63684 36032 63736 36038
rect 63684 35974 63736 35980
rect 63696 12442 63724 35974
rect 64156 34134 64184 86702
rect 64328 83496 64380 83502
rect 64328 83438 64380 83444
rect 64236 70508 64288 70514
rect 64236 70450 64288 70456
rect 64144 34128 64196 34134
rect 64144 34070 64196 34076
rect 63960 31680 64012 31686
rect 63960 31622 64012 31628
rect 63972 31142 64000 31622
rect 64144 31408 64196 31414
rect 64144 31350 64196 31356
rect 64156 31210 64184 31350
rect 64144 31204 64196 31210
rect 64144 31146 64196 31152
rect 63960 31136 64012 31142
rect 63960 31078 64012 31084
rect 64052 31136 64104 31142
rect 64052 31078 64104 31084
rect 63960 28960 64012 28966
rect 63960 28902 64012 28908
rect 63972 28694 64000 28902
rect 63960 28688 64012 28694
rect 63960 28630 64012 28636
rect 63776 13184 63828 13190
rect 63776 13126 63828 13132
rect 63684 12436 63736 12442
rect 63684 12378 63736 12384
rect 63592 12096 63644 12102
rect 63592 12038 63644 12044
rect 63684 10192 63736 10198
rect 63420 10140 63684 10146
rect 63420 10134 63736 10140
rect 63420 10118 63724 10134
rect 63420 10062 63448 10118
rect 63408 10056 63460 10062
rect 63408 9998 63460 10004
rect 63592 9988 63644 9994
rect 63592 9930 63644 9936
rect 63604 9897 63632 9930
rect 63590 9888 63646 9897
rect 63590 9823 63646 9832
rect 63408 9512 63460 9518
rect 63408 9454 63460 9460
rect 63132 2576 63184 2582
rect 63132 2518 63184 2524
rect 63420 2514 63448 9454
rect 63788 8362 63816 13126
rect 63868 10056 63920 10062
rect 63866 10024 63868 10033
rect 63920 10024 63922 10033
rect 63866 9959 63922 9968
rect 63776 8356 63828 8362
rect 63776 8298 63828 8304
rect 63684 3596 63736 3602
rect 63684 3538 63736 3544
rect 63500 3528 63552 3534
rect 63500 3470 63552 3476
rect 63408 2508 63460 2514
rect 63408 2450 63460 2456
rect 63316 2372 63368 2378
rect 63316 2314 63368 2320
rect 63328 800 63356 2314
rect 63512 800 63540 3470
rect 63696 800 63724 3538
rect 64064 2582 64092 31078
rect 64248 20602 64276 70450
rect 64340 43926 64368 83438
rect 64512 57316 64564 57322
rect 64512 57258 64564 57264
rect 64524 56982 64552 57258
rect 64512 56976 64564 56982
rect 64512 56918 64564 56924
rect 64604 56908 64656 56914
rect 64604 56850 64656 56856
rect 64616 53174 64644 56850
rect 64604 53168 64656 53174
rect 64604 53110 64656 53116
rect 64420 52352 64472 52358
rect 64420 52294 64472 52300
rect 64328 43920 64380 43926
rect 64328 43862 64380 43868
rect 64328 31340 64380 31346
rect 64328 31282 64380 31288
rect 64340 30802 64368 31282
rect 64328 30796 64380 30802
rect 64328 30738 64380 30744
rect 64432 21962 64460 52294
rect 64512 48272 64564 48278
rect 64512 48214 64564 48220
rect 64420 21956 64472 21962
rect 64420 21898 64472 21904
rect 64524 21554 64552 48214
rect 64616 31754 64644 53110
rect 64696 50448 64748 50454
rect 64696 50390 64748 50396
rect 64708 47122 64736 50390
rect 64696 47116 64748 47122
rect 64696 47058 64748 47064
rect 64800 44878 64828 96426
rect 65660 95772 65956 95792
rect 65716 95770 65740 95772
rect 65796 95770 65820 95772
rect 65876 95770 65900 95772
rect 65738 95718 65740 95770
rect 65802 95718 65814 95770
rect 65876 95718 65878 95770
rect 65716 95716 65740 95718
rect 65796 95716 65820 95718
rect 65876 95716 65900 95718
rect 65660 95696 65956 95716
rect 65660 94684 65956 94704
rect 65716 94682 65740 94684
rect 65796 94682 65820 94684
rect 65876 94682 65900 94684
rect 65738 94630 65740 94682
rect 65802 94630 65814 94682
rect 65876 94630 65878 94682
rect 65716 94628 65740 94630
rect 65796 94628 65820 94630
rect 65876 94628 65900 94630
rect 65660 94608 65956 94628
rect 65660 93596 65956 93616
rect 65716 93594 65740 93596
rect 65796 93594 65820 93596
rect 65876 93594 65900 93596
rect 65738 93542 65740 93594
rect 65802 93542 65814 93594
rect 65876 93542 65878 93594
rect 65716 93540 65740 93542
rect 65796 93540 65820 93542
rect 65876 93540 65900 93542
rect 65660 93520 65956 93540
rect 65660 92508 65956 92528
rect 65716 92506 65740 92508
rect 65796 92506 65820 92508
rect 65876 92506 65900 92508
rect 65738 92454 65740 92506
rect 65802 92454 65814 92506
rect 65876 92454 65878 92506
rect 65716 92452 65740 92454
rect 65796 92452 65820 92454
rect 65876 92452 65900 92454
rect 65660 92432 65956 92452
rect 65248 91860 65300 91866
rect 65248 91802 65300 91808
rect 64880 59696 64932 59702
rect 64880 59638 64932 59644
rect 64892 59566 64920 59638
rect 64880 59560 64932 59566
rect 64880 59502 64932 59508
rect 64788 44872 64840 44878
rect 64708 44832 64788 44860
rect 64708 36242 64736 44832
rect 64788 44814 64840 44820
rect 64696 36236 64748 36242
rect 64696 36178 64748 36184
rect 64616 31726 64736 31754
rect 64604 31476 64656 31482
rect 64604 31418 64656 31424
rect 64616 31142 64644 31418
rect 64604 31136 64656 31142
rect 64604 31078 64656 31084
rect 64708 27402 64736 31726
rect 64696 27396 64748 27402
rect 64696 27338 64748 27344
rect 64512 21548 64564 21554
rect 64512 21490 64564 21496
rect 64236 20596 64288 20602
rect 64236 20538 64288 20544
rect 64696 19984 64748 19990
rect 64696 19926 64748 19932
rect 64420 8016 64472 8022
rect 64420 7958 64472 7964
rect 64432 7546 64460 7958
rect 64420 7540 64472 7546
rect 64420 7482 64472 7488
rect 64144 4072 64196 4078
rect 64144 4014 64196 4020
rect 64052 2576 64104 2582
rect 64052 2518 64104 2524
rect 63868 2440 63920 2446
rect 63868 2382 63920 2388
rect 63880 800 63908 2382
rect 64156 2122 64184 4014
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 64064 2094 64184 2122
rect 64064 800 64092 2094
rect 64340 800 64368 3538
rect 64708 2990 64736 19926
rect 64892 18902 64920 59502
rect 65064 50312 65116 50318
rect 65064 50254 65116 50260
rect 65076 48686 65104 50254
rect 65064 48680 65116 48686
rect 65064 48622 65116 48628
rect 65076 47122 65104 48622
rect 65064 47116 65116 47122
rect 65064 47058 65116 47064
rect 65260 46986 65288 91802
rect 65660 91420 65956 91440
rect 65716 91418 65740 91420
rect 65796 91418 65820 91420
rect 65876 91418 65900 91420
rect 65738 91366 65740 91418
rect 65802 91366 65814 91418
rect 65876 91366 65878 91418
rect 65716 91364 65740 91366
rect 65796 91364 65820 91366
rect 65876 91364 65900 91366
rect 65660 91344 65956 91364
rect 65660 90332 65956 90352
rect 65716 90330 65740 90332
rect 65796 90330 65820 90332
rect 65876 90330 65900 90332
rect 65738 90278 65740 90330
rect 65802 90278 65814 90330
rect 65876 90278 65878 90330
rect 65716 90276 65740 90278
rect 65796 90276 65820 90278
rect 65876 90276 65900 90278
rect 65660 90256 65956 90276
rect 65660 89244 65956 89264
rect 65716 89242 65740 89244
rect 65796 89242 65820 89244
rect 65876 89242 65900 89244
rect 65738 89190 65740 89242
rect 65802 89190 65814 89242
rect 65876 89190 65878 89242
rect 65716 89188 65740 89190
rect 65796 89188 65820 89190
rect 65876 89188 65900 89190
rect 65660 89168 65956 89188
rect 65660 88156 65956 88176
rect 65716 88154 65740 88156
rect 65796 88154 65820 88156
rect 65876 88154 65900 88156
rect 65738 88102 65740 88154
rect 65802 88102 65814 88154
rect 65876 88102 65878 88154
rect 65716 88100 65740 88102
rect 65796 88100 65820 88102
rect 65876 88100 65900 88102
rect 65660 88080 65956 88100
rect 65660 87068 65956 87088
rect 65716 87066 65740 87068
rect 65796 87066 65820 87068
rect 65876 87066 65900 87068
rect 65738 87014 65740 87066
rect 65802 87014 65814 87066
rect 65876 87014 65878 87066
rect 65716 87012 65740 87014
rect 65796 87012 65820 87014
rect 65876 87012 65900 87014
rect 65660 86992 65956 87012
rect 65660 85980 65956 86000
rect 65716 85978 65740 85980
rect 65796 85978 65820 85980
rect 65876 85978 65900 85980
rect 65738 85926 65740 85978
rect 65802 85926 65814 85978
rect 65876 85926 65878 85978
rect 65716 85924 65740 85926
rect 65796 85924 65820 85926
rect 65876 85924 65900 85926
rect 65660 85904 65956 85924
rect 65660 84892 65956 84912
rect 65716 84890 65740 84892
rect 65796 84890 65820 84892
rect 65876 84890 65900 84892
rect 65738 84838 65740 84890
rect 65802 84838 65814 84890
rect 65876 84838 65878 84890
rect 65716 84836 65740 84838
rect 65796 84836 65820 84838
rect 65876 84836 65900 84838
rect 65660 84816 65956 84836
rect 65996 84182 66024 96970
rect 66076 94852 66128 94858
rect 66076 94794 66128 94800
rect 65984 84176 66036 84182
rect 65984 84118 66036 84124
rect 65524 83904 65576 83910
rect 65524 83846 65576 83852
rect 65432 71528 65484 71534
rect 65432 71470 65484 71476
rect 65444 71398 65472 71470
rect 65432 71392 65484 71398
rect 65432 71334 65484 71340
rect 65444 59702 65472 71334
rect 65432 59696 65484 59702
rect 65432 59638 65484 59644
rect 65340 59424 65392 59430
rect 65340 59366 65392 59372
rect 65248 46980 65300 46986
rect 65248 46922 65300 46928
rect 65156 25356 65208 25362
rect 65156 25298 65208 25304
rect 64972 24132 65024 24138
rect 64972 24074 65024 24080
rect 64984 19922 65012 24074
rect 65168 20058 65196 25298
rect 65156 20052 65208 20058
rect 65156 19994 65208 20000
rect 64972 19916 65024 19922
rect 64972 19858 65024 19864
rect 64880 18896 64932 18902
rect 64880 18838 64932 18844
rect 65352 18834 65380 59366
rect 65432 34944 65484 34950
rect 65432 34886 65484 34892
rect 65444 34678 65472 34886
rect 65432 34672 65484 34678
rect 65432 34614 65484 34620
rect 65432 34468 65484 34474
rect 65432 34410 65484 34416
rect 65444 34202 65472 34410
rect 65432 34196 65484 34202
rect 65432 34138 65484 34144
rect 65432 33584 65484 33590
rect 65432 33526 65484 33532
rect 65444 18970 65472 33526
rect 65536 22166 65564 83846
rect 65660 83804 65956 83824
rect 65716 83802 65740 83804
rect 65796 83802 65820 83804
rect 65876 83802 65900 83804
rect 65738 83750 65740 83802
rect 65802 83750 65814 83802
rect 65876 83750 65878 83802
rect 65716 83748 65740 83750
rect 65796 83748 65820 83750
rect 65876 83748 65900 83750
rect 65660 83728 65956 83748
rect 65660 82716 65956 82736
rect 65716 82714 65740 82716
rect 65796 82714 65820 82716
rect 65876 82714 65900 82716
rect 65738 82662 65740 82714
rect 65802 82662 65814 82714
rect 65876 82662 65878 82714
rect 65716 82660 65740 82662
rect 65796 82660 65820 82662
rect 65876 82660 65900 82662
rect 65660 82640 65956 82660
rect 65984 82408 66036 82414
rect 65984 82350 66036 82356
rect 65660 81628 65956 81648
rect 65716 81626 65740 81628
rect 65796 81626 65820 81628
rect 65876 81626 65900 81628
rect 65738 81574 65740 81626
rect 65802 81574 65814 81626
rect 65876 81574 65878 81626
rect 65716 81572 65740 81574
rect 65796 81572 65820 81574
rect 65876 81572 65900 81574
rect 65660 81552 65956 81572
rect 65660 80540 65956 80560
rect 65716 80538 65740 80540
rect 65796 80538 65820 80540
rect 65876 80538 65900 80540
rect 65738 80486 65740 80538
rect 65802 80486 65814 80538
rect 65876 80486 65878 80538
rect 65716 80484 65740 80486
rect 65796 80484 65820 80486
rect 65876 80484 65900 80486
rect 65660 80464 65956 80484
rect 65660 79452 65956 79472
rect 65716 79450 65740 79452
rect 65796 79450 65820 79452
rect 65876 79450 65900 79452
rect 65738 79398 65740 79450
rect 65802 79398 65814 79450
rect 65876 79398 65878 79450
rect 65716 79396 65740 79398
rect 65796 79396 65820 79398
rect 65876 79396 65900 79398
rect 65660 79376 65956 79396
rect 65660 78364 65956 78384
rect 65716 78362 65740 78364
rect 65796 78362 65820 78364
rect 65876 78362 65900 78364
rect 65738 78310 65740 78362
rect 65802 78310 65814 78362
rect 65876 78310 65878 78362
rect 65716 78308 65740 78310
rect 65796 78308 65820 78310
rect 65876 78308 65900 78310
rect 65660 78288 65956 78308
rect 65660 77276 65956 77296
rect 65716 77274 65740 77276
rect 65796 77274 65820 77276
rect 65876 77274 65900 77276
rect 65738 77222 65740 77274
rect 65802 77222 65814 77274
rect 65876 77222 65878 77274
rect 65716 77220 65740 77222
rect 65796 77220 65820 77222
rect 65876 77220 65900 77222
rect 65660 77200 65956 77220
rect 65660 76188 65956 76208
rect 65716 76186 65740 76188
rect 65796 76186 65820 76188
rect 65876 76186 65900 76188
rect 65738 76134 65740 76186
rect 65802 76134 65814 76186
rect 65876 76134 65878 76186
rect 65716 76132 65740 76134
rect 65796 76132 65820 76134
rect 65876 76132 65900 76134
rect 65660 76112 65956 76132
rect 65660 75100 65956 75120
rect 65716 75098 65740 75100
rect 65796 75098 65820 75100
rect 65876 75098 65900 75100
rect 65738 75046 65740 75098
rect 65802 75046 65814 75098
rect 65876 75046 65878 75098
rect 65716 75044 65740 75046
rect 65796 75044 65820 75046
rect 65876 75044 65900 75046
rect 65660 75024 65956 75044
rect 65660 74012 65956 74032
rect 65716 74010 65740 74012
rect 65796 74010 65820 74012
rect 65876 74010 65900 74012
rect 65738 73958 65740 74010
rect 65802 73958 65814 74010
rect 65876 73958 65878 74010
rect 65716 73956 65740 73958
rect 65796 73956 65820 73958
rect 65876 73956 65900 73958
rect 65660 73936 65956 73956
rect 65660 72924 65956 72944
rect 65716 72922 65740 72924
rect 65796 72922 65820 72924
rect 65876 72922 65900 72924
rect 65738 72870 65740 72922
rect 65802 72870 65814 72922
rect 65876 72870 65878 72922
rect 65716 72868 65740 72870
rect 65796 72868 65820 72870
rect 65876 72868 65900 72870
rect 65660 72848 65956 72868
rect 65660 71836 65956 71856
rect 65716 71834 65740 71836
rect 65796 71834 65820 71836
rect 65876 71834 65900 71836
rect 65738 71782 65740 71834
rect 65802 71782 65814 71834
rect 65876 71782 65878 71834
rect 65716 71780 65740 71782
rect 65796 71780 65820 71782
rect 65876 71780 65900 71782
rect 65660 71760 65956 71780
rect 65660 70748 65956 70768
rect 65716 70746 65740 70748
rect 65796 70746 65820 70748
rect 65876 70746 65900 70748
rect 65738 70694 65740 70746
rect 65802 70694 65814 70746
rect 65876 70694 65878 70746
rect 65716 70692 65740 70694
rect 65796 70692 65820 70694
rect 65876 70692 65900 70694
rect 65660 70672 65956 70692
rect 65660 69660 65956 69680
rect 65716 69658 65740 69660
rect 65796 69658 65820 69660
rect 65876 69658 65900 69660
rect 65738 69606 65740 69658
rect 65802 69606 65814 69658
rect 65876 69606 65878 69658
rect 65716 69604 65740 69606
rect 65796 69604 65820 69606
rect 65876 69604 65900 69606
rect 65660 69584 65956 69604
rect 65660 68572 65956 68592
rect 65716 68570 65740 68572
rect 65796 68570 65820 68572
rect 65876 68570 65900 68572
rect 65738 68518 65740 68570
rect 65802 68518 65814 68570
rect 65876 68518 65878 68570
rect 65716 68516 65740 68518
rect 65796 68516 65820 68518
rect 65876 68516 65900 68518
rect 65660 68496 65956 68516
rect 65660 67484 65956 67504
rect 65716 67482 65740 67484
rect 65796 67482 65820 67484
rect 65876 67482 65900 67484
rect 65738 67430 65740 67482
rect 65802 67430 65814 67482
rect 65876 67430 65878 67482
rect 65716 67428 65740 67430
rect 65796 67428 65820 67430
rect 65876 67428 65900 67430
rect 65660 67408 65956 67428
rect 65660 66396 65956 66416
rect 65716 66394 65740 66396
rect 65796 66394 65820 66396
rect 65876 66394 65900 66396
rect 65738 66342 65740 66394
rect 65802 66342 65814 66394
rect 65876 66342 65878 66394
rect 65716 66340 65740 66342
rect 65796 66340 65820 66342
rect 65876 66340 65900 66342
rect 65660 66320 65956 66340
rect 65660 65308 65956 65328
rect 65716 65306 65740 65308
rect 65796 65306 65820 65308
rect 65876 65306 65900 65308
rect 65738 65254 65740 65306
rect 65802 65254 65814 65306
rect 65876 65254 65878 65306
rect 65716 65252 65740 65254
rect 65796 65252 65820 65254
rect 65876 65252 65900 65254
rect 65660 65232 65956 65252
rect 65660 64220 65956 64240
rect 65716 64218 65740 64220
rect 65796 64218 65820 64220
rect 65876 64218 65900 64220
rect 65738 64166 65740 64218
rect 65802 64166 65814 64218
rect 65876 64166 65878 64218
rect 65716 64164 65740 64166
rect 65796 64164 65820 64166
rect 65876 64164 65900 64166
rect 65660 64144 65956 64164
rect 65660 63132 65956 63152
rect 65716 63130 65740 63132
rect 65796 63130 65820 63132
rect 65876 63130 65900 63132
rect 65738 63078 65740 63130
rect 65802 63078 65814 63130
rect 65876 63078 65878 63130
rect 65716 63076 65740 63078
rect 65796 63076 65820 63078
rect 65876 63076 65900 63078
rect 65660 63056 65956 63076
rect 65628 62478 65840 62506
rect 65628 62354 65656 62478
rect 65708 62416 65760 62422
rect 65708 62358 65760 62364
rect 65616 62348 65668 62354
rect 65616 62290 65668 62296
rect 65720 62286 65748 62358
rect 65812 62354 65840 62478
rect 65800 62348 65852 62354
rect 65800 62290 65852 62296
rect 65708 62280 65760 62286
rect 65708 62222 65760 62228
rect 65660 62044 65956 62064
rect 65716 62042 65740 62044
rect 65796 62042 65820 62044
rect 65876 62042 65900 62044
rect 65738 61990 65740 62042
rect 65802 61990 65814 62042
rect 65876 61990 65878 62042
rect 65716 61988 65740 61990
rect 65796 61988 65820 61990
rect 65876 61988 65900 61990
rect 65660 61968 65956 61988
rect 65660 60956 65956 60976
rect 65716 60954 65740 60956
rect 65796 60954 65820 60956
rect 65876 60954 65900 60956
rect 65738 60902 65740 60954
rect 65802 60902 65814 60954
rect 65876 60902 65878 60954
rect 65716 60900 65740 60902
rect 65796 60900 65820 60902
rect 65876 60900 65900 60902
rect 65660 60880 65956 60900
rect 65660 59868 65956 59888
rect 65716 59866 65740 59868
rect 65796 59866 65820 59868
rect 65876 59866 65900 59868
rect 65738 59814 65740 59866
rect 65802 59814 65814 59866
rect 65876 59814 65878 59866
rect 65716 59812 65740 59814
rect 65796 59812 65820 59814
rect 65876 59812 65900 59814
rect 65660 59792 65956 59812
rect 65660 58780 65956 58800
rect 65716 58778 65740 58780
rect 65796 58778 65820 58780
rect 65876 58778 65900 58780
rect 65738 58726 65740 58778
rect 65802 58726 65814 58778
rect 65876 58726 65878 58778
rect 65716 58724 65740 58726
rect 65796 58724 65820 58726
rect 65876 58724 65900 58726
rect 65660 58704 65956 58724
rect 65660 57692 65956 57712
rect 65716 57690 65740 57692
rect 65796 57690 65820 57692
rect 65876 57690 65900 57692
rect 65738 57638 65740 57690
rect 65802 57638 65814 57690
rect 65876 57638 65878 57690
rect 65716 57636 65740 57638
rect 65796 57636 65820 57638
rect 65876 57636 65900 57638
rect 65660 57616 65956 57636
rect 65660 56604 65956 56624
rect 65716 56602 65740 56604
rect 65796 56602 65820 56604
rect 65876 56602 65900 56604
rect 65738 56550 65740 56602
rect 65802 56550 65814 56602
rect 65876 56550 65878 56602
rect 65716 56548 65740 56550
rect 65796 56548 65820 56550
rect 65876 56548 65900 56550
rect 65660 56528 65956 56548
rect 65660 55516 65956 55536
rect 65716 55514 65740 55516
rect 65796 55514 65820 55516
rect 65876 55514 65900 55516
rect 65738 55462 65740 55514
rect 65802 55462 65814 55514
rect 65876 55462 65878 55514
rect 65716 55460 65740 55462
rect 65796 55460 65820 55462
rect 65876 55460 65900 55462
rect 65660 55440 65956 55460
rect 65660 54428 65956 54448
rect 65716 54426 65740 54428
rect 65796 54426 65820 54428
rect 65876 54426 65900 54428
rect 65738 54374 65740 54426
rect 65802 54374 65814 54426
rect 65876 54374 65878 54426
rect 65716 54372 65740 54374
rect 65796 54372 65820 54374
rect 65876 54372 65900 54374
rect 65660 54352 65956 54372
rect 65660 53340 65956 53360
rect 65716 53338 65740 53340
rect 65796 53338 65820 53340
rect 65876 53338 65900 53340
rect 65738 53286 65740 53338
rect 65802 53286 65814 53338
rect 65876 53286 65878 53338
rect 65716 53284 65740 53286
rect 65796 53284 65820 53286
rect 65876 53284 65900 53286
rect 65660 53264 65956 53284
rect 65660 52252 65956 52272
rect 65716 52250 65740 52252
rect 65796 52250 65820 52252
rect 65876 52250 65900 52252
rect 65738 52198 65740 52250
rect 65802 52198 65814 52250
rect 65876 52198 65878 52250
rect 65716 52196 65740 52198
rect 65796 52196 65820 52198
rect 65876 52196 65900 52198
rect 65660 52176 65956 52196
rect 65660 51164 65956 51184
rect 65716 51162 65740 51164
rect 65796 51162 65820 51164
rect 65876 51162 65900 51164
rect 65738 51110 65740 51162
rect 65802 51110 65814 51162
rect 65876 51110 65878 51162
rect 65716 51108 65740 51110
rect 65796 51108 65820 51110
rect 65876 51108 65900 51110
rect 65660 51088 65956 51108
rect 65660 50076 65956 50096
rect 65716 50074 65740 50076
rect 65796 50074 65820 50076
rect 65876 50074 65900 50076
rect 65738 50022 65740 50074
rect 65802 50022 65814 50074
rect 65876 50022 65878 50074
rect 65716 50020 65740 50022
rect 65796 50020 65820 50022
rect 65876 50020 65900 50022
rect 65660 50000 65956 50020
rect 65660 48988 65956 49008
rect 65716 48986 65740 48988
rect 65796 48986 65820 48988
rect 65876 48986 65900 48988
rect 65738 48934 65740 48986
rect 65802 48934 65814 48986
rect 65876 48934 65878 48986
rect 65716 48932 65740 48934
rect 65796 48932 65820 48934
rect 65876 48932 65900 48934
rect 65660 48912 65956 48932
rect 65660 47900 65956 47920
rect 65716 47898 65740 47900
rect 65796 47898 65820 47900
rect 65876 47898 65900 47900
rect 65738 47846 65740 47898
rect 65802 47846 65814 47898
rect 65876 47846 65878 47898
rect 65716 47844 65740 47846
rect 65796 47844 65820 47846
rect 65876 47844 65900 47846
rect 65660 47824 65956 47844
rect 65660 46812 65956 46832
rect 65716 46810 65740 46812
rect 65796 46810 65820 46812
rect 65876 46810 65900 46812
rect 65738 46758 65740 46810
rect 65802 46758 65814 46810
rect 65876 46758 65878 46810
rect 65716 46756 65740 46758
rect 65796 46756 65820 46758
rect 65876 46756 65900 46758
rect 65660 46736 65956 46756
rect 65660 45724 65956 45744
rect 65716 45722 65740 45724
rect 65796 45722 65820 45724
rect 65876 45722 65900 45724
rect 65738 45670 65740 45722
rect 65802 45670 65814 45722
rect 65876 45670 65878 45722
rect 65716 45668 65740 45670
rect 65796 45668 65820 45670
rect 65876 45668 65900 45670
rect 65660 45648 65956 45668
rect 65660 44636 65956 44656
rect 65716 44634 65740 44636
rect 65796 44634 65820 44636
rect 65876 44634 65900 44636
rect 65738 44582 65740 44634
rect 65802 44582 65814 44634
rect 65876 44582 65878 44634
rect 65716 44580 65740 44582
rect 65796 44580 65820 44582
rect 65876 44580 65900 44582
rect 65660 44560 65956 44580
rect 65660 43548 65956 43568
rect 65716 43546 65740 43548
rect 65796 43546 65820 43548
rect 65876 43546 65900 43548
rect 65738 43494 65740 43546
rect 65802 43494 65814 43546
rect 65876 43494 65878 43546
rect 65716 43492 65740 43494
rect 65796 43492 65820 43494
rect 65876 43492 65900 43494
rect 65660 43472 65956 43492
rect 65660 42460 65956 42480
rect 65716 42458 65740 42460
rect 65796 42458 65820 42460
rect 65876 42458 65900 42460
rect 65738 42406 65740 42458
rect 65802 42406 65814 42458
rect 65876 42406 65878 42458
rect 65716 42404 65740 42406
rect 65796 42404 65820 42406
rect 65876 42404 65900 42406
rect 65660 42384 65956 42404
rect 65660 41372 65956 41392
rect 65716 41370 65740 41372
rect 65796 41370 65820 41372
rect 65876 41370 65900 41372
rect 65738 41318 65740 41370
rect 65802 41318 65814 41370
rect 65876 41318 65878 41370
rect 65716 41316 65740 41318
rect 65796 41316 65820 41318
rect 65876 41316 65900 41318
rect 65660 41296 65956 41316
rect 65660 40284 65956 40304
rect 65716 40282 65740 40284
rect 65796 40282 65820 40284
rect 65876 40282 65900 40284
rect 65738 40230 65740 40282
rect 65802 40230 65814 40282
rect 65876 40230 65878 40282
rect 65716 40228 65740 40230
rect 65796 40228 65820 40230
rect 65876 40228 65900 40230
rect 65660 40208 65956 40228
rect 65660 39196 65956 39216
rect 65716 39194 65740 39196
rect 65796 39194 65820 39196
rect 65876 39194 65900 39196
rect 65738 39142 65740 39194
rect 65802 39142 65814 39194
rect 65876 39142 65878 39194
rect 65716 39140 65740 39142
rect 65796 39140 65820 39142
rect 65876 39140 65900 39142
rect 65660 39120 65956 39140
rect 65660 38108 65956 38128
rect 65716 38106 65740 38108
rect 65796 38106 65820 38108
rect 65876 38106 65900 38108
rect 65738 38054 65740 38106
rect 65802 38054 65814 38106
rect 65876 38054 65878 38106
rect 65716 38052 65740 38054
rect 65796 38052 65820 38054
rect 65876 38052 65900 38054
rect 65660 38032 65956 38052
rect 65660 37020 65956 37040
rect 65716 37018 65740 37020
rect 65796 37018 65820 37020
rect 65876 37018 65900 37020
rect 65738 36966 65740 37018
rect 65802 36966 65814 37018
rect 65876 36966 65878 37018
rect 65716 36964 65740 36966
rect 65796 36964 65820 36966
rect 65876 36964 65900 36966
rect 65660 36944 65956 36964
rect 65660 35932 65956 35952
rect 65716 35930 65740 35932
rect 65796 35930 65820 35932
rect 65876 35930 65900 35932
rect 65738 35878 65740 35930
rect 65802 35878 65814 35930
rect 65876 35878 65878 35930
rect 65716 35876 65740 35878
rect 65796 35876 65820 35878
rect 65876 35876 65900 35878
rect 65660 35856 65956 35876
rect 65660 34844 65956 34864
rect 65716 34842 65740 34844
rect 65796 34842 65820 34844
rect 65876 34842 65900 34844
rect 65738 34790 65740 34842
rect 65802 34790 65814 34842
rect 65876 34790 65878 34842
rect 65716 34788 65740 34790
rect 65796 34788 65820 34790
rect 65876 34788 65900 34790
rect 65660 34768 65956 34788
rect 65616 34400 65668 34406
rect 65616 34342 65668 34348
rect 65628 34066 65656 34342
rect 65616 34060 65668 34066
rect 65616 34002 65668 34008
rect 65660 33756 65956 33776
rect 65716 33754 65740 33756
rect 65796 33754 65820 33756
rect 65876 33754 65900 33756
rect 65738 33702 65740 33754
rect 65802 33702 65814 33754
rect 65876 33702 65878 33754
rect 65716 33700 65740 33702
rect 65796 33700 65820 33702
rect 65876 33700 65900 33702
rect 65660 33680 65956 33700
rect 65660 32668 65956 32688
rect 65716 32666 65740 32668
rect 65796 32666 65820 32668
rect 65876 32666 65900 32668
rect 65738 32614 65740 32666
rect 65802 32614 65814 32666
rect 65876 32614 65878 32666
rect 65716 32612 65740 32614
rect 65796 32612 65820 32614
rect 65876 32612 65900 32614
rect 65660 32592 65956 32612
rect 65660 31580 65956 31600
rect 65716 31578 65740 31580
rect 65796 31578 65820 31580
rect 65876 31578 65900 31580
rect 65738 31526 65740 31578
rect 65802 31526 65814 31578
rect 65876 31526 65878 31578
rect 65716 31524 65740 31526
rect 65796 31524 65820 31526
rect 65876 31524 65900 31526
rect 65660 31504 65956 31524
rect 65660 30492 65956 30512
rect 65716 30490 65740 30492
rect 65796 30490 65820 30492
rect 65876 30490 65900 30492
rect 65738 30438 65740 30490
rect 65802 30438 65814 30490
rect 65876 30438 65878 30490
rect 65716 30436 65740 30438
rect 65796 30436 65820 30438
rect 65876 30436 65900 30438
rect 65660 30416 65956 30436
rect 65660 29404 65956 29424
rect 65716 29402 65740 29404
rect 65796 29402 65820 29404
rect 65876 29402 65900 29404
rect 65738 29350 65740 29402
rect 65802 29350 65814 29402
rect 65876 29350 65878 29402
rect 65716 29348 65740 29350
rect 65796 29348 65820 29350
rect 65876 29348 65900 29350
rect 65660 29328 65956 29348
rect 65660 28316 65956 28336
rect 65716 28314 65740 28316
rect 65796 28314 65820 28316
rect 65876 28314 65900 28316
rect 65738 28262 65740 28314
rect 65802 28262 65814 28314
rect 65876 28262 65878 28314
rect 65716 28260 65740 28262
rect 65796 28260 65820 28262
rect 65876 28260 65900 28262
rect 65660 28240 65956 28260
rect 65660 27228 65956 27248
rect 65716 27226 65740 27228
rect 65796 27226 65820 27228
rect 65876 27226 65900 27228
rect 65738 27174 65740 27226
rect 65802 27174 65814 27226
rect 65876 27174 65878 27226
rect 65716 27172 65740 27174
rect 65796 27172 65820 27174
rect 65876 27172 65900 27174
rect 65660 27152 65956 27172
rect 65660 26140 65956 26160
rect 65716 26138 65740 26140
rect 65796 26138 65820 26140
rect 65876 26138 65900 26140
rect 65738 26086 65740 26138
rect 65802 26086 65814 26138
rect 65876 26086 65878 26138
rect 65716 26084 65740 26086
rect 65796 26084 65820 26086
rect 65876 26084 65900 26086
rect 65660 26064 65956 26084
rect 65660 25052 65956 25072
rect 65716 25050 65740 25052
rect 65796 25050 65820 25052
rect 65876 25050 65900 25052
rect 65738 24998 65740 25050
rect 65802 24998 65814 25050
rect 65876 24998 65878 25050
rect 65716 24996 65740 24998
rect 65796 24996 65820 24998
rect 65876 24996 65900 24998
rect 65660 24976 65956 24996
rect 65660 23964 65956 23984
rect 65716 23962 65740 23964
rect 65796 23962 65820 23964
rect 65876 23962 65900 23964
rect 65738 23910 65740 23962
rect 65802 23910 65814 23962
rect 65876 23910 65878 23962
rect 65716 23908 65740 23910
rect 65796 23908 65820 23910
rect 65876 23908 65900 23910
rect 65660 23888 65956 23908
rect 65660 22876 65956 22896
rect 65716 22874 65740 22876
rect 65796 22874 65820 22876
rect 65876 22874 65900 22876
rect 65738 22822 65740 22874
rect 65802 22822 65814 22874
rect 65876 22822 65878 22874
rect 65716 22820 65740 22822
rect 65796 22820 65820 22822
rect 65876 22820 65900 22822
rect 65660 22800 65956 22820
rect 65524 22160 65576 22166
rect 65524 22102 65576 22108
rect 65660 21788 65956 21808
rect 65716 21786 65740 21788
rect 65796 21786 65820 21788
rect 65876 21786 65900 21788
rect 65738 21734 65740 21786
rect 65802 21734 65814 21786
rect 65876 21734 65878 21786
rect 65716 21732 65740 21734
rect 65796 21732 65820 21734
rect 65876 21732 65900 21734
rect 65660 21712 65956 21732
rect 65660 20700 65956 20720
rect 65716 20698 65740 20700
rect 65796 20698 65820 20700
rect 65876 20698 65900 20700
rect 65738 20646 65740 20698
rect 65802 20646 65814 20698
rect 65876 20646 65878 20698
rect 65716 20644 65740 20646
rect 65796 20644 65820 20646
rect 65876 20644 65900 20646
rect 65660 20624 65956 20644
rect 65660 19612 65956 19632
rect 65716 19610 65740 19612
rect 65796 19610 65820 19612
rect 65876 19610 65900 19612
rect 65738 19558 65740 19610
rect 65802 19558 65814 19610
rect 65876 19558 65878 19610
rect 65716 19556 65740 19558
rect 65796 19556 65820 19558
rect 65876 19556 65900 19558
rect 65660 19536 65956 19556
rect 65432 18964 65484 18970
rect 65432 18906 65484 18912
rect 65340 18828 65392 18834
rect 65340 18770 65392 18776
rect 65660 18524 65956 18544
rect 65716 18522 65740 18524
rect 65796 18522 65820 18524
rect 65876 18522 65900 18524
rect 65738 18470 65740 18522
rect 65802 18470 65814 18522
rect 65876 18470 65878 18522
rect 65716 18468 65740 18470
rect 65796 18468 65820 18470
rect 65876 18468 65900 18470
rect 65660 18448 65956 18468
rect 65660 17436 65956 17456
rect 65716 17434 65740 17436
rect 65796 17434 65820 17436
rect 65876 17434 65900 17436
rect 65738 17382 65740 17434
rect 65802 17382 65814 17434
rect 65876 17382 65878 17434
rect 65716 17380 65740 17382
rect 65796 17380 65820 17382
rect 65876 17380 65900 17382
rect 65660 17360 65956 17380
rect 65996 16574 66024 82350
rect 66088 78606 66116 94794
rect 66168 94444 66220 94450
rect 66168 94386 66220 94392
rect 66076 78600 66128 78606
rect 66076 78542 66128 78548
rect 66088 59430 66116 78542
rect 66180 78266 66208 94386
rect 66168 78260 66220 78266
rect 66168 78202 66220 78208
rect 66180 71602 66208 78202
rect 66168 71596 66220 71602
rect 66168 71538 66220 71544
rect 66352 64116 66404 64122
rect 66352 64058 66404 64064
rect 66364 64025 66392 64058
rect 66350 64016 66406 64025
rect 66350 63951 66406 63960
rect 66548 60734 66576 97106
rect 67284 96626 67312 99200
rect 68204 97170 68232 99200
rect 68560 97504 68612 97510
rect 68560 97446 68612 97452
rect 68572 97238 68600 97446
rect 69032 97238 69060 99200
rect 69952 97238 69980 99200
rect 68560 97232 68612 97238
rect 68560 97174 68612 97180
rect 69020 97232 69072 97238
rect 69020 97174 69072 97180
rect 69940 97232 69992 97238
rect 69940 97174 69992 97180
rect 68192 97164 68244 97170
rect 68192 97106 68244 97112
rect 69296 97164 69348 97170
rect 69296 97106 69348 97112
rect 67272 96620 67324 96626
rect 67272 96562 67324 96568
rect 66904 95464 66956 95470
rect 66904 95406 66956 95412
rect 66916 83910 66944 95406
rect 69308 93838 69336 97106
rect 69664 97096 69716 97102
rect 69664 97038 69716 97044
rect 69296 93832 69348 93838
rect 69296 93774 69348 93780
rect 69308 93158 69336 93774
rect 69296 93152 69348 93158
rect 69296 93094 69348 93100
rect 68928 92336 68980 92342
rect 68928 92278 68980 92284
rect 68940 91730 68968 92278
rect 68468 91724 68520 91730
rect 68468 91666 68520 91672
rect 68928 91724 68980 91730
rect 68928 91666 68980 91672
rect 68284 88392 68336 88398
rect 68284 88334 68336 88340
rect 66904 83904 66956 83910
rect 66904 83846 66956 83852
rect 67548 83904 67600 83910
rect 67548 83846 67600 83852
rect 66628 71528 66680 71534
rect 66628 71470 66680 71476
rect 66272 60706 66576 60734
rect 66076 59424 66128 59430
rect 66076 59366 66128 59372
rect 66272 55162 66300 60706
rect 66180 55134 66300 55162
rect 66640 55146 66668 71470
rect 67088 64320 67140 64326
rect 67088 64262 67140 64268
rect 66996 64048 67048 64054
rect 66994 64016 66996 64025
rect 67048 64016 67050 64025
rect 66994 63951 67050 63960
rect 66352 55140 66404 55146
rect 66076 53032 66128 53038
rect 66076 52974 66128 52980
rect 66088 25702 66116 52974
rect 66180 46442 66208 55134
rect 66352 55082 66404 55088
rect 66628 55140 66680 55146
rect 66628 55082 66680 55088
rect 66364 51950 66392 55082
rect 66904 53168 66956 53174
rect 66904 53110 66956 53116
rect 66352 51944 66404 51950
rect 66352 51886 66404 51892
rect 66168 46436 66220 46442
rect 66168 46378 66220 46384
rect 66180 40390 66208 46378
rect 66720 43920 66772 43926
rect 66720 43862 66772 43868
rect 66168 40384 66220 40390
rect 66168 40326 66220 40332
rect 66180 33590 66208 40326
rect 66260 35012 66312 35018
rect 66260 34954 66312 34960
rect 66272 34542 66300 34954
rect 66444 34944 66496 34950
rect 66444 34886 66496 34892
rect 66456 34746 66484 34886
rect 66444 34740 66496 34746
rect 66444 34682 66496 34688
rect 66456 34542 66484 34682
rect 66628 34672 66680 34678
rect 66628 34614 66680 34620
rect 66640 34542 66668 34614
rect 66260 34536 66312 34542
rect 66260 34478 66312 34484
rect 66444 34536 66496 34542
rect 66444 34478 66496 34484
rect 66628 34536 66680 34542
rect 66628 34478 66680 34484
rect 66168 33584 66220 33590
rect 66168 33526 66220 33532
rect 66272 33318 66300 34478
rect 66260 33312 66312 33318
rect 66260 33254 66312 33260
rect 66076 25696 66128 25702
rect 66076 25638 66128 25644
rect 66260 25696 66312 25702
rect 66260 25638 66312 25644
rect 66272 25498 66300 25638
rect 66260 25492 66312 25498
rect 66260 25434 66312 25440
rect 66260 20596 66312 20602
rect 66260 20538 66312 20544
rect 65996 16546 66116 16574
rect 65660 16348 65956 16368
rect 65716 16346 65740 16348
rect 65796 16346 65820 16348
rect 65876 16346 65900 16348
rect 65738 16294 65740 16346
rect 65802 16294 65814 16346
rect 65876 16294 65878 16346
rect 65716 16292 65740 16294
rect 65796 16292 65820 16294
rect 65876 16292 65900 16294
rect 65660 16272 65956 16292
rect 65660 15260 65956 15280
rect 65716 15258 65740 15260
rect 65796 15258 65820 15260
rect 65876 15258 65900 15260
rect 65738 15206 65740 15258
rect 65802 15206 65814 15258
rect 65876 15206 65878 15258
rect 65716 15204 65740 15206
rect 65796 15204 65820 15206
rect 65876 15204 65900 15206
rect 65660 15184 65956 15204
rect 65660 14172 65956 14192
rect 65716 14170 65740 14172
rect 65796 14170 65820 14172
rect 65876 14170 65900 14172
rect 65738 14118 65740 14170
rect 65802 14118 65814 14170
rect 65876 14118 65878 14170
rect 65716 14116 65740 14118
rect 65796 14116 65820 14118
rect 65876 14116 65900 14118
rect 65660 14096 65956 14116
rect 65660 13084 65956 13104
rect 65716 13082 65740 13084
rect 65796 13082 65820 13084
rect 65876 13082 65900 13084
rect 65738 13030 65740 13082
rect 65802 13030 65814 13082
rect 65876 13030 65878 13082
rect 65716 13028 65740 13030
rect 65796 13028 65820 13030
rect 65876 13028 65900 13030
rect 65660 13008 65956 13028
rect 65660 11996 65956 12016
rect 65716 11994 65740 11996
rect 65796 11994 65820 11996
rect 65876 11994 65900 11996
rect 65738 11942 65740 11994
rect 65802 11942 65814 11994
rect 65876 11942 65878 11994
rect 65716 11940 65740 11942
rect 65796 11940 65820 11942
rect 65876 11940 65900 11942
rect 65660 11920 65956 11940
rect 65660 10908 65956 10928
rect 65716 10906 65740 10908
rect 65796 10906 65820 10908
rect 65876 10906 65900 10908
rect 65738 10854 65740 10906
rect 65802 10854 65814 10906
rect 65876 10854 65878 10906
rect 65716 10852 65740 10854
rect 65796 10852 65820 10854
rect 65876 10852 65900 10854
rect 65660 10832 65956 10852
rect 65660 9820 65956 9840
rect 65716 9818 65740 9820
rect 65796 9818 65820 9820
rect 65876 9818 65900 9820
rect 65738 9766 65740 9818
rect 65802 9766 65814 9818
rect 65876 9766 65878 9818
rect 65716 9764 65740 9766
rect 65796 9764 65820 9766
rect 65876 9764 65900 9766
rect 65660 9744 65956 9764
rect 65660 8732 65956 8752
rect 65716 8730 65740 8732
rect 65796 8730 65820 8732
rect 65876 8730 65900 8732
rect 65738 8678 65740 8730
rect 65802 8678 65814 8730
rect 65876 8678 65878 8730
rect 65716 8676 65740 8678
rect 65796 8676 65820 8678
rect 65876 8676 65900 8678
rect 65660 8656 65956 8676
rect 65660 7644 65956 7664
rect 65716 7642 65740 7644
rect 65796 7642 65820 7644
rect 65876 7642 65900 7644
rect 65738 7590 65740 7642
rect 65802 7590 65814 7642
rect 65876 7590 65878 7642
rect 65716 7588 65740 7590
rect 65796 7588 65820 7590
rect 65876 7588 65900 7590
rect 65660 7568 65956 7588
rect 65660 6556 65956 6576
rect 65716 6554 65740 6556
rect 65796 6554 65820 6556
rect 65876 6554 65900 6556
rect 65738 6502 65740 6554
rect 65802 6502 65814 6554
rect 65876 6502 65878 6554
rect 65716 6500 65740 6502
rect 65796 6500 65820 6502
rect 65876 6500 65900 6502
rect 65660 6480 65956 6500
rect 65660 5468 65956 5488
rect 65716 5466 65740 5468
rect 65796 5466 65820 5468
rect 65876 5466 65900 5468
rect 65738 5414 65740 5466
rect 65802 5414 65814 5466
rect 65876 5414 65878 5466
rect 65716 5412 65740 5414
rect 65796 5412 65820 5414
rect 65876 5412 65900 5414
rect 65660 5392 65956 5412
rect 65156 4480 65208 4486
rect 65156 4422 65208 4428
rect 65168 4282 65196 4422
rect 65660 4380 65956 4400
rect 65716 4378 65740 4380
rect 65796 4378 65820 4380
rect 65876 4378 65900 4380
rect 65738 4326 65740 4378
rect 65802 4326 65814 4378
rect 65876 4326 65878 4378
rect 65716 4324 65740 4326
rect 65796 4324 65820 4326
rect 65876 4324 65900 4326
rect 65660 4304 65956 4324
rect 65156 4276 65208 4282
rect 65156 4218 65208 4224
rect 64788 4072 64840 4078
rect 64788 4014 64840 4020
rect 65984 4072 66036 4078
rect 65984 4014 66036 4020
rect 64696 2984 64748 2990
rect 64696 2926 64748 2932
rect 64512 2916 64564 2922
rect 64512 2858 64564 2864
rect 64524 800 64552 2858
rect 64800 2122 64828 4014
rect 65340 3596 65392 3602
rect 65340 3538 65392 3544
rect 64880 2984 64932 2990
rect 64880 2926 64932 2932
rect 64708 2094 64828 2122
rect 64708 800 64736 2094
rect 64892 800 64920 2926
rect 65064 2304 65116 2310
rect 65064 2246 65116 2252
rect 65076 800 65104 2246
rect 65352 800 65380 3538
rect 65660 3292 65956 3312
rect 65716 3290 65740 3292
rect 65796 3290 65820 3292
rect 65876 3290 65900 3292
rect 65738 3238 65740 3290
rect 65802 3238 65814 3290
rect 65876 3238 65878 3290
rect 65716 3236 65740 3238
rect 65796 3236 65820 3238
rect 65876 3236 65900 3238
rect 65660 3216 65956 3236
rect 65524 2984 65576 2990
rect 65524 2926 65576 2932
rect 65536 800 65564 2926
rect 65660 2204 65956 2224
rect 65716 2202 65740 2204
rect 65796 2202 65820 2204
rect 65876 2202 65900 2204
rect 65738 2150 65740 2202
rect 65802 2150 65814 2202
rect 65876 2150 65878 2202
rect 65716 2148 65740 2150
rect 65796 2148 65820 2150
rect 65876 2148 65900 2150
rect 65660 2128 65956 2148
rect 65996 1986 66024 4014
rect 66088 2582 66116 16546
rect 66168 3052 66220 3058
rect 66168 2994 66220 3000
rect 66076 2576 66128 2582
rect 66076 2518 66128 2524
rect 65904 1958 66024 1986
rect 65708 1420 65760 1426
rect 65708 1362 65760 1368
rect 65720 800 65748 1362
rect 65904 800 65932 1958
rect 66180 800 66208 2994
rect 66272 2650 66300 20538
rect 66628 13252 66680 13258
rect 66628 13194 66680 13200
rect 66352 13184 66404 13190
rect 66352 13126 66404 13132
rect 66364 12782 66392 13126
rect 66640 12782 66668 13194
rect 66352 12776 66404 12782
rect 66352 12718 66404 12724
rect 66628 12776 66680 12782
rect 66628 12718 66680 12724
rect 66536 4072 66588 4078
rect 66536 4014 66588 4020
rect 66260 2644 66312 2650
rect 66260 2586 66312 2592
rect 66352 2508 66404 2514
rect 66352 2450 66404 2456
rect 66364 800 66392 2450
rect 66444 2372 66496 2378
rect 66444 2314 66496 2320
rect 66456 1426 66484 2314
rect 66444 1420 66496 1426
rect 66444 1362 66496 1368
rect 66548 800 66576 4014
rect 66732 3194 66760 43862
rect 66916 41274 66944 53110
rect 66996 53032 67048 53038
rect 66996 52974 67048 52980
rect 66904 41268 66956 41274
rect 66904 41210 66956 41216
rect 66916 40934 66944 41210
rect 66904 40928 66956 40934
rect 66904 40870 66956 40876
rect 67008 39302 67036 52974
rect 66996 39296 67048 39302
rect 66996 39238 67048 39244
rect 66812 36372 66864 36378
rect 66812 36314 66864 36320
rect 66824 34490 66852 36314
rect 66904 35012 66956 35018
rect 66904 34954 66956 34960
rect 66916 34678 66944 34954
rect 66904 34672 66956 34678
rect 66904 34614 66956 34620
rect 66904 34536 66956 34542
rect 66824 34484 66904 34490
rect 66824 34478 66956 34484
rect 66824 34462 66944 34478
rect 66904 33312 66956 33318
rect 66904 33254 66956 33260
rect 66916 23730 66944 33254
rect 67008 29238 67036 39238
rect 67100 32434 67128 64262
rect 67454 64016 67510 64025
rect 67272 63980 67324 63986
rect 67454 63951 67510 63960
rect 67272 63922 67324 63928
rect 67284 63889 67312 63922
rect 67270 63880 67326 63889
rect 67270 63815 67326 63824
rect 67468 63782 67496 63951
rect 67456 63776 67508 63782
rect 67456 63718 67508 63724
rect 67560 60654 67588 83846
rect 68100 71052 68152 71058
rect 68100 70994 68152 71000
rect 68112 60858 68140 70994
rect 68100 60852 68152 60858
rect 68100 60794 68152 60800
rect 67548 60648 67600 60654
rect 67824 60648 67876 60654
rect 67548 60590 67600 60596
rect 67652 60608 67824 60636
rect 67180 59968 67232 59974
rect 67180 59910 67232 59916
rect 67088 32428 67140 32434
rect 67088 32370 67140 32376
rect 67088 31136 67140 31142
rect 67088 31078 67140 31084
rect 67100 30598 67128 31078
rect 67088 30592 67140 30598
rect 67088 30534 67140 30540
rect 66996 29232 67048 29238
rect 66996 29174 67048 29180
rect 67100 28914 67128 30534
rect 67008 28886 67128 28914
rect 66904 23724 66956 23730
rect 66904 23666 66956 23672
rect 67008 22778 67036 28886
rect 67088 25696 67140 25702
rect 67088 25638 67140 25644
rect 66996 22772 67048 22778
rect 66996 22714 67048 22720
rect 66996 17876 67048 17882
rect 66996 17818 67048 17824
rect 67008 17202 67036 17818
rect 66996 17196 67048 17202
rect 66996 17138 67048 17144
rect 66812 14816 66864 14822
rect 66812 14758 66864 14764
rect 66824 12782 66852 14758
rect 67008 12782 67036 17138
rect 67100 12782 67128 25638
rect 67192 14346 67220 59910
rect 67364 52896 67416 52902
rect 67364 52838 67416 52844
rect 67376 52698 67404 52838
rect 67364 52692 67416 52698
rect 67364 52634 67416 52640
rect 67376 52358 67404 52634
rect 67364 52352 67416 52358
rect 67364 52294 67416 52300
rect 67560 48754 67588 60590
rect 67652 60246 67680 60608
rect 67824 60590 67876 60596
rect 68008 60648 68060 60654
rect 68008 60590 68060 60596
rect 68020 60314 68048 60590
rect 68008 60308 68060 60314
rect 68008 60250 68060 60256
rect 67640 60240 67692 60246
rect 67640 60182 67692 60188
rect 67652 49910 67680 60182
rect 67640 49904 67692 49910
rect 67640 49846 67692 49852
rect 67548 48748 67600 48754
rect 67548 48690 67600 48696
rect 67732 48680 67784 48686
rect 67732 48622 67784 48628
rect 67744 40526 67772 48622
rect 67732 40520 67784 40526
rect 67732 40462 67784 40468
rect 67744 40118 67772 40462
rect 67732 40112 67784 40118
rect 67732 40054 67784 40060
rect 67824 34536 67876 34542
rect 67824 34478 67876 34484
rect 67836 33930 67864 34478
rect 67824 33924 67876 33930
rect 67824 33866 67876 33872
rect 67824 31476 67876 31482
rect 67824 31418 67876 31424
rect 67836 30802 67864 31418
rect 67916 30864 67968 30870
rect 67916 30806 67968 30812
rect 67824 30796 67876 30802
rect 67824 30738 67876 30744
rect 67836 30394 67864 30738
rect 67928 30394 67956 30806
rect 67824 30388 67876 30394
rect 67824 30330 67876 30336
rect 67916 30388 67968 30394
rect 67916 30330 67968 30336
rect 67640 19304 67692 19310
rect 67640 19246 67692 19252
rect 67652 18358 67680 19246
rect 67640 18352 67692 18358
rect 67640 18294 67692 18300
rect 67730 18320 67786 18329
rect 67548 16448 67600 16454
rect 67548 16390 67600 16396
rect 67180 14340 67232 14346
rect 67180 14282 67232 14288
rect 67364 13388 67416 13394
rect 67364 13330 67416 13336
rect 66812 12776 66864 12782
rect 66812 12718 66864 12724
rect 66996 12776 67048 12782
rect 66996 12718 67048 12724
rect 67088 12776 67140 12782
rect 67088 12718 67140 12724
rect 67088 8356 67140 8362
rect 67088 8298 67140 8304
rect 66812 3596 66864 3602
rect 66812 3538 66864 3544
rect 66720 3188 66772 3194
rect 66720 3130 66772 3136
rect 66732 2990 66760 3130
rect 66720 2984 66772 2990
rect 66720 2926 66772 2932
rect 66824 1850 66852 3538
rect 66904 2916 66956 2922
rect 66904 2858 66956 2864
rect 66732 1822 66852 1850
rect 66732 800 66760 1822
rect 66916 800 66944 2858
rect 67100 2582 67128 8298
rect 67376 5302 67404 13330
rect 67560 12782 67588 16390
rect 67548 12776 67600 12782
rect 67548 12718 67600 12724
rect 67652 12442 67680 18294
rect 67730 18255 67732 18264
rect 67784 18255 67786 18264
rect 67732 18226 67784 18232
rect 67640 12436 67692 12442
rect 67640 12378 67692 12384
rect 67744 12374 67772 18226
rect 67732 12368 67784 12374
rect 67732 12310 67784 12316
rect 68296 9518 68324 88334
rect 68376 75336 68428 75342
rect 68376 75278 68428 75284
rect 68388 19922 68416 75278
rect 68480 64122 68508 91666
rect 68560 91316 68612 91322
rect 68560 91258 68612 91264
rect 68572 75478 68600 91258
rect 69676 89714 69704 97038
rect 70780 96558 70808 99200
rect 71700 97186 71728 99200
rect 71044 97164 71096 97170
rect 71700 97158 71820 97186
rect 71044 97106 71096 97112
rect 70768 96552 70820 96558
rect 70768 96494 70820 96500
rect 70860 96416 70912 96422
rect 70860 96358 70912 96364
rect 69848 90636 69900 90642
rect 69848 90578 69900 90584
rect 69676 89686 69796 89714
rect 69768 87786 69796 89686
rect 69756 87780 69808 87786
rect 69756 87722 69808 87728
rect 68836 82476 68888 82482
rect 68836 82418 68888 82424
rect 68560 75472 68612 75478
rect 68560 75414 68612 75420
rect 68468 64116 68520 64122
rect 68468 64058 68520 64064
rect 68376 19916 68428 19922
rect 68376 19858 68428 19864
rect 68376 16788 68428 16794
rect 68376 16730 68428 16736
rect 68284 9512 68336 9518
rect 68284 9454 68336 9460
rect 67364 5296 67416 5302
rect 67364 5238 67416 5244
rect 67180 4072 67232 4078
rect 67180 4014 67232 4020
rect 67732 4072 67784 4078
rect 67732 4014 67784 4020
rect 67088 2576 67140 2582
rect 67088 2518 67140 2524
rect 67192 800 67220 4014
rect 67364 2916 67416 2922
rect 67364 2858 67416 2864
rect 67376 800 67404 2858
rect 67548 2440 67600 2446
rect 67548 2382 67600 2388
rect 67560 800 67588 2382
rect 67744 800 67772 4014
rect 67916 3596 67968 3602
rect 67916 3538 67968 3544
rect 67928 800 67956 3538
rect 68388 2582 68416 16730
rect 68480 5370 68508 64058
rect 68744 56908 68796 56914
rect 68744 56850 68796 56856
rect 68756 55758 68784 56850
rect 68744 55752 68796 55758
rect 68744 55694 68796 55700
rect 68560 40724 68612 40730
rect 68560 40666 68612 40672
rect 68572 40526 68600 40666
rect 68560 40520 68612 40526
rect 68560 40462 68612 40468
rect 68572 30784 68600 40462
rect 68652 40112 68704 40118
rect 68652 40054 68704 40060
rect 68664 31346 68692 40054
rect 68652 31340 68704 31346
rect 68652 31282 68704 31288
rect 68744 31136 68796 31142
rect 68744 31078 68796 31084
rect 68652 30796 68704 30802
rect 68572 30756 68652 30784
rect 68652 30738 68704 30744
rect 68468 5364 68520 5370
rect 68468 5306 68520 5312
rect 68468 4072 68520 4078
rect 68468 4014 68520 4020
rect 68376 2576 68428 2582
rect 68376 2518 68428 2524
rect 68480 2122 68508 4014
rect 68664 3738 68692 30738
rect 68756 30734 68784 31078
rect 68744 30728 68796 30734
rect 68744 30670 68796 30676
rect 68652 3732 68704 3738
rect 68652 3674 68704 3680
rect 68560 3596 68612 3602
rect 68560 3538 68612 3544
rect 68388 2094 68508 2122
rect 68192 1420 68244 1426
rect 68192 1362 68244 1368
rect 68204 800 68232 1362
rect 68388 800 68416 2094
rect 68572 800 68600 3538
rect 68848 2650 68876 82418
rect 69664 49428 69716 49434
rect 69664 49370 69716 49376
rect 68928 47048 68980 47054
rect 68928 46990 68980 46996
rect 68940 40526 68968 46990
rect 69572 44192 69624 44198
rect 69572 44134 69624 44140
rect 69204 43716 69256 43722
rect 69204 43658 69256 43664
rect 68928 40520 68980 40526
rect 68928 40462 68980 40468
rect 69020 39500 69072 39506
rect 69020 39442 69072 39448
rect 68928 39296 68980 39302
rect 68928 39238 68980 39244
rect 68940 39098 68968 39238
rect 68928 39092 68980 39098
rect 68928 39034 68980 39040
rect 69032 26790 69060 39442
rect 69216 39370 69244 43658
rect 69204 39364 69256 39370
rect 69204 39306 69256 39312
rect 69480 31680 69532 31686
rect 69480 31622 69532 31628
rect 69492 30870 69520 31622
rect 69480 30864 69532 30870
rect 69480 30806 69532 30812
rect 69020 26784 69072 26790
rect 69020 26726 69072 26732
rect 69480 26036 69532 26042
rect 69480 25978 69532 25984
rect 68928 4072 68980 4078
rect 68928 4014 68980 4020
rect 68836 2644 68888 2650
rect 68836 2586 68888 2592
rect 68744 1488 68796 1494
rect 68744 1430 68796 1436
rect 68756 800 68784 1430
rect 68940 800 68968 4014
rect 69204 3596 69256 3602
rect 69204 3538 69256 3544
rect 69112 2372 69164 2378
rect 69112 2314 69164 2320
rect 69124 1426 69152 2314
rect 69112 1420 69164 1426
rect 69112 1362 69164 1368
rect 69216 800 69244 3538
rect 69388 2916 69440 2922
rect 69388 2858 69440 2864
rect 69400 800 69428 2858
rect 69492 2650 69520 25978
rect 69584 21690 69612 44134
rect 69676 30802 69704 49370
rect 69664 30796 69716 30802
rect 69664 30738 69716 30744
rect 69768 30122 69796 87722
rect 69860 56370 69888 90578
rect 70308 90568 70360 90574
rect 70308 90510 70360 90516
rect 70216 73228 70268 73234
rect 70216 73170 70268 73176
rect 70124 71460 70176 71466
rect 70124 71402 70176 71408
rect 70032 70644 70084 70650
rect 70032 70586 70084 70592
rect 69848 56364 69900 56370
rect 69848 56306 69900 56312
rect 69940 54528 69992 54534
rect 69940 54470 69992 54476
rect 69848 31952 69900 31958
rect 69848 31894 69900 31900
rect 69756 30116 69808 30122
rect 69756 30058 69808 30064
rect 69768 27962 69796 30058
rect 69676 27934 69796 27962
rect 69572 21684 69624 21690
rect 69572 21626 69624 21632
rect 69676 5778 69704 27934
rect 69756 26784 69808 26790
rect 69756 26726 69808 26732
rect 69768 15910 69796 26726
rect 69860 17882 69888 31894
rect 69848 17876 69900 17882
rect 69848 17818 69900 17824
rect 69756 15904 69808 15910
rect 69756 15846 69808 15852
rect 69756 13320 69808 13326
rect 69756 13262 69808 13268
rect 69768 12986 69796 13262
rect 69756 12980 69808 12986
rect 69756 12922 69808 12928
rect 69664 5772 69716 5778
rect 69664 5714 69716 5720
rect 69952 4282 69980 54470
rect 70044 39642 70072 70586
rect 70136 49434 70164 71402
rect 70228 67114 70256 73170
rect 70216 67108 70268 67114
rect 70216 67050 70268 67056
rect 70124 49428 70176 49434
rect 70124 49370 70176 49376
rect 70032 39636 70084 39642
rect 70032 39578 70084 39584
rect 70228 31958 70256 67050
rect 70320 62286 70348 90510
rect 70768 89412 70820 89418
rect 70768 89354 70820 89360
rect 70676 71528 70728 71534
rect 70676 71470 70728 71476
rect 70308 62280 70360 62286
rect 70308 62222 70360 62228
rect 70320 36038 70348 62222
rect 70688 45082 70716 71470
rect 70676 45076 70728 45082
rect 70676 45018 70728 45024
rect 70492 44396 70544 44402
rect 70492 44338 70544 44344
rect 70308 36032 70360 36038
rect 70308 35974 70360 35980
rect 70320 34746 70348 35974
rect 70308 34740 70360 34746
rect 70308 34682 70360 34688
rect 70216 31952 70268 31958
rect 70216 31894 70268 31900
rect 70032 31408 70084 31414
rect 70032 31350 70084 31356
rect 70044 30802 70072 31350
rect 70504 30802 70532 44338
rect 70032 30796 70084 30802
rect 70032 30738 70084 30744
rect 70492 30796 70544 30802
rect 70492 30738 70544 30744
rect 70032 30592 70084 30598
rect 70032 30534 70084 30540
rect 70044 30394 70072 30534
rect 70032 30388 70084 30394
rect 70032 30330 70084 30336
rect 70400 27328 70452 27334
rect 70400 27270 70452 27276
rect 70412 26926 70440 27270
rect 70400 26920 70452 26926
rect 70400 26862 70452 26868
rect 70584 18896 70636 18902
rect 70584 18838 70636 18844
rect 70596 18222 70624 18838
rect 70584 18216 70636 18222
rect 70490 18184 70546 18193
rect 70584 18158 70636 18164
rect 70490 18119 70492 18128
rect 70544 18119 70546 18128
rect 70492 18090 70544 18096
rect 70780 9450 70808 89354
rect 70872 71534 70900 96358
rect 71056 83706 71084 97106
rect 71792 96966 71820 97158
rect 71872 97164 71924 97170
rect 71872 97106 71924 97112
rect 72332 97164 72384 97170
rect 72332 97106 72384 97112
rect 71136 96960 71188 96966
rect 71136 96902 71188 96908
rect 71780 96960 71832 96966
rect 71780 96902 71832 96908
rect 71148 96626 71176 96902
rect 71136 96620 71188 96626
rect 71136 96562 71188 96568
rect 71884 94246 71912 97106
rect 71872 94240 71924 94246
rect 71872 94182 71924 94188
rect 71136 88868 71188 88874
rect 71136 88810 71188 88816
rect 71044 83700 71096 83706
rect 71044 83642 71096 83648
rect 71056 82278 71084 83642
rect 71148 83502 71176 88810
rect 71136 83496 71188 83502
rect 71136 83438 71188 83444
rect 71044 82272 71096 82278
rect 71044 82214 71096 82220
rect 71148 71534 71176 83438
rect 71780 76560 71832 76566
rect 71780 76502 71832 76508
rect 71792 75954 71820 76502
rect 71780 75948 71832 75954
rect 71780 75890 71832 75896
rect 72240 74792 72292 74798
rect 72240 74734 72292 74740
rect 71228 71664 71280 71670
rect 71228 71606 71280 71612
rect 70860 71528 70912 71534
rect 70860 71470 70912 71476
rect 71136 71528 71188 71534
rect 71136 71470 71188 71476
rect 70952 71460 71004 71466
rect 70952 71402 71004 71408
rect 70964 33114 70992 71402
rect 71148 53174 71176 71470
rect 71136 53168 71188 53174
rect 71136 53110 71188 53116
rect 71148 52562 71176 53110
rect 71136 52556 71188 52562
rect 71136 52498 71188 52504
rect 71044 52352 71096 52358
rect 71044 52294 71096 52300
rect 70952 33108 71004 33114
rect 70952 33050 71004 33056
rect 70768 9444 70820 9450
rect 70768 9386 70820 9392
rect 71056 6254 71084 52294
rect 71240 47734 71268 71606
rect 71688 63844 71740 63850
rect 71688 63786 71740 63792
rect 71320 61736 71372 61742
rect 71320 61678 71372 61684
rect 71332 55214 71360 61678
rect 71332 55186 71636 55214
rect 71608 50250 71636 55186
rect 71700 53106 71728 63786
rect 71688 53100 71740 53106
rect 71688 53042 71740 53048
rect 71596 50244 71648 50250
rect 71596 50186 71648 50192
rect 71228 47728 71280 47734
rect 71228 47670 71280 47676
rect 71228 46368 71280 46374
rect 71228 46310 71280 46316
rect 71136 43104 71188 43110
rect 71136 43046 71188 43052
rect 71148 22098 71176 43046
rect 71136 22092 71188 22098
rect 71136 22034 71188 22040
rect 71136 18352 71188 18358
rect 71134 18320 71136 18329
rect 71188 18320 71190 18329
rect 71134 18255 71190 18264
rect 71240 17270 71268 46310
rect 71504 39976 71556 39982
rect 71504 39918 71556 39924
rect 71320 33108 71372 33114
rect 71320 33050 71372 33056
rect 71332 31822 71360 33050
rect 71320 31816 71372 31822
rect 71320 31758 71372 31764
rect 71332 25498 71360 31758
rect 71412 31136 71464 31142
rect 71412 31078 71464 31084
rect 71424 27334 71452 31078
rect 71412 27328 71464 27334
rect 71412 27270 71464 27276
rect 71320 25492 71372 25498
rect 71320 25434 71372 25440
rect 71412 24948 71464 24954
rect 71412 24890 71464 24896
rect 71320 20800 71372 20806
rect 71320 20742 71372 20748
rect 71332 18358 71360 20742
rect 71320 18352 71372 18358
rect 71320 18294 71372 18300
rect 71318 18184 71374 18193
rect 71318 18119 71320 18128
rect 71372 18119 71374 18128
rect 71320 18090 71372 18096
rect 71228 17264 71280 17270
rect 71228 17206 71280 17212
rect 71424 16046 71452 24890
rect 71412 16040 71464 16046
rect 71412 15982 71464 15988
rect 71044 6248 71096 6254
rect 71044 6190 71096 6196
rect 69940 4276 69992 4282
rect 69940 4218 69992 4224
rect 70676 4208 70728 4214
rect 70676 4150 70728 4156
rect 69940 4140 69992 4146
rect 69940 4082 69992 4088
rect 69572 4004 69624 4010
rect 69572 3946 69624 3952
rect 69480 2644 69532 2650
rect 69480 2586 69532 2592
rect 69584 800 69612 3946
rect 69756 3596 69808 3602
rect 69756 3538 69808 3544
rect 69768 800 69796 3538
rect 69952 2990 69980 4082
rect 70400 3596 70452 3602
rect 70400 3538 70452 3544
rect 70216 3528 70268 3534
rect 70216 3470 70268 3476
rect 69940 2984 69992 2990
rect 69940 2926 69992 2932
rect 69848 2508 69900 2514
rect 69848 2450 69900 2456
rect 69860 1494 69888 2450
rect 70032 2304 70084 2310
rect 70032 2246 70084 2252
rect 69848 1488 69900 1494
rect 69848 1430 69900 1436
rect 70044 800 70072 2246
rect 70228 800 70256 3470
rect 70412 800 70440 3538
rect 70584 2916 70636 2922
rect 70584 2858 70636 2864
rect 70596 800 70624 2858
rect 70688 2650 70716 4150
rect 70768 4072 70820 4078
rect 70768 4014 70820 4020
rect 71412 4072 71464 4078
rect 71412 4014 71464 4020
rect 70676 2644 70728 2650
rect 70676 2586 70728 2592
rect 70780 800 70808 4014
rect 71044 2984 71096 2990
rect 71044 2926 71096 2932
rect 71056 800 71084 2926
rect 71228 2508 71280 2514
rect 71228 2450 71280 2456
rect 71240 800 71268 2450
rect 71424 800 71452 4014
rect 71516 2650 71544 39918
rect 71608 31278 71636 50186
rect 71700 49774 71728 53042
rect 71780 52896 71832 52902
rect 71780 52838 71832 52844
rect 71688 49768 71740 49774
rect 71688 49710 71740 49716
rect 71688 48000 71740 48006
rect 71688 47942 71740 47948
rect 71700 44402 71728 47942
rect 71792 46578 71820 52838
rect 71780 46572 71832 46578
rect 71780 46514 71832 46520
rect 71688 44396 71740 44402
rect 71688 44338 71740 44344
rect 72056 39976 72108 39982
rect 72056 39918 72108 39924
rect 71596 31272 71648 31278
rect 71596 31214 71648 31220
rect 72068 23050 72096 39918
rect 72252 38350 72280 74734
rect 72344 60042 72372 97106
rect 72528 96966 72556 99200
rect 73356 97170 73384 99200
rect 74276 97238 74304 99200
rect 74264 97232 74316 97238
rect 74264 97174 74316 97180
rect 73344 97164 73396 97170
rect 73344 97106 73396 97112
rect 74448 97164 74500 97170
rect 74448 97106 74500 97112
rect 72516 96960 72568 96966
rect 72516 96902 72568 96908
rect 72424 94240 72476 94246
rect 72424 94182 72476 94188
rect 72436 74866 72464 94182
rect 74460 93294 74488 97106
rect 75104 96626 75132 99200
rect 76024 97238 76052 99200
rect 76852 97238 76880 99200
rect 76012 97232 76064 97238
rect 76012 97174 76064 97180
rect 76840 97232 76892 97238
rect 76840 97174 76892 97180
rect 75184 97164 75236 97170
rect 75184 97106 75236 97112
rect 77300 97164 77352 97170
rect 77300 97106 77352 97112
rect 75092 96620 75144 96626
rect 75092 96562 75144 96568
rect 74540 96484 74592 96490
rect 74540 96426 74592 96432
rect 74448 93288 74500 93294
rect 74448 93230 74500 93236
rect 73620 91724 73672 91730
rect 73620 91666 73672 91672
rect 74172 91724 74224 91730
rect 74172 91666 74224 91672
rect 73528 87372 73580 87378
rect 73528 87314 73580 87320
rect 72516 85196 72568 85202
rect 72516 85138 72568 85144
rect 72528 76566 72556 85138
rect 72516 76560 72568 76566
rect 72516 76502 72568 76508
rect 72424 74860 72476 74866
rect 72424 74802 72476 74808
rect 72700 74792 72752 74798
rect 72700 74734 72752 74740
rect 72884 74792 72936 74798
rect 72884 74734 72936 74740
rect 72976 74792 73028 74798
rect 72976 74734 73028 74740
rect 72712 74534 72740 74734
rect 72712 74506 72832 74534
rect 72700 67176 72752 67182
rect 72700 67118 72752 67124
rect 72712 65550 72740 67118
rect 72700 65544 72752 65550
rect 72700 65486 72752 65492
rect 72424 62416 72476 62422
rect 72424 62358 72476 62364
rect 72436 62150 72464 62358
rect 72424 62144 72476 62150
rect 72424 62086 72476 62092
rect 72712 60246 72740 65486
rect 72700 60240 72752 60246
rect 72700 60182 72752 60188
rect 72332 60036 72384 60042
rect 72332 59978 72384 59984
rect 72516 45008 72568 45014
rect 72516 44950 72568 44956
rect 72424 43988 72476 43994
rect 72424 43930 72476 43936
rect 72436 42906 72464 43930
rect 72424 42900 72476 42906
rect 72424 42842 72476 42848
rect 72240 38344 72292 38350
rect 72240 38286 72292 38292
rect 72332 34944 72384 34950
rect 72332 34886 72384 34892
rect 72344 26246 72372 34886
rect 72332 26240 72384 26246
rect 72332 26182 72384 26188
rect 72344 25226 72372 26182
rect 72332 25220 72384 25226
rect 72332 25162 72384 25168
rect 72056 23044 72108 23050
rect 72056 22986 72108 22992
rect 72240 22160 72292 22166
rect 72240 22102 72292 22108
rect 71688 20052 71740 20058
rect 71688 19994 71740 20000
rect 71700 19378 71728 19994
rect 71688 19372 71740 19378
rect 71688 19314 71740 19320
rect 71700 18222 71728 19314
rect 71688 18216 71740 18222
rect 71688 18158 71740 18164
rect 72056 4072 72108 4078
rect 72056 4014 72108 4020
rect 71596 3596 71648 3602
rect 71596 3538 71648 3544
rect 71504 2644 71556 2650
rect 71504 2586 71556 2592
rect 71608 800 71636 3538
rect 71872 2372 71924 2378
rect 71872 2314 71924 2320
rect 71884 1170 71912 2314
rect 71792 1142 71912 1170
rect 71792 800 71820 1142
rect 72068 800 72096 4014
rect 72252 3194 72280 22102
rect 72436 17270 72464 42842
rect 72528 42702 72556 44950
rect 72516 42696 72568 42702
rect 72516 42638 72568 42644
rect 72516 42356 72568 42362
rect 72516 42298 72568 42304
rect 72528 41750 72556 42298
rect 72516 41744 72568 41750
rect 72516 41686 72568 41692
rect 72424 17264 72476 17270
rect 72424 17206 72476 17212
rect 72528 17202 72556 41686
rect 72804 25906 72832 74506
rect 72896 42362 72924 74734
rect 72988 43994 73016 74734
rect 73540 67658 73568 87314
rect 73528 67652 73580 67658
rect 73528 67594 73580 67600
rect 73632 61402 73660 91666
rect 73988 91656 74040 91662
rect 73988 91598 74040 91604
rect 74000 91322 74028 91598
rect 73988 91316 74040 91322
rect 73988 91258 74040 91264
rect 73804 89548 73856 89554
rect 73804 89490 73856 89496
rect 73712 87304 73764 87310
rect 73712 87246 73764 87252
rect 73620 61396 73672 61402
rect 73620 61338 73672 61344
rect 73252 46912 73304 46918
rect 73252 46854 73304 46860
rect 73160 44940 73212 44946
rect 73160 44882 73212 44888
rect 72976 43988 73028 43994
rect 72976 43930 73028 43936
rect 73068 42696 73120 42702
rect 73172 42650 73200 44882
rect 73120 42644 73200 42650
rect 73068 42638 73200 42644
rect 73080 42622 73200 42638
rect 72884 42356 72936 42362
rect 72884 42298 72936 42304
rect 73160 39840 73212 39846
rect 73160 39782 73212 39788
rect 73172 39030 73200 39782
rect 73160 39024 73212 39030
rect 73160 38966 73212 38972
rect 73068 38344 73120 38350
rect 73068 38286 73120 38292
rect 73080 32230 73108 38286
rect 73264 37398 73292 46854
rect 73528 42764 73580 42770
rect 73528 42706 73580 42712
rect 73540 42566 73568 42706
rect 73528 42560 73580 42566
rect 73528 42502 73580 42508
rect 73620 40044 73672 40050
rect 73620 39986 73672 39992
rect 73344 39908 73396 39914
rect 73344 39850 73396 39856
rect 73356 38486 73384 39850
rect 73344 38480 73396 38486
rect 73396 38428 73568 38434
rect 73344 38422 73568 38428
rect 73356 38406 73568 38422
rect 73540 38350 73568 38406
rect 73528 38344 73580 38350
rect 73528 38286 73580 38292
rect 73632 38214 73660 39986
rect 73620 38208 73672 38214
rect 73620 38150 73672 38156
rect 73528 37664 73580 37670
rect 73528 37606 73580 37612
rect 73252 37392 73304 37398
rect 73252 37334 73304 37340
rect 73436 35828 73488 35834
rect 73436 35770 73488 35776
rect 73448 34542 73476 35770
rect 73436 34536 73488 34542
rect 73436 34478 73488 34484
rect 73252 34196 73304 34202
rect 73252 34138 73304 34144
rect 73068 32224 73120 32230
rect 73068 32166 73120 32172
rect 72792 25900 72844 25906
rect 72792 25842 72844 25848
rect 72700 25220 72752 25226
rect 72700 25162 72752 25168
rect 72608 17332 72660 17338
rect 72608 17274 72660 17280
rect 72516 17196 72568 17202
rect 72516 17138 72568 17144
rect 72620 6914 72648 17274
rect 72528 6886 72648 6914
rect 72240 3188 72292 3194
rect 72240 3130 72292 3136
rect 72252 2990 72280 3130
rect 72240 2984 72292 2990
rect 72240 2926 72292 2932
rect 72424 2916 72476 2922
rect 72424 2858 72476 2864
rect 72240 2848 72292 2854
rect 72240 2790 72292 2796
rect 72252 800 72280 2790
rect 72436 800 72464 2858
rect 72528 2582 72556 6886
rect 72712 6118 72740 25162
rect 72804 24954 72832 25842
rect 72792 24948 72844 24954
rect 72792 24890 72844 24896
rect 72884 23520 72936 23526
rect 72884 23462 72936 23468
rect 72896 19922 72924 23462
rect 73264 19922 73292 34138
rect 73344 27532 73396 27538
rect 73344 27474 73396 27480
rect 72884 19916 72936 19922
rect 72884 19858 72936 19864
rect 73252 19916 73304 19922
rect 73252 19858 73304 19864
rect 73356 18426 73384 27474
rect 73448 19174 73476 34478
rect 73436 19168 73488 19174
rect 73436 19110 73488 19116
rect 73448 18902 73476 19110
rect 73436 18896 73488 18902
rect 73436 18838 73488 18844
rect 73344 18420 73396 18426
rect 73344 18362 73396 18368
rect 73540 6186 73568 37606
rect 73724 17678 73752 87246
rect 73816 86290 73844 89490
rect 73896 87372 73948 87378
rect 73896 87314 73948 87320
rect 73804 86284 73856 86290
rect 73804 86226 73856 86232
rect 73816 82006 73844 86226
rect 73804 82000 73856 82006
rect 73804 81942 73856 81948
rect 73804 81524 73856 81530
rect 73804 81466 73856 81472
rect 73816 35630 73844 81466
rect 73908 67386 73936 87314
rect 74080 81932 74132 81938
rect 74080 81874 74132 81880
rect 74092 80918 74120 81874
rect 74184 81530 74212 91666
rect 74356 91588 74408 91594
rect 74356 91530 74408 91536
rect 74368 90438 74396 91530
rect 74356 90432 74408 90438
rect 74356 90374 74408 90380
rect 74552 87378 74580 96426
rect 74632 89480 74684 89486
rect 74632 89422 74684 89428
rect 74540 87372 74592 87378
rect 74540 87314 74592 87320
rect 74644 86358 74672 89422
rect 74908 89412 74960 89418
rect 74908 89354 74960 89360
rect 74632 86352 74684 86358
rect 74632 86294 74684 86300
rect 74920 85338 74948 89354
rect 74908 85332 74960 85338
rect 74908 85274 74960 85280
rect 74172 81524 74224 81530
rect 74172 81466 74224 81472
rect 74080 80912 74132 80918
rect 74080 80854 74132 80860
rect 74540 72480 74592 72486
rect 74540 72422 74592 72428
rect 74080 67652 74132 67658
rect 74080 67594 74132 67600
rect 73896 67380 73948 67386
rect 73896 67322 73948 67328
rect 73908 47598 73936 67322
rect 73988 62348 74040 62354
rect 73988 62290 74040 62296
rect 74000 47802 74028 62290
rect 73988 47796 74040 47802
rect 73988 47738 74040 47744
rect 73896 47592 73948 47598
rect 73896 47534 73948 47540
rect 74000 35834 74028 47738
rect 74092 47190 74120 67594
rect 74448 62348 74500 62354
rect 74448 62290 74500 62296
rect 74264 62280 74316 62286
rect 74264 62222 74316 62228
rect 74080 47184 74132 47190
rect 74080 47126 74132 47132
rect 74276 46578 74304 62222
rect 74460 55214 74488 62290
rect 74368 55186 74488 55214
rect 74264 46572 74316 46578
rect 74264 46514 74316 46520
rect 74276 46374 74304 46514
rect 74264 46368 74316 46374
rect 74264 46310 74316 46316
rect 74264 45348 74316 45354
rect 74264 45290 74316 45296
rect 74276 45014 74304 45290
rect 74264 45008 74316 45014
rect 74264 44950 74316 44956
rect 74080 43988 74132 43994
rect 74080 43930 74132 43936
rect 74092 40526 74120 43930
rect 74368 41414 74396 55186
rect 74448 52556 74500 52562
rect 74448 52498 74500 52504
rect 74460 44946 74488 52498
rect 74448 44940 74500 44946
rect 74448 44882 74500 44888
rect 74460 42770 74488 44882
rect 74448 42764 74500 42770
rect 74448 42706 74500 42712
rect 74276 41386 74396 41414
rect 74080 40520 74132 40526
rect 74080 40462 74132 40468
rect 74092 37330 74120 40462
rect 74080 37324 74132 37330
rect 74080 37266 74132 37272
rect 74276 36174 74304 41386
rect 74448 38276 74500 38282
rect 74448 38218 74500 38224
rect 74460 37262 74488 38218
rect 74552 37330 74580 72422
rect 75196 71466 75224 97106
rect 76380 96960 76432 96966
rect 76380 96902 76432 96908
rect 75276 90024 75328 90030
rect 75276 89966 75328 89972
rect 75828 90024 75880 90030
rect 75828 89966 75880 89972
rect 75184 71460 75236 71466
rect 75184 71402 75236 71408
rect 75000 65612 75052 65618
rect 75000 65554 75052 65560
rect 75012 64122 75040 65554
rect 75000 64116 75052 64122
rect 75000 64058 75052 64064
rect 75012 61946 75040 64058
rect 75288 64054 75316 89966
rect 75736 89888 75788 89894
rect 75736 89830 75788 89836
rect 75368 87372 75420 87378
rect 75368 87314 75420 87320
rect 75380 70394 75408 87314
rect 75644 82952 75696 82958
rect 75644 82894 75696 82900
rect 75656 80102 75684 82894
rect 75644 80096 75696 80102
rect 75644 80038 75696 80044
rect 75380 70366 75500 70394
rect 75472 68202 75500 70366
rect 75460 68196 75512 68202
rect 75460 68138 75512 68144
rect 75368 64456 75420 64462
rect 75368 64398 75420 64404
rect 75276 64048 75328 64054
rect 75276 63990 75328 63996
rect 75000 61940 75052 61946
rect 75000 61882 75052 61888
rect 74816 61396 74868 61402
rect 74816 61338 74868 61344
rect 74828 60178 74856 61338
rect 75288 60734 75316 63990
rect 75380 63918 75408 64398
rect 75368 63912 75420 63918
rect 75368 63854 75420 63860
rect 75196 60706 75316 60734
rect 74816 60172 74868 60178
rect 74816 60114 74868 60120
rect 74828 58970 74856 60114
rect 74828 58942 75040 58970
rect 74816 55276 74868 55282
rect 74816 55218 74868 55224
rect 74632 44736 74684 44742
rect 74632 44678 74684 44684
rect 74540 37324 74592 37330
rect 74540 37266 74592 37272
rect 74448 37256 74500 37262
rect 74448 37198 74500 37204
rect 74264 36168 74316 36174
rect 74264 36110 74316 36116
rect 73988 35828 74040 35834
rect 73988 35770 74040 35776
rect 73804 35624 73856 35630
rect 73804 35566 73856 35572
rect 73816 35018 73844 35566
rect 73896 35488 73948 35494
rect 73896 35430 73948 35436
rect 73804 35012 73856 35018
rect 73804 34954 73856 34960
rect 73908 25770 73936 35430
rect 74276 34610 74304 36110
rect 74264 34604 74316 34610
rect 74264 34546 74316 34552
rect 74460 34066 74488 37198
rect 74448 34060 74500 34066
rect 74448 34002 74500 34008
rect 74460 27538 74488 34002
rect 74644 28082 74672 44678
rect 74828 41414 74856 55218
rect 74736 41386 74856 41414
rect 74736 38350 74764 41386
rect 74724 38344 74776 38350
rect 74724 38286 74776 38292
rect 75012 36718 75040 58942
rect 75196 50318 75224 60706
rect 75380 50454 75408 63854
rect 75472 61130 75500 68138
rect 75460 61124 75512 61130
rect 75460 61066 75512 61072
rect 75748 60314 75776 89830
rect 75840 64462 75868 89966
rect 76196 89956 76248 89962
rect 76196 89898 76248 89904
rect 76012 82952 76064 82958
rect 76012 82894 76064 82900
rect 76024 79558 76052 82894
rect 76012 79552 76064 79558
rect 76012 79494 76064 79500
rect 76208 67114 76236 89898
rect 76288 89888 76340 89894
rect 76288 89830 76340 89836
rect 76196 67108 76248 67114
rect 76196 67050 76248 67056
rect 75828 64456 75880 64462
rect 75828 64398 75880 64404
rect 75920 60648 75972 60654
rect 75920 60590 75972 60596
rect 75736 60308 75788 60314
rect 75736 60250 75788 60256
rect 75828 56228 75880 56234
rect 75828 56170 75880 56176
rect 75840 55282 75868 56170
rect 75828 55276 75880 55282
rect 75828 55218 75880 55224
rect 75368 50448 75420 50454
rect 75368 50390 75420 50396
rect 75184 50312 75236 50318
rect 75184 50254 75236 50260
rect 75828 46708 75880 46714
rect 75828 46650 75880 46656
rect 75840 36718 75868 46650
rect 75000 36712 75052 36718
rect 75000 36654 75052 36660
rect 75184 36712 75236 36718
rect 75184 36654 75236 36660
rect 75368 36712 75420 36718
rect 75368 36654 75420 36660
rect 75736 36712 75788 36718
rect 75736 36654 75788 36660
rect 75828 36712 75880 36718
rect 75828 36654 75880 36660
rect 75092 29096 75144 29102
rect 75092 29038 75144 29044
rect 74632 28076 74684 28082
rect 74632 28018 74684 28024
rect 74448 27532 74500 27538
rect 74448 27474 74500 27480
rect 75000 25832 75052 25838
rect 75000 25774 75052 25780
rect 73896 25764 73948 25770
rect 73896 25706 73948 25712
rect 73804 25152 73856 25158
rect 73804 25094 73856 25100
rect 73712 17672 73764 17678
rect 73712 17614 73764 17620
rect 73816 9450 73844 25094
rect 74172 20256 74224 20262
rect 74172 20198 74224 20204
rect 73804 9444 73856 9450
rect 73804 9386 73856 9392
rect 73528 6180 73580 6186
rect 73528 6122 73580 6128
rect 72700 6112 72752 6118
rect 72700 6054 72752 6060
rect 73712 5092 73764 5098
rect 73712 5034 73764 5040
rect 72608 4072 72660 4078
rect 72608 4014 72660 4020
rect 73252 4072 73304 4078
rect 73252 4014 73304 4020
rect 72516 2576 72568 2582
rect 72516 2518 72568 2524
rect 72620 800 72648 4014
rect 72792 3596 72844 3602
rect 72792 3538 72844 3544
rect 72804 800 72832 3538
rect 73068 2440 73120 2446
rect 73068 2382 73120 2388
rect 73080 800 73108 2382
rect 73264 800 73292 4014
rect 73436 2984 73488 2990
rect 73436 2926 73488 2932
rect 73448 800 73476 2926
rect 73620 2848 73672 2854
rect 73620 2790 73672 2796
rect 73632 800 73660 2790
rect 73724 2514 73752 5034
rect 73804 4684 73856 4690
rect 73804 4626 73856 4632
rect 73712 2508 73764 2514
rect 73712 2450 73764 2456
rect 73816 800 73844 4626
rect 74080 3596 74132 3602
rect 74080 3538 74132 3544
rect 74092 800 74120 3538
rect 74184 2650 74212 20198
rect 75012 14482 75040 25774
rect 75000 14476 75052 14482
rect 75000 14418 75052 14424
rect 75104 8430 75132 29038
rect 75196 10538 75224 36654
rect 75380 36310 75408 36654
rect 75748 36378 75776 36654
rect 75736 36372 75788 36378
rect 75736 36314 75788 36320
rect 75932 36310 75960 60590
rect 76104 53644 76156 53650
rect 76104 53586 76156 53592
rect 76012 47116 76064 47122
rect 76012 47058 76064 47064
rect 76024 46714 76052 47058
rect 76012 46708 76064 46714
rect 76012 46650 76064 46656
rect 76116 41414 76144 53586
rect 76196 49292 76248 49298
rect 76196 49234 76248 49240
rect 76024 41386 76144 41414
rect 76024 36378 76052 41386
rect 76208 36922 76236 49234
rect 76300 47122 76328 89830
rect 76288 47116 76340 47122
rect 76288 47058 76340 47064
rect 76392 37330 76420 96902
rect 76564 83020 76616 83026
rect 76564 82962 76616 82968
rect 76472 82952 76524 82958
rect 76472 82894 76524 82900
rect 76484 79762 76512 82894
rect 76472 79756 76524 79762
rect 76472 79698 76524 79704
rect 76576 73302 76604 82962
rect 76748 77920 76800 77926
rect 76748 77862 76800 77868
rect 76564 73296 76616 73302
rect 76564 73238 76616 73244
rect 76576 59090 76604 73238
rect 76656 67108 76708 67114
rect 76656 67050 76708 67056
rect 76668 61130 76696 67050
rect 76656 61124 76708 61130
rect 76656 61066 76708 61072
rect 76564 59084 76616 59090
rect 76564 59026 76616 59032
rect 76668 55826 76696 61066
rect 76656 55820 76708 55826
rect 76656 55762 76708 55768
rect 76668 55214 76696 55762
rect 76576 55186 76696 55214
rect 76380 37324 76432 37330
rect 76380 37266 76432 37272
rect 76196 36916 76248 36922
rect 76196 36858 76248 36864
rect 76012 36372 76064 36378
rect 76012 36314 76064 36320
rect 75368 36304 75420 36310
rect 75368 36246 75420 36252
rect 75920 36304 75972 36310
rect 75920 36246 75972 36252
rect 75920 25764 75972 25770
rect 75920 25706 75972 25712
rect 75932 25158 75960 25706
rect 75920 25152 75972 25158
rect 75920 25094 75972 25100
rect 76576 22166 76604 55186
rect 76760 54670 76788 77862
rect 76840 73636 76892 73642
rect 76840 73578 76892 73584
rect 76852 67250 76880 73578
rect 76932 73568 76984 73574
rect 76932 73510 76984 73516
rect 76840 67244 76892 67250
rect 76840 67186 76892 67192
rect 76944 60654 76972 73510
rect 77312 70378 77340 97106
rect 77772 96490 77800 99200
rect 78600 97152 78628 99200
rect 79520 97238 79548 99200
rect 79508 97232 79560 97238
rect 79508 97174 79560 97180
rect 78680 97164 78732 97170
rect 78600 97124 78680 97152
rect 78680 97106 78732 97112
rect 79968 97164 80020 97170
rect 79968 97106 80020 97112
rect 79140 97096 79192 97102
rect 79140 97038 79192 97044
rect 79152 96762 79180 97038
rect 79140 96756 79192 96762
rect 79140 96698 79192 96704
rect 77760 96484 77812 96490
rect 77760 96426 77812 96432
rect 77484 88256 77536 88262
rect 77484 88198 77536 88204
rect 77496 87854 77524 88198
rect 77668 87984 77720 87990
rect 77668 87926 77720 87932
rect 77484 87848 77536 87854
rect 77484 87790 77536 87796
rect 77576 87848 77628 87854
rect 77576 87790 77628 87796
rect 77680 87802 77708 87926
rect 77760 87848 77812 87854
rect 77680 87796 77760 87802
rect 77680 87790 77812 87796
rect 77588 87514 77616 87790
rect 77680 87774 77800 87790
rect 77576 87508 77628 87514
rect 77576 87450 77628 87456
rect 77680 84194 77708 87774
rect 79508 85128 79560 85134
rect 79508 85070 79560 85076
rect 77680 84166 77800 84194
rect 77300 70372 77352 70378
rect 77300 70314 77352 70320
rect 77208 69760 77260 69766
rect 77208 69702 77260 69708
rect 76932 60648 76984 60654
rect 76932 60590 76984 60596
rect 76748 54664 76800 54670
rect 76748 54606 76800 54612
rect 76656 47592 76708 47598
rect 76656 47534 76708 47540
rect 76668 25158 76696 47534
rect 77116 47116 77168 47122
rect 77116 47058 77168 47064
rect 76840 39636 76892 39642
rect 76840 39578 76892 39584
rect 76748 36304 76800 36310
rect 76748 36246 76800 36252
rect 76656 25152 76708 25158
rect 76656 25094 76708 25100
rect 76564 22160 76616 22166
rect 76564 22102 76616 22108
rect 76564 21616 76616 21622
rect 76564 21558 76616 21564
rect 75184 10532 75236 10538
rect 75184 10474 75236 10480
rect 75092 8424 75144 8430
rect 75092 8366 75144 8372
rect 74816 8084 74868 8090
rect 74816 8026 74868 8032
rect 74448 4072 74500 4078
rect 74448 4014 74500 4020
rect 74172 2644 74224 2650
rect 74172 2586 74224 2592
rect 74264 2508 74316 2514
rect 74264 2450 74316 2456
rect 74276 800 74304 2450
rect 74460 800 74488 4014
rect 74632 3596 74684 3602
rect 74632 3538 74684 3544
rect 74644 800 74672 3538
rect 74724 2848 74776 2854
rect 74724 2790 74776 2796
rect 74736 2310 74764 2790
rect 74828 2650 74856 8026
rect 75092 4072 75144 4078
rect 75736 4072 75788 4078
rect 75092 4014 75144 4020
rect 75656 4032 75736 4060
rect 74908 2916 74960 2922
rect 74908 2858 74960 2864
rect 74816 2644 74868 2650
rect 74816 2586 74868 2592
rect 74724 2304 74776 2310
rect 74724 2246 74776 2252
rect 74920 800 74948 2858
rect 75104 800 75132 4014
rect 75184 3460 75236 3466
rect 75184 3402 75236 3408
rect 75196 2990 75224 3402
rect 75184 2984 75236 2990
rect 75184 2926 75236 2932
rect 75276 2984 75328 2990
rect 75276 2926 75328 2932
rect 75288 800 75316 2926
rect 75460 2372 75512 2378
rect 75460 2314 75512 2320
rect 75472 800 75500 2314
rect 75656 800 75684 4032
rect 76380 4072 76432 4078
rect 75736 4014 75788 4020
rect 76300 4032 76380 4060
rect 75920 3596 75972 3602
rect 75920 3538 75972 3544
rect 75932 800 75960 3538
rect 76104 2848 76156 2854
rect 76104 2790 76156 2796
rect 76116 800 76144 2790
rect 76300 800 76328 4032
rect 76380 4014 76432 4020
rect 76472 3596 76524 3602
rect 76472 3538 76524 3544
rect 76484 800 76512 3538
rect 76576 2582 76604 21558
rect 76760 21554 76788 36246
rect 76748 21548 76800 21554
rect 76748 21490 76800 21496
rect 76852 2990 76880 39578
rect 76932 36372 76984 36378
rect 76932 36314 76984 36320
rect 76944 21622 76972 36314
rect 77128 26234 77156 47058
rect 77036 26206 77156 26234
rect 77036 24954 77064 26206
rect 77024 24948 77076 24954
rect 77024 24890 77076 24896
rect 76932 21616 76984 21622
rect 76932 21558 76984 21564
rect 77036 14414 77064 24890
rect 77024 14408 77076 14414
rect 77024 14350 77076 14356
rect 77116 12096 77168 12102
rect 77116 12038 77168 12044
rect 77128 11694 77156 12038
rect 77116 11688 77168 11694
rect 77116 11630 77168 11636
rect 77024 4072 77076 4078
rect 76944 4032 77024 4060
rect 76840 2984 76892 2990
rect 76840 2926 76892 2932
rect 76656 2916 76708 2922
rect 76656 2858 76708 2864
rect 76564 2576 76616 2582
rect 76564 2518 76616 2524
rect 76668 800 76696 2858
rect 76944 800 76972 4032
rect 77024 4014 77076 4020
rect 77116 3596 77168 3602
rect 77116 3538 77168 3544
rect 77128 800 77156 3538
rect 77220 2582 77248 69702
rect 77312 65958 77340 70314
rect 77300 65952 77352 65958
rect 77300 65894 77352 65900
rect 77484 55888 77536 55894
rect 77484 55830 77536 55836
rect 77300 47592 77352 47598
rect 77300 47534 77352 47540
rect 77312 47190 77340 47534
rect 77300 47184 77352 47190
rect 77300 47126 77352 47132
rect 77300 2848 77352 2854
rect 77300 2790 77352 2796
rect 77312 2582 77340 2790
rect 77496 2650 77524 55830
rect 77668 45824 77720 45830
rect 77668 45766 77720 45772
rect 77680 45558 77708 45766
rect 77668 45552 77720 45558
rect 77668 45494 77720 45500
rect 77668 40384 77720 40390
rect 77668 40326 77720 40332
rect 77680 40186 77708 40326
rect 77668 40180 77720 40186
rect 77668 40122 77720 40128
rect 77576 38208 77628 38214
rect 77576 38150 77628 38156
rect 77588 27402 77616 38150
rect 77772 30258 77800 84166
rect 79324 84040 79376 84046
rect 79324 83982 79376 83988
rect 79336 83706 79364 83982
rect 79324 83700 79376 83706
rect 79324 83642 79376 83648
rect 78128 79688 78180 79694
rect 78128 79630 78180 79636
rect 78140 77042 78168 79630
rect 78128 77036 78180 77042
rect 78128 76978 78180 76984
rect 78140 74534 78168 76978
rect 79416 76832 79468 76838
rect 79416 76774 79468 76780
rect 79324 74724 79376 74730
rect 79324 74666 79376 74672
rect 78312 74656 78364 74662
rect 78312 74598 78364 74604
rect 78140 74506 78260 74534
rect 78232 68882 78260 74506
rect 78324 74322 78352 74598
rect 78312 74316 78364 74322
rect 78312 74258 78364 74264
rect 78496 74248 78548 74254
rect 78496 74190 78548 74196
rect 78508 73778 78536 74190
rect 78496 73772 78548 73778
rect 78496 73714 78548 73720
rect 78588 72616 78640 72622
rect 78588 72558 78640 72564
rect 78600 71942 78628 72558
rect 78680 72140 78732 72146
rect 78680 72082 78732 72088
rect 78692 71942 78720 72082
rect 78864 72072 78916 72078
rect 78864 72014 78916 72020
rect 78588 71936 78640 71942
rect 78588 71878 78640 71884
rect 78680 71936 78732 71942
rect 78680 71878 78732 71884
rect 78692 69970 78720 71878
rect 78680 69964 78732 69970
rect 78680 69906 78732 69912
rect 78312 69012 78364 69018
rect 78312 68954 78364 68960
rect 78220 68876 78272 68882
rect 78220 68818 78272 68824
rect 78324 68814 78352 68954
rect 78496 68876 78548 68882
rect 78496 68818 78548 68824
rect 78312 68808 78364 68814
rect 78312 68750 78364 68756
rect 77944 66496 77996 66502
rect 77944 66438 77996 66444
rect 77956 61878 77984 66438
rect 77944 61872 77996 61878
rect 77944 61814 77996 61820
rect 78324 60734 78352 68750
rect 78232 60706 78352 60734
rect 78128 54664 78180 54670
rect 78128 54606 78180 54612
rect 78036 49224 78088 49230
rect 78036 49166 78088 49172
rect 77852 45620 77904 45626
rect 77852 45562 77904 45568
rect 77864 45490 77892 45562
rect 77852 45484 77904 45490
rect 77852 45426 77904 45432
rect 78048 37262 78076 49166
rect 78140 43994 78168 54606
rect 78128 43988 78180 43994
rect 78128 43930 78180 43936
rect 78036 37256 78088 37262
rect 78036 37198 78088 37204
rect 77944 36168 77996 36174
rect 77944 36110 77996 36116
rect 77956 31754 77984 36110
rect 77864 31726 77984 31754
rect 77864 31346 77892 31726
rect 77852 31340 77904 31346
rect 77852 31282 77904 31288
rect 77760 30252 77812 30258
rect 77760 30194 77812 30200
rect 77668 28620 77720 28626
rect 77668 28562 77720 28568
rect 77680 28422 77708 28562
rect 77944 28552 77996 28558
rect 77944 28494 77996 28500
rect 77668 28416 77720 28422
rect 77668 28358 77720 28364
rect 77576 27396 77628 27402
rect 77576 27338 77628 27344
rect 77680 21146 77708 28358
rect 77956 28218 77984 28494
rect 77944 28212 77996 28218
rect 77944 28154 77996 28160
rect 78048 26234 78076 37198
rect 78232 29170 78260 60706
rect 78312 39568 78364 39574
rect 78312 39510 78364 39516
rect 78324 36242 78352 39510
rect 78404 39364 78456 39370
rect 78404 39306 78456 39312
rect 78416 38010 78444 39306
rect 78404 38004 78456 38010
rect 78404 37946 78456 37952
rect 78312 36236 78364 36242
rect 78312 36178 78364 36184
rect 78508 30258 78536 68818
rect 78772 68740 78824 68746
rect 78772 68682 78824 68688
rect 78588 58948 78640 58954
rect 78588 58890 78640 58896
rect 78600 37806 78628 58890
rect 78680 42764 78732 42770
rect 78680 42706 78732 42712
rect 78692 42090 78720 42706
rect 78680 42084 78732 42090
rect 78680 42026 78732 42032
rect 78588 37800 78640 37806
rect 78588 37742 78640 37748
rect 78496 30252 78548 30258
rect 78496 30194 78548 30200
rect 78784 29306 78812 68682
rect 78876 66094 78904 72014
rect 79336 67046 79364 74666
rect 79324 67040 79376 67046
rect 79324 66982 79376 66988
rect 78864 66088 78916 66094
rect 78864 66030 78916 66036
rect 78876 63850 78904 66030
rect 78864 63844 78916 63850
rect 78864 63786 78916 63792
rect 79324 61056 79376 61062
rect 79324 60998 79376 61004
rect 78956 54596 79008 54602
rect 78956 54538 79008 54544
rect 78968 37874 78996 54538
rect 78956 37868 79008 37874
rect 78956 37810 79008 37816
rect 78864 37800 78916 37806
rect 78864 37742 78916 37748
rect 79140 37800 79192 37806
rect 79140 37742 79192 37748
rect 78772 29300 78824 29306
rect 78772 29242 78824 29248
rect 78220 29164 78272 29170
rect 78220 29106 78272 29112
rect 78220 27396 78272 27402
rect 78220 27338 78272 27344
rect 77864 26206 78076 26234
rect 77864 23662 77892 26206
rect 78232 25294 78260 27338
rect 78220 25288 78272 25294
rect 78220 25230 78272 25236
rect 78496 25288 78548 25294
rect 78496 25230 78548 25236
rect 77852 23656 77904 23662
rect 77852 23598 77904 23604
rect 78232 23186 78260 25230
rect 78220 23180 78272 23186
rect 78220 23122 78272 23128
rect 77944 23112 77996 23118
rect 77944 23054 77996 23060
rect 77668 21140 77720 21146
rect 77668 21082 77720 21088
rect 77668 21004 77720 21010
rect 77668 20946 77720 20952
rect 77680 17610 77708 20946
rect 77956 18698 77984 23054
rect 78128 20392 78180 20398
rect 78128 20334 78180 20340
rect 77944 18692 77996 18698
rect 77944 18634 77996 18640
rect 77668 17604 77720 17610
rect 77668 17546 77720 17552
rect 78036 6656 78088 6662
rect 78036 6598 78088 6604
rect 78048 6458 78076 6598
rect 78036 6452 78088 6458
rect 78036 6394 78088 6400
rect 78140 4162 78168 20334
rect 78508 7818 78536 25230
rect 78772 23316 78824 23322
rect 78772 23258 78824 23264
rect 78496 7812 78548 7818
rect 78496 7754 78548 7760
rect 78784 6914 78812 23258
rect 78876 10742 78904 37742
rect 78864 10736 78916 10742
rect 78864 10678 78916 10684
rect 79152 8022 79180 37742
rect 79232 37664 79284 37670
rect 79232 37606 79284 37612
rect 79140 8016 79192 8022
rect 79140 7958 79192 7964
rect 79244 7886 79272 37606
rect 79232 7880 79284 7886
rect 79232 7822 79284 7828
rect 78784 6886 78904 6914
rect 78772 4684 78824 4690
rect 78772 4626 78824 4632
rect 78048 4134 78168 4162
rect 77668 4072 77720 4078
rect 77588 4032 77668 4060
rect 77484 2644 77536 2650
rect 77484 2586 77536 2592
rect 77208 2576 77260 2582
rect 77208 2518 77260 2524
rect 77300 2576 77352 2582
rect 77300 2518 77352 2524
rect 77300 2440 77352 2446
rect 77300 2382 77352 2388
rect 77312 800 77340 2382
rect 77588 2122 77616 4032
rect 77668 4014 77720 4020
rect 77760 3596 77812 3602
rect 77496 2094 77616 2122
rect 77680 3556 77760 3584
rect 77496 800 77524 2094
rect 77680 800 77708 3556
rect 77760 3538 77812 3544
rect 78048 2922 78076 4134
rect 78128 4004 78180 4010
rect 78128 3946 78180 3952
rect 77944 2916 77996 2922
rect 77944 2858 77996 2864
rect 78036 2916 78088 2922
rect 78036 2858 78088 2864
rect 77956 800 77984 2858
rect 78140 800 78168 3946
rect 78220 3936 78272 3942
rect 78220 3878 78272 3884
rect 78232 2990 78260 3878
rect 78404 3596 78456 3602
rect 78324 3556 78404 3584
rect 78220 2984 78272 2990
rect 78220 2926 78272 2932
rect 78324 800 78352 3556
rect 78404 3538 78456 3544
rect 78496 2372 78548 2378
rect 78496 2314 78548 2320
rect 78508 800 78536 2314
rect 78784 800 78812 4626
rect 78876 2650 78904 6886
rect 79336 4826 79364 60998
rect 79428 41414 79456 76774
rect 79520 46918 79548 85070
rect 79784 76560 79836 76566
rect 79784 76502 79836 76508
rect 79600 67040 79652 67046
rect 79600 66982 79652 66988
rect 79612 51074 79640 66982
rect 79692 63232 79744 63238
rect 79692 63174 79744 63180
rect 79704 54738 79732 63174
rect 79796 55214 79824 76502
rect 79980 72486 80008 97106
rect 80348 96626 80376 99200
rect 81268 97594 81296 99200
rect 81268 97566 81388 97594
rect 81020 97404 81316 97424
rect 81076 97402 81100 97404
rect 81156 97402 81180 97404
rect 81236 97402 81260 97404
rect 81098 97350 81100 97402
rect 81162 97350 81174 97402
rect 81236 97350 81238 97402
rect 81076 97348 81100 97350
rect 81156 97348 81180 97350
rect 81236 97348 81260 97350
rect 81020 97328 81316 97348
rect 80704 97028 80756 97034
rect 80704 96970 80756 96976
rect 80336 96620 80388 96626
rect 80336 96562 80388 96568
rect 79968 72480 80020 72486
rect 79968 72422 80020 72428
rect 79980 72282 80008 72422
rect 79968 72276 80020 72282
rect 79968 72218 80020 72224
rect 80244 71936 80296 71942
rect 80244 71878 80296 71884
rect 80256 64598 80284 71878
rect 80716 68338 80744 96970
rect 81360 96558 81388 97566
rect 82096 97238 82124 99200
rect 82924 97322 82952 99200
rect 82924 97294 83044 97322
rect 82084 97232 82136 97238
rect 82084 97174 82136 97180
rect 82176 97164 82228 97170
rect 82176 97106 82228 97112
rect 82912 97164 82964 97170
rect 82912 97106 82964 97112
rect 81348 96552 81400 96558
rect 81348 96494 81400 96500
rect 81440 96416 81492 96422
rect 81440 96358 81492 96364
rect 81020 96316 81316 96336
rect 81076 96314 81100 96316
rect 81156 96314 81180 96316
rect 81236 96314 81260 96316
rect 81098 96262 81100 96314
rect 81162 96262 81174 96314
rect 81236 96262 81238 96314
rect 81076 96260 81100 96262
rect 81156 96260 81180 96262
rect 81236 96260 81260 96262
rect 81020 96240 81316 96260
rect 81020 95228 81316 95248
rect 81076 95226 81100 95228
rect 81156 95226 81180 95228
rect 81236 95226 81260 95228
rect 81098 95174 81100 95226
rect 81162 95174 81174 95226
rect 81236 95174 81238 95226
rect 81076 95172 81100 95174
rect 81156 95172 81180 95174
rect 81236 95172 81260 95174
rect 81020 95152 81316 95172
rect 81020 94140 81316 94160
rect 81076 94138 81100 94140
rect 81156 94138 81180 94140
rect 81236 94138 81260 94140
rect 81098 94086 81100 94138
rect 81162 94086 81174 94138
rect 81236 94086 81238 94138
rect 81076 94084 81100 94086
rect 81156 94084 81180 94086
rect 81236 94084 81260 94086
rect 81020 94064 81316 94084
rect 81020 93052 81316 93072
rect 81076 93050 81100 93052
rect 81156 93050 81180 93052
rect 81236 93050 81260 93052
rect 81098 92998 81100 93050
rect 81162 92998 81174 93050
rect 81236 92998 81238 93050
rect 81076 92996 81100 92998
rect 81156 92996 81180 92998
rect 81236 92996 81260 92998
rect 81020 92976 81316 92996
rect 81020 91964 81316 91984
rect 81076 91962 81100 91964
rect 81156 91962 81180 91964
rect 81236 91962 81260 91964
rect 81098 91910 81100 91962
rect 81162 91910 81174 91962
rect 81236 91910 81238 91962
rect 81076 91908 81100 91910
rect 81156 91908 81180 91910
rect 81236 91908 81260 91910
rect 81020 91888 81316 91908
rect 81020 90876 81316 90896
rect 81076 90874 81100 90876
rect 81156 90874 81180 90876
rect 81236 90874 81260 90876
rect 81098 90822 81100 90874
rect 81162 90822 81174 90874
rect 81236 90822 81238 90874
rect 81076 90820 81100 90822
rect 81156 90820 81180 90822
rect 81236 90820 81260 90822
rect 81020 90800 81316 90820
rect 81020 89788 81316 89808
rect 81076 89786 81100 89788
rect 81156 89786 81180 89788
rect 81236 89786 81260 89788
rect 81098 89734 81100 89786
rect 81162 89734 81174 89786
rect 81236 89734 81238 89786
rect 81076 89732 81100 89734
rect 81156 89732 81180 89734
rect 81236 89732 81260 89734
rect 81020 89712 81316 89732
rect 81452 89554 81480 96358
rect 81440 89548 81492 89554
rect 81440 89490 81492 89496
rect 82188 89010 82216 97106
rect 82820 96960 82872 96966
rect 82820 96902 82872 96908
rect 82832 96490 82860 96902
rect 82820 96484 82872 96490
rect 82820 96426 82872 96432
rect 82176 89004 82228 89010
rect 82176 88946 82228 88952
rect 81020 88700 81316 88720
rect 81076 88698 81100 88700
rect 81156 88698 81180 88700
rect 81236 88698 81260 88700
rect 81098 88646 81100 88698
rect 81162 88646 81174 88698
rect 81236 88646 81238 88698
rect 81076 88644 81100 88646
rect 81156 88644 81180 88646
rect 81236 88644 81260 88646
rect 81020 88624 81316 88644
rect 81020 87612 81316 87632
rect 81076 87610 81100 87612
rect 81156 87610 81180 87612
rect 81236 87610 81260 87612
rect 81098 87558 81100 87610
rect 81162 87558 81174 87610
rect 81236 87558 81238 87610
rect 81076 87556 81100 87558
rect 81156 87556 81180 87558
rect 81236 87556 81260 87558
rect 81020 87536 81316 87556
rect 81020 86524 81316 86544
rect 81076 86522 81100 86524
rect 81156 86522 81180 86524
rect 81236 86522 81260 86524
rect 81098 86470 81100 86522
rect 81162 86470 81174 86522
rect 81236 86470 81238 86522
rect 81076 86468 81100 86470
rect 81156 86468 81180 86470
rect 81236 86468 81260 86470
rect 81020 86448 81316 86468
rect 82820 86080 82872 86086
rect 82820 86022 82872 86028
rect 82084 85672 82136 85678
rect 82084 85614 82136 85620
rect 81020 85436 81316 85456
rect 81076 85434 81100 85436
rect 81156 85434 81180 85436
rect 81236 85434 81260 85436
rect 81098 85382 81100 85434
rect 81162 85382 81174 85434
rect 81236 85382 81238 85434
rect 81076 85380 81100 85382
rect 81156 85380 81180 85382
rect 81236 85380 81260 85382
rect 81020 85360 81316 85380
rect 81020 84348 81316 84368
rect 81076 84346 81100 84348
rect 81156 84346 81180 84348
rect 81236 84346 81260 84348
rect 81098 84294 81100 84346
rect 81162 84294 81174 84346
rect 81236 84294 81238 84346
rect 81076 84292 81100 84294
rect 81156 84292 81180 84294
rect 81236 84292 81260 84294
rect 81020 84272 81316 84292
rect 81020 83260 81316 83280
rect 81076 83258 81100 83260
rect 81156 83258 81180 83260
rect 81236 83258 81260 83260
rect 81098 83206 81100 83258
rect 81162 83206 81174 83258
rect 81236 83206 81238 83258
rect 81076 83204 81100 83206
rect 81156 83204 81180 83206
rect 81236 83204 81260 83206
rect 81020 83184 81316 83204
rect 81020 82172 81316 82192
rect 81076 82170 81100 82172
rect 81156 82170 81180 82172
rect 81236 82170 81260 82172
rect 81098 82118 81100 82170
rect 81162 82118 81174 82170
rect 81236 82118 81238 82170
rect 81076 82116 81100 82118
rect 81156 82116 81180 82118
rect 81236 82116 81260 82118
rect 81020 82096 81316 82116
rect 81020 81084 81316 81104
rect 81076 81082 81100 81084
rect 81156 81082 81180 81084
rect 81236 81082 81260 81084
rect 81098 81030 81100 81082
rect 81162 81030 81174 81082
rect 81236 81030 81238 81082
rect 81076 81028 81100 81030
rect 81156 81028 81180 81030
rect 81236 81028 81260 81030
rect 81020 81008 81316 81028
rect 81020 79996 81316 80016
rect 81076 79994 81100 79996
rect 81156 79994 81180 79996
rect 81236 79994 81260 79996
rect 81098 79942 81100 79994
rect 81162 79942 81174 79994
rect 81236 79942 81238 79994
rect 81076 79940 81100 79942
rect 81156 79940 81180 79942
rect 81236 79940 81260 79942
rect 81020 79920 81316 79940
rect 80796 79620 80848 79626
rect 80796 79562 80848 79568
rect 80808 77110 80836 79562
rect 81020 78908 81316 78928
rect 81076 78906 81100 78908
rect 81156 78906 81180 78908
rect 81236 78906 81260 78908
rect 81098 78854 81100 78906
rect 81162 78854 81174 78906
rect 81236 78854 81238 78906
rect 81076 78852 81100 78854
rect 81156 78852 81180 78854
rect 81236 78852 81260 78854
rect 81020 78832 81316 78852
rect 81020 77820 81316 77840
rect 81076 77818 81100 77820
rect 81156 77818 81180 77820
rect 81236 77818 81260 77820
rect 81098 77766 81100 77818
rect 81162 77766 81174 77818
rect 81236 77766 81238 77818
rect 81076 77764 81100 77766
rect 81156 77764 81180 77766
rect 81236 77764 81260 77766
rect 81020 77744 81316 77764
rect 80796 77104 80848 77110
rect 80796 77046 80848 77052
rect 80808 68814 80836 77046
rect 81020 76732 81316 76752
rect 81076 76730 81100 76732
rect 81156 76730 81180 76732
rect 81236 76730 81260 76732
rect 81098 76678 81100 76730
rect 81162 76678 81174 76730
rect 81236 76678 81238 76730
rect 81076 76676 81100 76678
rect 81156 76676 81180 76678
rect 81236 76676 81260 76678
rect 81020 76656 81316 76676
rect 81020 75644 81316 75664
rect 81076 75642 81100 75644
rect 81156 75642 81180 75644
rect 81236 75642 81260 75644
rect 81098 75590 81100 75642
rect 81162 75590 81174 75642
rect 81236 75590 81238 75642
rect 81076 75588 81100 75590
rect 81156 75588 81180 75590
rect 81236 75588 81260 75590
rect 81020 75568 81316 75588
rect 81020 74556 81316 74576
rect 81076 74554 81100 74556
rect 81156 74554 81180 74556
rect 81236 74554 81260 74556
rect 81098 74502 81100 74554
rect 81162 74502 81174 74554
rect 81236 74502 81238 74554
rect 81076 74500 81100 74502
rect 81156 74500 81180 74502
rect 81236 74500 81260 74502
rect 81020 74480 81316 74500
rect 81020 73468 81316 73488
rect 81076 73466 81100 73468
rect 81156 73466 81180 73468
rect 81236 73466 81260 73468
rect 81098 73414 81100 73466
rect 81162 73414 81174 73466
rect 81236 73414 81238 73466
rect 81076 73412 81100 73414
rect 81156 73412 81180 73414
rect 81236 73412 81260 73414
rect 81020 73392 81316 73412
rect 81020 72380 81316 72400
rect 81076 72378 81100 72380
rect 81156 72378 81180 72380
rect 81236 72378 81260 72380
rect 81098 72326 81100 72378
rect 81162 72326 81174 72378
rect 81236 72326 81238 72378
rect 81076 72324 81100 72326
rect 81156 72324 81180 72326
rect 81236 72324 81260 72326
rect 81020 72304 81316 72324
rect 81020 71292 81316 71312
rect 81076 71290 81100 71292
rect 81156 71290 81180 71292
rect 81236 71290 81260 71292
rect 81098 71238 81100 71290
rect 81162 71238 81174 71290
rect 81236 71238 81238 71290
rect 81076 71236 81100 71238
rect 81156 71236 81180 71238
rect 81236 71236 81260 71238
rect 81020 71216 81316 71236
rect 81020 70204 81316 70224
rect 81076 70202 81100 70204
rect 81156 70202 81180 70204
rect 81236 70202 81260 70204
rect 81098 70150 81100 70202
rect 81162 70150 81174 70202
rect 81236 70150 81238 70202
rect 81076 70148 81100 70150
rect 81156 70148 81180 70150
rect 81236 70148 81260 70150
rect 81020 70128 81316 70148
rect 81020 69116 81316 69136
rect 81076 69114 81100 69116
rect 81156 69114 81180 69116
rect 81236 69114 81260 69116
rect 81098 69062 81100 69114
rect 81162 69062 81174 69114
rect 81236 69062 81238 69114
rect 81076 69060 81100 69062
rect 81156 69060 81180 69062
rect 81236 69060 81260 69062
rect 81020 69040 81316 69060
rect 80796 68808 80848 68814
rect 80796 68750 80848 68756
rect 80704 68332 80756 68338
rect 80704 68274 80756 68280
rect 80520 66088 80572 66094
rect 80520 66030 80572 66036
rect 80336 65204 80388 65210
rect 80336 65146 80388 65152
rect 80348 64874 80376 65146
rect 80348 64846 80468 64874
rect 80244 64592 80296 64598
rect 80244 64534 80296 64540
rect 80152 60716 80204 60722
rect 80152 60658 80204 60664
rect 80164 59158 80192 60658
rect 80440 60178 80468 64846
rect 80428 60172 80480 60178
rect 80428 60114 80480 60120
rect 80152 59152 80204 59158
rect 80152 59094 80204 59100
rect 79796 55186 80008 55214
rect 79692 54732 79744 54738
rect 79692 54674 79744 54680
rect 79980 53650 80008 55186
rect 79968 53644 80020 53650
rect 79968 53586 80020 53592
rect 79612 51046 79732 51074
rect 79508 46912 79560 46918
rect 79508 46854 79560 46860
rect 79428 41386 79548 41414
rect 79416 22976 79468 22982
rect 79416 22918 79468 22924
rect 79428 22506 79456 22918
rect 79520 22710 79548 41386
rect 79704 37330 79732 51046
rect 79980 42770 80008 53586
rect 80164 52562 80192 59094
rect 80440 55842 80468 60114
rect 80532 55962 80560 66030
rect 80520 55956 80572 55962
rect 80520 55898 80572 55904
rect 80440 55814 80560 55842
rect 80532 52562 80560 55814
rect 80612 55752 80664 55758
rect 80612 55694 80664 55700
rect 80152 52556 80204 52562
rect 80152 52498 80204 52504
rect 80520 52556 80572 52562
rect 80520 52498 80572 52504
rect 80520 51876 80572 51882
rect 80520 51818 80572 51824
rect 80532 45554 80560 51818
rect 80256 45526 80560 45554
rect 79968 42764 80020 42770
rect 79968 42706 80020 42712
rect 80060 41812 80112 41818
rect 80060 41754 80112 41760
rect 80072 41478 80100 41754
rect 80060 41472 80112 41478
rect 80060 41414 80112 41420
rect 79692 37324 79744 37330
rect 79692 37266 79744 37272
rect 79600 25152 79652 25158
rect 79600 25094 79652 25100
rect 79508 22704 79560 22710
rect 79508 22646 79560 22652
rect 79416 22500 79468 22506
rect 79416 22442 79468 22448
rect 79428 18902 79456 22442
rect 79416 18896 79468 18902
rect 79416 18838 79468 18844
rect 79612 18170 79640 25094
rect 79428 18142 79640 18170
rect 79428 16590 79456 18142
rect 79416 16584 79468 16590
rect 79416 16526 79468 16532
rect 79428 15910 79456 16526
rect 79416 15904 79468 15910
rect 79416 15846 79468 15852
rect 79508 9376 79560 9382
rect 79508 9318 79560 9324
rect 79324 4820 79376 4826
rect 79324 4762 79376 4768
rect 79324 4684 79376 4690
rect 79324 4626 79376 4632
rect 79048 3596 79100 3602
rect 78968 3556 79048 3584
rect 78864 2644 78916 2650
rect 78864 2586 78916 2592
rect 78968 800 78996 3556
rect 79048 3538 79100 3544
rect 79232 2848 79284 2854
rect 79232 2790 79284 2796
rect 79244 1442 79272 2790
rect 79152 1414 79272 1442
rect 79152 800 79180 1414
rect 79336 800 79364 4626
rect 79520 2650 79548 9318
rect 79704 7886 79732 37266
rect 80256 31754 80284 45526
rect 80428 41812 80480 41818
rect 80428 41754 80480 41760
rect 80072 31726 80284 31754
rect 80440 31754 80468 41754
rect 80440 31726 80560 31754
rect 80072 24070 80100 31726
rect 80152 25900 80204 25906
rect 80152 25842 80204 25848
rect 80164 25430 80192 25842
rect 80152 25424 80204 25430
rect 80152 25366 80204 25372
rect 80244 25288 80296 25294
rect 80244 25230 80296 25236
rect 80256 24954 80284 25230
rect 80244 24948 80296 24954
rect 80244 24890 80296 24896
rect 80060 24064 80112 24070
rect 80060 24006 80112 24012
rect 79876 17264 79928 17270
rect 80152 17264 80204 17270
rect 79928 17212 80152 17218
rect 79876 17206 80204 17212
rect 79888 17190 80192 17206
rect 80336 15972 80388 15978
rect 80336 15914 80388 15920
rect 79692 7880 79744 7886
rect 79692 7822 79744 7828
rect 80244 5704 80296 5710
rect 80244 5646 80296 5652
rect 80152 4752 80204 4758
rect 80152 4694 80204 4700
rect 80060 4684 80112 4690
rect 80060 4626 80112 4632
rect 79692 3596 79744 3602
rect 79612 3556 79692 3584
rect 79508 2644 79560 2650
rect 79508 2586 79560 2592
rect 79612 1850 79640 3556
rect 79692 3538 79744 3544
rect 79968 3528 80020 3534
rect 79968 3470 80020 3476
rect 79980 3058 80008 3470
rect 79968 3052 80020 3058
rect 79968 2994 80020 3000
rect 79784 2916 79836 2922
rect 79784 2858 79836 2864
rect 79520 1822 79640 1850
rect 79520 800 79548 1822
rect 79796 800 79824 2858
rect 80072 2802 80100 4626
rect 80164 3618 80192 4694
rect 80256 4078 80284 5646
rect 80348 4078 80376 15914
rect 80532 11830 80560 31726
rect 80624 21486 80652 55694
rect 80704 53032 80756 53038
rect 80704 52974 80756 52980
rect 80716 42634 80744 52974
rect 80704 42628 80756 42634
rect 80704 42570 80756 42576
rect 80808 24750 80836 68750
rect 81020 68028 81316 68048
rect 81076 68026 81100 68028
rect 81156 68026 81180 68028
rect 81236 68026 81260 68028
rect 81098 67974 81100 68026
rect 81162 67974 81174 68026
rect 81236 67974 81238 68026
rect 81076 67972 81100 67974
rect 81156 67972 81180 67974
rect 81236 67972 81260 67974
rect 81020 67952 81316 67972
rect 81020 66940 81316 66960
rect 81076 66938 81100 66940
rect 81156 66938 81180 66940
rect 81236 66938 81260 66940
rect 81098 66886 81100 66938
rect 81162 66886 81174 66938
rect 81236 66886 81238 66938
rect 81076 66884 81100 66886
rect 81156 66884 81180 66886
rect 81236 66884 81260 66886
rect 81020 66864 81316 66884
rect 81992 66088 82044 66094
rect 81992 66030 82044 66036
rect 81020 65852 81316 65872
rect 81076 65850 81100 65852
rect 81156 65850 81180 65852
rect 81236 65850 81260 65852
rect 81098 65798 81100 65850
rect 81162 65798 81174 65850
rect 81236 65798 81238 65850
rect 81076 65796 81100 65798
rect 81156 65796 81180 65798
rect 81236 65796 81260 65798
rect 81020 65776 81316 65796
rect 80888 65068 80940 65074
rect 80888 65010 80940 65016
rect 80900 60586 80928 65010
rect 81716 64864 81768 64870
rect 81716 64806 81768 64812
rect 81020 64764 81316 64784
rect 81076 64762 81100 64764
rect 81156 64762 81180 64764
rect 81236 64762 81260 64764
rect 81098 64710 81100 64762
rect 81162 64710 81174 64762
rect 81236 64710 81238 64762
rect 81076 64708 81100 64710
rect 81156 64708 81180 64710
rect 81236 64708 81260 64710
rect 81020 64688 81316 64708
rect 81728 63850 81756 64806
rect 81716 63844 81768 63850
rect 81716 63786 81768 63792
rect 81020 63676 81316 63696
rect 81076 63674 81100 63676
rect 81156 63674 81180 63676
rect 81236 63674 81260 63676
rect 81098 63622 81100 63674
rect 81162 63622 81174 63674
rect 81236 63622 81238 63674
rect 81076 63620 81100 63622
rect 81156 63620 81180 63622
rect 81236 63620 81260 63622
rect 81020 63600 81316 63620
rect 81020 62588 81316 62608
rect 81076 62586 81100 62588
rect 81156 62586 81180 62588
rect 81236 62586 81260 62588
rect 81098 62534 81100 62586
rect 81162 62534 81174 62586
rect 81236 62534 81238 62586
rect 81076 62532 81100 62534
rect 81156 62532 81180 62534
rect 81236 62532 81260 62534
rect 81020 62512 81316 62532
rect 81020 61500 81316 61520
rect 81076 61498 81100 61500
rect 81156 61498 81180 61500
rect 81236 61498 81260 61500
rect 81098 61446 81100 61498
rect 81162 61446 81174 61498
rect 81236 61446 81238 61498
rect 81076 61444 81100 61446
rect 81156 61444 81180 61446
rect 81236 61444 81260 61446
rect 81020 61424 81316 61444
rect 80888 60580 80940 60586
rect 80888 60522 80940 60528
rect 80900 52562 80928 60522
rect 81020 60412 81316 60432
rect 81076 60410 81100 60412
rect 81156 60410 81180 60412
rect 81236 60410 81260 60412
rect 81098 60358 81100 60410
rect 81162 60358 81174 60410
rect 81236 60358 81238 60410
rect 81076 60356 81100 60358
rect 81156 60356 81180 60358
rect 81236 60356 81260 60358
rect 81020 60336 81316 60356
rect 81020 59324 81316 59344
rect 81076 59322 81100 59324
rect 81156 59322 81180 59324
rect 81236 59322 81260 59324
rect 81098 59270 81100 59322
rect 81162 59270 81174 59322
rect 81236 59270 81238 59322
rect 81076 59268 81100 59270
rect 81156 59268 81180 59270
rect 81236 59268 81260 59270
rect 81020 59248 81316 59268
rect 81348 58336 81400 58342
rect 81348 58278 81400 58284
rect 81020 58236 81316 58256
rect 81076 58234 81100 58236
rect 81156 58234 81180 58236
rect 81236 58234 81260 58236
rect 81098 58182 81100 58234
rect 81162 58182 81174 58234
rect 81236 58182 81238 58234
rect 81076 58180 81100 58182
rect 81156 58180 81180 58182
rect 81236 58180 81260 58182
rect 81020 58160 81316 58180
rect 81020 57148 81316 57168
rect 81076 57146 81100 57148
rect 81156 57146 81180 57148
rect 81236 57146 81260 57148
rect 81098 57094 81100 57146
rect 81162 57094 81174 57146
rect 81236 57094 81238 57146
rect 81076 57092 81100 57094
rect 81156 57092 81180 57094
rect 81236 57092 81260 57094
rect 81020 57072 81316 57092
rect 81020 56060 81316 56080
rect 81076 56058 81100 56060
rect 81156 56058 81180 56060
rect 81236 56058 81260 56060
rect 81098 56006 81100 56058
rect 81162 56006 81174 56058
rect 81236 56006 81238 56058
rect 81076 56004 81100 56006
rect 81156 56004 81180 56006
rect 81236 56004 81260 56006
rect 81020 55984 81316 56004
rect 81020 54972 81316 54992
rect 81076 54970 81100 54972
rect 81156 54970 81180 54972
rect 81236 54970 81260 54972
rect 81098 54918 81100 54970
rect 81162 54918 81174 54970
rect 81236 54918 81238 54970
rect 81076 54916 81100 54918
rect 81156 54916 81180 54918
rect 81236 54916 81260 54918
rect 81020 54896 81316 54916
rect 81020 53884 81316 53904
rect 81076 53882 81100 53884
rect 81156 53882 81180 53884
rect 81236 53882 81260 53884
rect 81098 53830 81100 53882
rect 81162 53830 81174 53882
rect 81236 53830 81238 53882
rect 81076 53828 81100 53830
rect 81156 53828 81180 53830
rect 81236 53828 81260 53830
rect 81020 53808 81316 53828
rect 81072 53508 81124 53514
rect 81072 53450 81124 53456
rect 81084 53106 81112 53450
rect 81072 53100 81124 53106
rect 81072 53042 81124 53048
rect 81020 52796 81316 52816
rect 81076 52794 81100 52796
rect 81156 52794 81180 52796
rect 81236 52794 81260 52796
rect 81098 52742 81100 52794
rect 81162 52742 81174 52794
rect 81236 52742 81238 52794
rect 81076 52740 81100 52742
rect 81156 52740 81180 52742
rect 81236 52740 81260 52742
rect 81020 52720 81316 52740
rect 80888 52556 80940 52562
rect 80888 52498 80940 52504
rect 80980 52488 81032 52494
rect 80980 52430 81032 52436
rect 80992 51882 81020 52430
rect 80980 51876 81032 51882
rect 80980 51818 81032 51824
rect 81020 51708 81316 51728
rect 81076 51706 81100 51708
rect 81156 51706 81180 51708
rect 81236 51706 81260 51708
rect 81098 51654 81100 51706
rect 81162 51654 81174 51706
rect 81236 51654 81238 51706
rect 81076 51652 81100 51654
rect 81156 51652 81180 51654
rect 81236 51652 81260 51654
rect 81020 51632 81316 51652
rect 81020 50620 81316 50640
rect 81076 50618 81100 50620
rect 81156 50618 81180 50620
rect 81236 50618 81260 50620
rect 81098 50566 81100 50618
rect 81162 50566 81174 50618
rect 81236 50566 81238 50618
rect 81076 50564 81100 50566
rect 81156 50564 81180 50566
rect 81236 50564 81260 50566
rect 81020 50544 81316 50564
rect 81020 49532 81316 49552
rect 81076 49530 81100 49532
rect 81156 49530 81180 49532
rect 81236 49530 81260 49532
rect 81098 49478 81100 49530
rect 81162 49478 81174 49530
rect 81236 49478 81238 49530
rect 81076 49476 81100 49478
rect 81156 49476 81180 49478
rect 81236 49476 81260 49478
rect 81020 49456 81316 49476
rect 81020 48444 81316 48464
rect 81076 48442 81100 48444
rect 81156 48442 81180 48444
rect 81236 48442 81260 48444
rect 81098 48390 81100 48442
rect 81162 48390 81174 48442
rect 81236 48390 81238 48442
rect 81076 48388 81100 48390
rect 81156 48388 81180 48390
rect 81236 48388 81260 48390
rect 81020 48368 81316 48388
rect 81020 47356 81316 47376
rect 81076 47354 81100 47356
rect 81156 47354 81180 47356
rect 81236 47354 81260 47356
rect 81098 47302 81100 47354
rect 81162 47302 81174 47354
rect 81236 47302 81238 47354
rect 81076 47300 81100 47302
rect 81156 47300 81180 47302
rect 81236 47300 81260 47302
rect 81020 47280 81316 47300
rect 81020 46268 81316 46288
rect 81076 46266 81100 46268
rect 81156 46266 81180 46268
rect 81236 46266 81260 46268
rect 81098 46214 81100 46266
rect 81162 46214 81174 46266
rect 81236 46214 81238 46266
rect 81076 46212 81100 46214
rect 81156 46212 81180 46214
rect 81236 46212 81260 46214
rect 81020 46192 81316 46212
rect 81020 45180 81316 45200
rect 81076 45178 81100 45180
rect 81156 45178 81180 45180
rect 81236 45178 81260 45180
rect 81098 45126 81100 45178
rect 81162 45126 81174 45178
rect 81236 45126 81238 45178
rect 81076 45124 81100 45126
rect 81156 45124 81180 45126
rect 81236 45124 81260 45126
rect 81020 45104 81316 45124
rect 81020 44092 81316 44112
rect 81076 44090 81100 44092
rect 81156 44090 81180 44092
rect 81236 44090 81260 44092
rect 81098 44038 81100 44090
rect 81162 44038 81174 44090
rect 81236 44038 81238 44090
rect 81076 44036 81100 44038
rect 81156 44036 81180 44038
rect 81236 44036 81260 44038
rect 81020 44016 81316 44036
rect 81020 43004 81316 43024
rect 81076 43002 81100 43004
rect 81156 43002 81180 43004
rect 81236 43002 81260 43004
rect 81098 42950 81100 43002
rect 81162 42950 81174 43002
rect 81236 42950 81238 43002
rect 81076 42948 81100 42950
rect 81156 42948 81180 42950
rect 81236 42948 81260 42950
rect 81020 42928 81316 42948
rect 80888 42832 80940 42838
rect 80888 42774 80940 42780
rect 80796 24744 80848 24750
rect 80796 24686 80848 24692
rect 80612 21480 80664 21486
rect 80612 21422 80664 21428
rect 80796 21480 80848 21486
rect 80796 21422 80848 21428
rect 80704 12096 80756 12102
rect 80704 12038 80756 12044
rect 80716 11830 80744 12038
rect 80520 11824 80572 11830
rect 80520 11766 80572 11772
rect 80704 11824 80756 11830
rect 80704 11766 80756 11772
rect 80808 11286 80836 21422
rect 80900 11762 80928 42774
rect 81020 41916 81316 41936
rect 81076 41914 81100 41916
rect 81156 41914 81180 41916
rect 81236 41914 81260 41916
rect 81098 41862 81100 41914
rect 81162 41862 81174 41914
rect 81236 41862 81238 41914
rect 81076 41860 81100 41862
rect 81156 41860 81180 41862
rect 81236 41860 81260 41862
rect 81020 41840 81316 41860
rect 81020 40828 81316 40848
rect 81076 40826 81100 40828
rect 81156 40826 81180 40828
rect 81236 40826 81260 40828
rect 81098 40774 81100 40826
rect 81162 40774 81174 40826
rect 81236 40774 81238 40826
rect 81076 40772 81100 40774
rect 81156 40772 81180 40774
rect 81236 40772 81260 40774
rect 81020 40752 81316 40772
rect 81020 39740 81316 39760
rect 81076 39738 81100 39740
rect 81156 39738 81180 39740
rect 81236 39738 81260 39740
rect 81098 39686 81100 39738
rect 81162 39686 81174 39738
rect 81236 39686 81238 39738
rect 81076 39684 81100 39686
rect 81156 39684 81180 39686
rect 81236 39684 81260 39686
rect 81020 39664 81316 39684
rect 81020 38652 81316 38672
rect 81076 38650 81100 38652
rect 81156 38650 81180 38652
rect 81236 38650 81260 38652
rect 81098 38598 81100 38650
rect 81162 38598 81174 38650
rect 81236 38598 81238 38650
rect 81076 38596 81100 38598
rect 81156 38596 81180 38598
rect 81236 38596 81260 38598
rect 81020 38576 81316 38596
rect 81164 38208 81216 38214
rect 81164 38150 81216 38156
rect 81176 38010 81204 38150
rect 81164 38004 81216 38010
rect 81164 37946 81216 37952
rect 81176 37874 81204 37946
rect 81164 37868 81216 37874
rect 81164 37810 81216 37816
rect 81020 37564 81316 37584
rect 81076 37562 81100 37564
rect 81156 37562 81180 37564
rect 81236 37562 81260 37564
rect 81098 37510 81100 37562
rect 81162 37510 81174 37562
rect 81236 37510 81238 37562
rect 81076 37508 81100 37510
rect 81156 37508 81180 37510
rect 81236 37508 81260 37510
rect 81020 37488 81316 37508
rect 81020 36476 81316 36496
rect 81076 36474 81100 36476
rect 81156 36474 81180 36476
rect 81236 36474 81260 36476
rect 81098 36422 81100 36474
rect 81162 36422 81174 36474
rect 81236 36422 81238 36474
rect 81076 36420 81100 36422
rect 81156 36420 81180 36422
rect 81236 36420 81260 36422
rect 81020 36400 81316 36420
rect 81020 35388 81316 35408
rect 81076 35386 81100 35388
rect 81156 35386 81180 35388
rect 81236 35386 81260 35388
rect 81098 35334 81100 35386
rect 81162 35334 81174 35386
rect 81236 35334 81238 35386
rect 81076 35332 81100 35334
rect 81156 35332 81180 35334
rect 81236 35332 81260 35334
rect 81020 35312 81316 35332
rect 81020 34300 81316 34320
rect 81076 34298 81100 34300
rect 81156 34298 81180 34300
rect 81236 34298 81260 34300
rect 81098 34246 81100 34298
rect 81162 34246 81174 34298
rect 81236 34246 81238 34298
rect 81076 34244 81100 34246
rect 81156 34244 81180 34246
rect 81236 34244 81260 34246
rect 81020 34224 81316 34244
rect 81020 33212 81316 33232
rect 81076 33210 81100 33212
rect 81156 33210 81180 33212
rect 81236 33210 81260 33212
rect 81098 33158 81100 33210
rect 81162 33158 81174 33210
rect 81236 33158 81238 33210
rect 81076 33156 81100 33158
rect 81156 33156 81180 33158
rect 81236 33156 81260 33158
rect 81020 33136 81316 33156
rect 81020 32124 81316 32144
rect 81076 32122 81100 32124
rect 81156 32122 81180 32124
rect 81236 32122 81260 32124
rect 81098 32070 81100 32122
rect 81162 32070 81174 32122
rect 81236 32070 81238 32122
rect 81076 32068 81100 32070
rect 81156 32068 81180 32070
rect 81236 32068 81260 32070
rect 81020 32048 81316 32068
rect 81020 31036 81316 31056
rect 81076 31034 81100 31036
rect 81156 31034 81180 31036
rect 81236 31034 81260 31036
rect 81098 30982 81100 31034
rect 81162 30982 81174 31034
rect 81236 30982 81238 31034
rect 81076 30980 81100 30982
rect 81156 30980 81180 30982
rect 81236 30980 81260 30982
rect 81020 30960 81316 30980
rect 81020 29948 81316 29968
rect 81076 29946 81100 29948
rect 81156 29946 81180 29948
rect 81236 29946 81260 29948
rect 81098 29894 81100 29946
rect 81162 29894 81174 29946
rect 81236 29894 81238 29946
rect 81076 29892 81100 29894
rect 81156 29892 81180 29894
rect 81236 29892 81260 29894
rect 81020 29872 81316 29892
rect 81020 28860 81316 28880
rect 81076 28858 81100 28860
rect 81156 28858 81180 28860
rect 81236 28858 81260 28860
rect 81098 28806 81100 28858
rect 81162 28806 81174 28858
rect 81236 28806 81238 28858
rect 81076 28804 81100 28806
rect 81156 28804 81180 28806
rect 81236 28804 81260 28806
rect 81020 28784 81316 28804
rect 81020 27772 81316 27792
rect 81076 27770 81100 27772
rect 81156 27770 81180 27772
rect 81236 27770 81260 27772
rect 81098 27718 81100 27770
rect 81162 27718 81174 27770
rect 81236 27718 81238 27770
rect 81076 27716 81100 27718
rect 81156 27716 81180 27718
rect 81236 27716 81260 27718
rect 81020 27696 81316 27716
rect 81020 26684 81316 26704
rect 81076 26682 81100 26684
rect 81156 26682 81180 26684
rect 81236 26682 81260 26684
rect 81098 26630 81100 26682
rect 81162 26630 81174 26682
rect 81236 26630 81238 26682
rect 81076 26628 81100 26630
rect 81156 26628 81180 26630
rect 81236 26628 81260 26630
rect 81020 26608 81316 26628
rect 81020 25596 81316 25616
rect 81076 25594 81100 25596
rect 81156 25594 81180 25596
rect 81236 25594 81260 25596
rect 81098 25542 81100 25594
rect 81162 25542 81174 25594
rect 81236 25542 81238 25594
rect 81076 25540 81100 25542
rect 81156 25540 81180 25542
rect 81236 25540 81260 25542
rect 81020 25520 81316 25540
rect 80980 25152 81032 25158
rect 80980 25094 81032 25100
rect 80992 24886 81020 25094
rect 80980 24880 81032 24886
rect 80980 24822 81032 24828
rect 81020 24508 81316 24528
rect 81076 24506 81100 24508
rect 81156 24506 81180 24508
rect 81236 24506 81260 24508
rect 81098 24454 81100 24506
rect 81162 24454 81174 24506
rect 81236 24454 81238 24506
rect 81076 24452 81100 24454
rect 81156 24452 81180 24454
rect 81236 24452 81260 24454
rect 81020 24432 81316 24452
rect 81020 23420 81316 23440
rect 81076 23418 81100 23420
rect 81156 23418 81180 23420
rect 81236 23418 81260 23420
rect 81098 23366 81100 23418
rect 81162 23366 81174 23418
rect 81236 23366 81238 23418
rect 81076 23364 81100 23366
rect 81156 23364 81180 23366
rect 81236 23364 81260 23366
rect 81020 23344 81316 23364
rect 81020 22332 81316 22352
rect 81076 22330 81100 22332
rect 81156 22330 81180 22332
rect 81236 22330 81260 22332
rect 81098 22278 81100 22330
rect 81162 22278 81174 22330
rect 81236 22278 81238 22330
rect 81076 22276 81100 22278
rect 81156 22276 81180 22278
rect 81236 22276 81260 22278
rect 81020 22256 81316 22276
rect 81020 21244 81316 21264
rect 81076 21242 81100 21244
rect 81156 21242 81180 21244
rect 81236 21242 81260 21244
rect 81098 21190 81100 21242
rect 81162 21190 81174 21242
rect 81236 21190 81238 21242
rect 81076 21188 81100 21190
rect 81156 21188 81180 21190
rect 81236 21188 81260 21190
rect 81020 21168 81316 21188
rect 81020 20156 81316 20176
rect 81076 20154 81100 20156
rect 81156 20154 81180 20156
rect 81236 20154 81260 20156
rect 81098 20102 81100 20154
rect 81162 20102 81174 20154
rect 81236 20102 81238 20154
rect 81076 20100 81100 20102
rect 81156 20100 81180 20102
rect 81236 20100 81260 20102
rect 81020 20080 81316 20100
rect 81020 19068 81316 19088
rect 81076 19066 81100 19068
rect 81156 19066 81180 19068
rect 81236 19066 81260 19068
rect 81098 19014 81100 19066
rect 81162 19014 81174 19066
rect 81236 19014 81238 19066
rect 81076 19012 81100 19014
rect 81156 19012 81180 19014
rect 81236 19012 81260 19014
rect 81020 18992 81316 19012
rect 81020 17980 81316 18000
rect 81076 17978 81100 17980
rect 81156 17978 81180 17980
rect 81236 17978 81260 17980
rect 81098 17926 81100 17978
rect 81162 17926 81174 17978
rect 81236 17926 81238 17978
rect 81076 17924 81100 17926
rect 81156 17924 81180 17926
rect 81236 17924 81260 17926
rect 81020 17904 81316 17924
rect 81020 16892 81316 16912
rect 81076 16890 81100 16892
rect 81156 16890 81180 16892
rect 81236 16890 81260 16892
rect 81098 16838 81100 16890
rect 81162 16838 81174 16890
rect 81236 16838 81238 16890
rect 81076 16836 81100 16838
rect 81156 16836 81180 16838
rect 81236 16836 81260 16838
rect 81020 16816 81316 16836
rect 81020 15804 81316 15824
rect 81076 15802 81100 15804
rect 81156 15802 81180 15804
rect 81236 15802 81260 15804
rect 81098 15750 81100 15802
rect 81162 15750 81174 15802
rect 81236 15750 81238 15802
rect 81076 15748 81100 15750
rect 81156 15748 81180 15750
rect 81236 15748 81260 15750
rect 81020 15728 81316 15748
rect 81020 14716 81316 14736
rect 81076 14714 81100 14716
rect 81156 14714 81180 14716
rect 81236 14714 81260 14716
rect 81098 14662 81100 14714
rect 81162 14662 81174 14714
rect 81236 14662 81238 14714
rect 81076 14660 81100 14662
rect 81156 14660 81180 14662
rect 81236 14660 81260 14662
rect 81020 14640 81316 14660
rect 81020 13628 81316 13648
rect 81076 13626 81100 13628
rect 81156 13626 81180 13628
rect 81236 13626 81260 13628
rect 81098 13574 81100 13626
rect 81162 13574 81174 13626
rect 81236 13574 81238 13626
rect 81076 13572 81100 13574
rect 81156 13572 81180 13574
rect 81236 13572 81260 13574
rect 81020 13552 81316 13572
rect 81020 12540 81316 12560
rect 81076 12538 81100 12540
rect 81156 12538 81180 12540
rect 81236 12538 81260 12540
rect 81098 12486 81100 12538
rect 81162 12486 81174 12538
rect 81236 12486 81238 12538
rect 81076 12484 81100 12486
rect 81156 12484 81180 12486
rect 81236 12484 81260 12486
rect 81020 12464 81316 12484
rect 80888 11756 80940 11762
rect 80888 11698 80940 11704
rect 80888 11552 80940 11558
rect 80888 11494 80940 11500
rect 80796 11280 80848 11286
rect 80796 11222 80848 11228
rect 80900 10130 80928 11494
rect 81020 11452 81316 11472
rect 81076 11450 81100 11452
rect 81156 11450 81180 11452
rect 81236 11450 81260 11452
rect 81098 11398 81100 11450
rect 81162 11398 81174 11450
rect 81236 11398 81238 11450
rect 81076 11396 81100 11398
rect 81156 11396 81180 11398
rect 81236 11396 81260 11398
rect 81020 11376 81316 11396
rect 81020 10364 81316 10384
rect 81076 10362 81100 10364
rect 81156 10362 81180 10364
rect 81236 10362 81260 10364
rect 81098 10310 81100 10362
rect 81162 10310 81174 10362
rect 81236 10310 81238 10362
rect 81076 10308 81100 10310
rect 81156 10308 81180 10310
rect 81236 10308 81260 10310
rect 81020 10288 81316 10308
rect 80888 10124 80940 10130
rect 80888 10066 80940 10072
rect 81020 9276 81316 9296
rect 81076 9274 81100 9276
rect 81156 9274 81180 9276
rect 81236 9274 81260 9276
rect 81098 9222 81100 9274
rect 81162 9222 81174 9274
rect 81236 9222 81238 9274
rect 81076 9220 81100 9222
rect 81156 9220 81180 9222
rect 81236 9220 81260 9222
rect 81020 9200 81316 9220
rect 81020 8188 81316 8208
rect 81076 8186 81100 8188
rect 81156 8186 81180 8188
rect 81236 8186 81260 8188
rect 81098 8134 81100 8186
rect 81162 8134 81174 8186
rect 81236 8134 81238 8186
rect 81076 8132 81100 8134
rect 81156 8132 81180 8134
rect 81236 8132 81260 8134
rect 81020 8112 81316 8132
rect 81020 7100 81316 7120
rect 81076 7098 81100 7100
rect 81156 7098 81180 7100
rect 81236 7098 81260 7100
rect 81098 7046 81100 7098
rect 81162 7046 81174 7098
rect 81236 7046 81238 7098
rect 81076 7044 81100 7046
rect 81156 7044 81180 7046
rect 81236 7044 81260 7046
rect 81020 7024 81316 7044
rect 81020 6012 81316 6032
rect 81076 6010 81100 6012
rect 81156 6010 81180 6012
rect 81236 6010 81260 6012
rect 81098 5958 81100 6010
rect 81162 5958 81174 6010
rect 81236 5958 81238 6010
rect 81076 5956 81100 5958
rect 81156 5956 81180 5958
rect 81236 5956 81260 5958
rect 81020 5936 81316 5956
rect 80612 5296 80664 5302
rect 80612 5238 80664 5244
rect 80520 5160 80572 5166
rect 80520 5102 80572 5108
rect 80244 4072 80296 4078
rect 80244 4014 80296 4020
rect 80336 4072 80388 4078
rect 80336 4014 80388 4020
rect 80164 3590 80284 3618
rect 80152 3528 80204 3534
rect 80152 3470 80204 3476
rect 79980 2774 80100 2802
rect 79980 800 80008 2774
rect 80164 800 80192 3470
rect 80256 3194 80284 3590
rect 80244 3188 80296 3194
rect 80244 3130 80296 3136
rect 80256 2938 80284 3130
rect 80256 2922 80468 2938
rect 80256 2916 80480 2922
rect 80256 2910 80428 2916
rect 80428 2858 80480 2864
rect 80336 2848 80388 2854
rect 80336 2790 80388 2796
rect 80348 800 80376 2790
rect 80532 800 80560 5102
rect 80624 2582 80652 5238
rect 81020 4924 81316 4944
rect 81076 4922 81100 4924
rect 81156 4922 81180 4924
rect 81236 4922 81260 4924
rect 81098 4870 81100 4922
rect 81162 4870 81174 4922
rect 81236 4870 81238 4922
rect 81076 4868 81100 4870
rect 81156 4868 81180 4870
rect 81236 4868 81260 4870
rect 81020 4848 81316 4868
rect 80796 4684 80848 4690
rect 80796 4626 80848 4632
rect 80612 2576 80664 2582
rect 80612 2518 80664 2524
rect 80808 800 80836 4626
rect 81020 3836 81316 3856
rect 81076 3834 81100 3836
rect 81156 3834 81180 3836
rect 81236 3834 81260 3836
rect 81098 3782 81100 3834
rect 81162 3782 81174 3834
rect 81236 3782 81238 3834
rect 81076 3780 81100 3782
rect 81156 3780 81180 3782
rect 81236 3780 81260 3782
rect 81020 3760 81316 3780
rect 80888 3188 80940 3194
rect 80888 3130 80940 3136
rect 80900 1442 80928 3130
rect 81360 2990 81388 58278
rect 82004 49366 82032 66030
rect 81992 49360 82044 49366
rect 81992 49302 82044 49308
rect 81532 46912 81584 46918
rect 81532 46854 81584 46860
rect 81544 46442 81572 46854
rect 81532 46436 81584 46442
rect 81532 46378 81584 46384
rect 81544 31278 81572 46378
rect 81532 31272 81584 31278
rect 81532 31214 81584 31220
rect 81544 30394 81572 31214
rect 81532 30388 81584 30394
rect 81532 30330 81584 30336
rect 81532 17332 81584 17338
rect 81532 17274 81584 17280
rect 81544 17202 81572 17274
rect 81532 17196 81584 17202
rect 81532 17138 81584 17144
rect 81624 14612 81676 14618
rect 81624 14554 81676 14560
rect 81532 4820 81584 4826
rect 81532 4762 81584 4768
rect 81440 4684 81492 4690
rect 81440 4626 81492 4632
rect 81348 2984 81400 2990
rect 81348 2926 81400 2932
rect 81452 2802 81480 4626
rect 81544 3670 81572 4762
rect 81636 4146 81664 14554
rect 82096 4826 82124 85614
rect 82636 85060 82688 85066
rect 82636 85002 82688 85008
rect 82176 80096 82228 80102
rect 82176 80038 82228 80044
rect 82188 12238 82216 80038
rect 82268 77988 82320 77994
rect 82268 77930 82320 77936
rect 82280 49842 82308 77930
rect 82544 66088 82596 66094
rect 82544 66030 82596 66036
rect 82452 64048 82504 64054
rect 82452 63990 82504 63996
rect 82464 61334 82492 63990
rect 82452 61328 82504 61334
rect 82452 61270 82504 61276
rect 82360 57248 82412 57254
rect 82360 57190 82412 57196
rect 82268 49836 82320 49842
rect 82268 49778 82320 49784
rect 82268 45348 82320 45354
rect 82268 45290 82320 45296
rect 82176 12232 82228 12238
rect 82176 12174 82228 12180
rect 82280 5370 82308 45290
rect 82372 43450 82400 57190
rect 82452 45280 82504 45286
rect 82452 45222 82504 45228
rect 82360 43444 82412 43450
rect 82360 43386 82412 43392
rect 82360 30388 82412 30394
rect 82360 30330 82412 30336
rect 82268 5364 82320 5370
rect 82268 5306 82320 5312
rect 82084 4820 82136 4826
rect 82084 4762 82136 4768
rect 82372 4214 82400 30330
rect 82464 5914 82492 45222
rect 82556 43314 82584 66030
rect 82544 43308 82596 43314
rect 82544 43250 82596 43256
rect 82544 37664 82596 37670
rect 82544 37606 82596 37612
rect 82556 12714 82584 37606
rect 82648 19922 82676 85002
rect 82832 79354 82860 86022
rect 82820 79348 82872 79354
rect 82820 79290 82872 79296
rect 82728 78668 82780 78674
rect 82728 78610 82780 78616
rect 82740 78062 82768 78610
rect 82728 78056 82780 78062
rect 82728 77998 82780 78004
rect 82924 72554 82952 97106
rect 83016 96422 83044 97294
rect 83844 96558 83872 99200
rect 84672 97238 84700 99200
rect 84660 97232 84712 97238
rect 84660 97174 84712 97180
rect 85028 97164 85080 97170
rect 85028 97106 85080 97112
rect 85488 97164 85540 97170
rect 85488 97106 85540 97112
rect 84108 97096 84160 97102
rect 84108 97038 84160 97044
rect 84120 96626 84148 97038
rect 85040 96966 85068 97106
rect 85028 96960 85080 96966
rect 85028 96902 85080 96908
rect 84108 96620 84160 96626
rect 84108 96562 84160 96568
rect 83832 96552 83884 96558
rect 83832 96494 83884 96500
rect 83004 96416 83056 96422
rect 83004 96358 83056 96364
rect 83464 96076 83516 96082
rect 83464 96018 83516 96024
rect 83476 93770 83504 96018
rect 83832 96008 83884 96014
rect 83832 95950 83884 95956
rect 83844 94042 83872 95950
rect 83924 95940 83976 95946
rect 83924 95882 83976 95888
rect 83832 94036 83884 94042
rect 83832 93978 83884 93984
rect 83464 93764 83516 93770
rect 83464 93706 83516 93712
rect 83096 86216 83148 86222
rect 83096 86158 83148 86164
rect 83004 81932 83056 81938
rect 83004 81874 83056 81880
rect 83016 81258 83044 81874
rect 83004 81252 83056 81258
rect 83004 81194 83056 81200
rect 83108 79082 83136 86158
rect 83096 79076 83148 79082
rect 83096 79018 83148 79024
rect 83096 78056 83148 78062
rect 83096 77998 83148 78004
rect 83108 77722 83136 77998
rect 83096 77716 83148 77722
rect 83096 77658 83148 77664
rect 83476 74534 83504 93706
rect 83844 88262 83872 93978
rect 83832 88256 83884 88262
rect 83832 88198 83884 88204
rect 83648 81252 83700 81258
rect 83648 81194 83700 81200
rect 83476 74506 83596 74534
rect 82912 72548 82964 72554
rect 82912 72490 82964 72496
rect 83464 70848 83516 70854
rect 83464 70790 83516 70796
rect 83096 66088 83148 66094
rect 83096 66030 83148 66036
rect 83280 66088 83332 66094
rect 83280 66030 83332 66036
rect 82912 56296 82964 56302
rect 82912 56238 82964 56244
rect 82924 52494 82952 56238
rect 82912 52488 82964 52494
rect 82912 52430 82964 52436
rect 82728 49428 82780 49434
rect 82728 49370 82780 49376
rect 82636 19916 82688 19922
rect 82636 19858 82688 19864
rect 82544 12708 82596 12714
rect 82544 12650 82596 12656
rect 82452 5908 82504 5914
rect 82452 5850 82504 5856
rect 82360 4208 82412 4214
rect 82360 4150 82412 4156
rect 81624 4140 81676 4146
rect 81624 4082 81676 4088
rect 81992 4072 82044 4078
rect 81992 4014 82044 4020
rect 81808 4004 81860 4010
rect 81808 3946 81860 3952
rect 81532 3664 81584 3670
rect 81532 3606 81584 3612
rect 81624 3596 81676 3602
rect 81624 3538 81676 3544
rect 81360 2774 81480 2802
rect 81020 2748 81316 2768
rect 81076 2746 81100 2748
rect 81156 2746 81180 2748
rect 81236 2746 81260 2748
rect 81098 2694 81100 2746
rect 81162 2694 81174 2746
rect 81236 2694 81238 2746
rect 81076 2692 81100 2694
rect 81156 2692 81180 2694
rect 81236 2692 81260 2694
rect 81020 2672 81316 2692
rect 81360 2446 81388 2774
rect 81164 2440 81216 2446
rect 81164 2382 81216 2388
rect 81348 2440 81400 2446
rect 81348 2382 81400 2388
rect 80900 1414 81020 1442
rect 80992 800 81020 1414
rect 81176 800 81204 2382
rect 81636 2258 81664 3538
rect 81716 3392 81768 3398
rect 81716 3334 81768 3340
rect 81360 2230 81664 2258
rect 81360 800 81388 2230
rect 81728 1714 81756 3334
rect 81544 1686 81756 1714
rect 81544 800 81572 1686
rect 81820 800 81848 3946
rect 82004 800 82032 4014
rect 82360 3052 82412 3058
rect 82360 2994 82412 3000
rect 82176 2848 82228 2854
rect 82176 2790 82228 2796
rect 82188 800 82216 2790
rect 82372 800 82400 2994
rect 82636 2984 82688 2990
rect 82636 2926 82688 2932
rect 82648 1578 82676 2926
rect 82740 2650 82768 49370
rect 82924 14482 82952 52430
rect 83108 48006 83136 66030
rect 83188 60648 83240 60654
rect 83188 60590 83240 60596
rect 83096 48000 83148 48006
rect 83096 47942 83148 47948
rect 83200 28150 83228 60590
rect 83292 52426 83320 66030
rect 83476 64874 83504 70790
rect 83568 68882 83596 74506
rect 83556 68876 83608 68882
rect 83556 68818 83608 68824
rect 83556 65952 83608 65958
rect 83556 65894 83608 65900
rect 83568 65754 83596 65894
rect 83556 65748 83608 65754
rect 83556 65690 83608 65696
rect 83476 64846 83596 64874
rect 83464 62348 83516 62354
rect 83464 62290 83516 62296
rect 83476 61674 83504 62290
rect 83464 61668 83516 61674
rect 83464 61610 83516 61616
rect 83372 60648 83424 60654
rect 83372 60590 83424 60596
rect 83384 60178 83412 60590
rect 83372 60172 83424 60178
rect 83372 60114 83424 60120
rect 83280 52420 83332 52426
rect 83280 52362 83332 52368
rect 83292 51610 83320 52362
rect 83280 51604 83332 51610
rect 83280 51546 83332 51552
rect 83188 28144 83240 28150
rect 83188 28086 83240 28092
rect 83464 28008 83516 28014
rect 83464 27950 83516 27956
rect 82912 14476 82964 14482
rect 82912 14418 82964 14424
rect 82820 9444 82872 9450
rect 82820 9386 82872 9392
rect 82728 2644 82780 2650
rect 82728 2586 82780 2592
rect 82832 2582 82860 9386
rect 83476 9382 83504 27950
rect 83464 9376 83516 9382
rect 83464 9318 83516 9324
rect 82912 4684 82964 4690
rect 82912 4626 82964 4632
rect 82924 3058 82952 4626
rect 83568 4146 83596 64846
rect 83660 60734 83688 81194
rect 83740 61124 83792 61130
rect 83740 61066 83792 61072
rect 83752 60858 83780 61066
rect 83740 60852 83792 60858
rect 83740 60794 83792 60800
rect 83660 60706 83780 60734
rect 83648 60648 83700 60654
rect 83648 60590 83700 60596
rect 83660 60314 83688 60590
rect 83648 60308 83700 60314
rect 83648 60250 83700 60256
rect 83752 55894 83780 60706
rect 83936 58886 83964 95882
rect 84292 92064 84344 92070
rect 84292 92006 84344 92012
rect 84304 80918 84332 92006
rect 84568 87508 84620 87514
rect 84568 87450 84620 87456
rect 84580 86222 84608 87450
rect 84568 86216 84620 86222
rect 84568 86158 84620 86164
rect 84292 80912 84344 80918
rect 84292 80854 84344 80860
rect 84384 80776 84436 80782
rect 84384 80718 84436 80724
rect 84200 77988 84252 77994
rect 84200 77930 84252 77936
rect 84212 72826 84240 77930
rect 84200 72820 84252 72826
rect 84200 72762 84252 72768
rect 83924 58880 83976 58886
rect 83924 58822 83976 58828
rect 83740 55888 83792 55894
rect 83740 55830 83792 55836
rect 84108 55208 84160 55214
rect 84108 55150 84160 55156
rect 84120 54806 84148 55150
rect 84108 54800 84160 54806
rect 84108 54742 84160 54748
rect 83648 54732 83700 54738
rect 83648 54674 83700 54680
rect 83660 48210 83688 54674
rect 83740 51604 83792 51610
rect 83740 51546 83792 51552
rect 83648 48204 83700 48210
rect 83648 48146 83700 48152
rect 83648 37120 83700 37126
rect 83648 37062 83700 37068
rect 83660 19990 83688 37062
rect 83752 32298 83780 51546
rect 84200 49224 84252 49230
rect 84200 49166 84252 49172
rect 84212 48890 84240 49166
rect 84200 48884 84252 48890
rect 84200 48826 84252 48832
rect 84396 34950 84424 80718
rect 84476 80640 84528 80646
rect 84476 80582 84528 80588
rect 84384 34944 84436 34950
rect 84384 34886 84436 34892
rect 83740 32292 83792 32298
rect 83740 32234 83792 32240
rect 84108 29504 84160 29510
rect 84108 29446 84160 29452
rect 83648 19984 83700 19990
rect 83648 19926 83700 19932
rect 84120 5778 84148 29446
rect 84384 26308 84436 26314
rect 84384 26250 84436 26256
rect 84396 15162 84424 26250
rect 84384 15156 84436 15162
rect 84384 15098 84436 15104
rect 84488 12646 84516 80582
rect 84580 77994 84608 86158
rect 84660 80776 84712 80782
rect 84660 80718 84712 80724
rect 84568 77988 84620 77994
rect 84568 77930 84620 77936
rect 84568 72820 84620 72826
rect 84568 72762 84620 72768
rect 84580 70514 84608 72762
rect 84568 70508 84620 70514
rect 84568 70450 84620 70456
rect 84580 68814 84608 70450
rect 84568 68808 84620 68814
rect 84568 68750 84620 68756
rect 84580 65482 84608 68750
rect 84568 65476 84620 65482
rect 84568 65418 84620 65424
rect 84568 54528 84620 54534
rect 84568 54470 84620 54476
rect 84580 50182 84608 54470
rect 84568 50176 84620 50182
rect 84568 50118 84620 50124
rect 84568 30388 84620 30394
rect 84568 30330 84620 30336
rect 84476 12640 84528 12646
rect 84476 12582 84528 12588
rect 84108 5772 84160 5778
rect 84108 5714 84160 5720
rect 84580 5250 84608 30330
rect 84672 6730 84700 80718
rect 84752 80640 84804 80646
rect 84752 80582 84804 80588
rect 84764 7342 84792 80582
rect 84844 68808 84896 68814
rect 84844 68750 84896 68756
rect 84856 68134 84884 68750
rect 84844 68128 84896 68134
rect 84844 68070 84896 68076
rect 84936 61668 84988 61674
rect 84936 61610 84988 61616
rect 84844 60648 84896 60654
rect 84844 60590 84896 60596
rect 84856 60246 84884 60590
rect 84844 60240 84896 60246
rect 84844 60182 84896 60188
rect 84844 54528 84896 54534
rect 84844 54470 84896 54476
rect 84856 49978 84884 54470
rect 84844 49972 84896 49978
rect 84844 49914 84896 49920
rect 84844 46368 84896 46374
rect 84844 46310 84896 46316
rect 84856 30938 84884 46310
rect 84948 44198 84976 61610
rect 84936 44192 84988 44198
rect 84936 44134 84988 44140
rect 85040 32026 85068 96902
rect 85304 84040 85356 84046
rect 85304 83982 85356 83988
rect 85212 70440 85264 70446
rect 85212 70382 85264 70388
rect 85224 50794 85252 70382
rect 85212 50788 85264 50794
rect 85212 50730 85264 50736
rect 85028 32020 85080 32026
rect 85028 31962 85080 31968
rect 84844 30932 84896 30938
rect 84844 30874 84896 30880
rect 84856 30394 84884 30874
rect 84844 30388 84896 30394
rect 84844 30330 84896 30336
rect 84936 29776 84988 29782
rect 84936 29718 84988 29724
rect 84948 28490 84976 29718
rect 84936 28484 84988 28490
rect 84936 28426 84988 28432
rect 84844 27328 84896 27334
rect 84844 27270 84896 27276
rect 84856 27130 84884 27270
rect 84844 27124 84896 27130
rect 84844 27066 84896 27072
rect 84948 23746 84976 28426
rect 85212 24608 85264 24614
rect 85212 24550 85264 24556
rect 85224 23866 85252 24550
rect 85212 23860 85264 23866
rect 85212 23802 85264 23808
rect 84948 23718 85252 23746
rect 85120 22976 85172 22982
rect 85120 22918 85172 22924
rect 84752 7336 84804 7342
rect 84752 7278 84804 7284
rect 84660 6724 84712 6730
rect 84660 6666 84712 6672
rect 84936 5908 84988 5914
rect 84936 5850 84988 5856
rect 84580 5222 84700 5250
rect 84568 4820 84620 4826
rect 84568 4762 84620 4768
rect 83556 4140 83608 4146
rect 83556 4082 83608 4088
rect 83648 4072 83700 4078
rect 83648 4014 83700 4020
rect 84200 4072 84252 4078
rect 84200 4014 84252 4020
rect 83004 3596 83056 3602
rect 83004 3538 83056 3544
rect 82912 3052 82964 3058
rect 82912 2994 82964 3000
rect 82820 2576 82872 2582
rect 82820 2518 82872 2524
rect 82820 2304 82872 2310
rect 82820 2246 82872 2252
rect 82556 1550 82676 1578
rect 82556 800 82584 1550
rect 82832 800 82860 2246
rect 83016 800 83044 3538
rect 83280 2984 83332 2990
rect 83280 2926 83332 2932
rect 83292 1578 83320 2926
rect 83372 2304 83424 2310
rect 83372 2246 83424 2252
rect 83200 1550 83320 1578
rect 83200 800 83228 1550
rect 83384 800 83412 2246
rect 83660 800 83688 4014
rect 83924 2984 83976 2990
rect 83924 2926 83976 2932
rect 83936 1578 83964 2926
rect 84016 2372 84068 2378
rect 84016 2314 84068 2320
rect 83844 1550 83964 1578
rect 83844 800 83872 1550
rect 84028 800 84056 2314
rect 84212 800 84240 4014
rect 84476 3596 84528 3602
rect 84476 3538 84528 3544
rect 84488 3482 84516 3538
rect 84304 3454 84516 3482
rect 84304 3398 84332 3454
rect 84292 3392 84344 3398
rect 84292 3334 84344 3340
rect 84304 1358 84332 3334
rect 84384 2916 84436 2922
rect 84384 2858 84436 2864
rect 84292 1352 84344 1358
rect 84292 1294 84344 1300
rect 84396 800 84424 2858
rect 84580 2650 84608 4762
rect 84672 3602 84700 5222
rect 84752 4208 84804 4214
rect 84752 4150 84804 4156
rect 84764 3602 84792 4150
rect 84844 4072 84896 4078
rect 84844 4014 84896 4020
rect 84660 3596 84712 3602
rect 84660 3538 84712 3544
rect 84752 3596 84804 3602
rect 84752 3538 84804 3544
rect 84568 2644 84620 2650
rect 84568 2586 84620 2592
rect 84660 2440 84712 2446
rect 84660 2382 84712 2388
rect 84672 800 84700 2382
rect 84856 800 84884 4014
rect 84948 3602 84976 5850
rect 85028 5364 85080 5370
rect 85028 5306 85080 5312
rect 85040 3738 85068 5306
rect 85028 3732 85080 3738
rect 85028 3674 85080 3680
rect 84936 3596 84988 3602
rect 84936 3538 84988 3544
rect 85028 3596 85080 3602
rect 85028 3538 85080 3544
rect 85040 800 85068 3538
rect 85132 3126 85160 22918
rect 85224 5914 85252 23718
rect 85316 11830 85344 83982
rect 85396 65476 85448 65482
rect 85396 65418 85448 65424
rect 85408 64938 85436 65418
rect 85396 64932 85448 64938
rect 85396 64874 85448 64880
rect 85500 56166 85528 97106
rect 85592 96626 85620 99200
rect 85580 96620 85632 96626
rect 85580 96562 85632 96568
rect 86420 96558 86448 99200
rect 87340 97238 87368 99200
rect 88168 97322 88196 99200
rect 88168 97294 88288 97322
rect 87328 97232 87380 97238
rect 87328 97174 87380 97180
rect 87512 97164 87564 97170
rect 87512 97106 87564 97112
rect 88156 97164 88208 97170
rect 88156 97106 88208 97112
rect 87524 96966 87552 97106
rect 87512 96960 87564 96966
rect 87512 96902 87564 96908
rect 86408 96552 86460 96558
rect 86408 96494 86460 96500
rect 85856 93152 85908 93158
rect 85856 93094 85908 93100
rect 85764 84584 85816 84590
rect 85764 84526 85816 84532
rect 85672 84040 85724 84046
rect 85672 83982 85724 83988
rect 85684 71602 85712 83982
rect 85672 71596 85724 71602
rect 85672 71538 85724 71544
rect 85580 70304 85632 70310
rect 85580 70246 85632 70252
rect 85488 56160 85540 56166
rect 85488 56102 85540 56108
rect 85592 42838 85620 70246
rect 85672 55888 85724 55894
rect 85672 55830 85724 55836
rect 85580 42832 85632 42838
rect 85580 42774 85632 42780
rect 85580 24744 85632 24750
rect 85408 24692 85580 24698
rect 85408 24686 85632 24692
rect 85408 24670 85620 24686
rect 85408 24614 85436 24670
rect 85396 24608 85448 24614
rect 85396 24550 85448 24556
rect 85684 12306 85712 55830
rect 85776 53174 85804 84526
rect 85868 69018 85896 93094
rect 85948 84448 86000 84454
rect 85948 84390 86000 84396
rect 85856 69012 85908 69018
rect 85856 68954 85908 68960
rect 85960 60734 85988 84390
rect 86224 84108 86276 84114
rect 86224 84050 86276 84056
rect 86132 84040 86184 84046
rect 86132 83982 86184 83988
rect 86144 83502 86172 83982
rect 86236 83570 86264 84050
rect 86224 83564 86276 83570
rect 86224 83506 86276 83512
rect 86132 83496 86184 83502
rect 86132 83438 86184 83444
rect 86236 79218 86264 83506
rect 86224 79212 86276 79218
rect 86224 79154 86276 79160
rect 86592 67108 86644 67114
rect 86592 67050 86644 67056
rect 85960 60706 86264 60734
rect 86236 58682 86264 60706
rect 86224 58676 86276 58682
rect 86224 58618 86276 58624
rect 85948 57452 86000 57458
rect 85948 57394 86000 57400
rect 85960 54534 85988 57394
rect 85948 54528 86000 54534
rect 85948 54470 86000 54476
rect 85764 53168 85816 53174
rect 85764 53110 85816 53116
rect 85960 49230 85988 54470
rect 85948 49224 86000 49230
rect 85948 49166 86000 49172
rect 85960 45830 85988 49166
rect 85948 45824 86000 45830
rect 85948 45766 86000 45772
rect 86236 42770 86264 58618
rect 86500 44192 86552 44198
rect 86500 44134 86552 44140
rect 86224 42764 86276 42770
rect 86224 42706 86276 42712
rect 86408 40724 86460 40730
rect 86408 40666 86460 40672
rect 86224 30184 86276 30190
rect 86224 30126 86276 30132
rect 86236 24750 86264 30126
rect 86420 24750 86448 40666
rect 86224 24744 86276 24750
rect 86224 24686 86276 24692
rect 86408 24744 86460 24750
rect 86408 24686 86460 24692
rect 85856 19916 85908 19922
rect 85856 19858 85908 19864
rect 85868 12306 85896 19858
rect 85948 16176 86000 16182
rect 85948 16118 86000 16124
rect 85672 12300 85724 12306
rect 85672 12242 85724 12248
rect 85856 12300 85908 12306
rect 85856 12242 85908 12248
rect 85304 11824 85356 11830
rect 85304 11766 85356 11772
rect 85580 7336 85632 7342
rect 85580 7278 85632 7284
rect 85212 5908 85264 5914
rect 85212 5850 85264 5856
rect 85396 4004 85448 4010
rect 85396 3946 85448 3952
rect 85120 3120 85172 3126
rect 85120 3062 85172 3068
rect 85212 2304 85264 2310
rect 85212 2246 85264 2252
rect 85224 800 85252 2246
rect 85408 800 85436 3946
rect 85592 2582 85620 7278
rect 85672 3596 85724 3602
rect 85672 3538 85724 3544
rect 85580 2576 85632 2582
rect 85580 2518 85632 2524
rect 85684 800 85712 3538
rect 85960 2582 85988 16118
rect 86512 12306 86540 44134
rect 86604 42566 86632 67050
rect 86960 64932 87012 64938
rect 86960 64874 87012 64880
rect 86972 60734 87000 64874
rect 86880 60706 87000 60734
rect 86880 59022 86908 60706
rect 86868 59016 86920 59022
rect 86868 58958 86920 58964
rect 86880 57458 86908 58958
rect 86868 57452 86920 57458
rect 86868 57394 86920 57400
rect 87524 48822 87552 96902
rect 88168 89622 88196 97106
rect 88260 96490 88288 97294
rect 88340 97028 88392 97034
rect 88340 96970 88392 96976
rect 88248 96484 88300 96490
rect 88248 96426 88300 96432
rect 88352 96422 88380 96970
rect 89088 96558 89116 99200
rect 89916 97238 89944 99200
rect 90456 97640 90508 97646
rect 90456 97582 90508 97588
rect 90468 97306 90496 97582
rect 90456 97300 90508 97306
rect 90456 97242 90508 97248
rect 89904 97232 89956 97238
rect 89904 97174 89956 97180
rect 89720 97164 89772 97170
rect 89720 97106 89772 97112
rect 89732 96966 89760 97106
rect 90640 97028 90692 97034
rect 90640 96970 90692 96976
rect 89720 96960 89772 96966
rect 89720 96902 89772 96908
rect 89076 96552 89128 96558
rect 89076 96494 89128 96500
rect 88340 96416 88392 96422
rect 88340 96358 88392 96364
rect 88984 95668 89036 95674
rect 88984 95610 89036 95616
rect 87972 89616 88024 89622
rect 87972 89558 88024 89564
rect 88156 89616 88208 89622
rect 88156 89558 88208 89564
rect 87880 75268 87932 75274
rect 87880 75210 87932 75216
rect 87696 64456 87748 64462
rect 87696 64398 87748 64404
rect 87512 48816 87564 48822
rect 87512 48758 87564 48764
rect 86960 47796 87012 47802
rect 86960 47738 87012 47744
rect 86684 47660 86736 47666
rect 86684 47602 86736 47608
rect 86696 47530 86724 47602
rect 86972 47598 87000 47738
rect 86868 47592 86920 47598
rect 86868 47534 86920 47540
rect 86960 47592 87012 47598
rect 86960 47534 87012 47540
rect 87328 47592 87380 47598
rect 87328 47534 87380 47540
rect 87420 47592 87472 47598
rect 87420 47534 87472 47540
rect 86684 47524 86736 47530
rect 86684 47466 86736 47472
rect 86880 47462 86908 47534
rect 86868 47456 86920 47462
rect 86868 47398 86920 47404
rect 87340 47122 87368 47534
rect 87432 47190 87460 47534
rect 87604 47524 87656 47530
rect 87604 47466 87656 47472
rect 87420 47184 87472 47190
rect 87420 47126 87472 47132
rect 87328 47116 87380 47122
rect 87328 47058 87380 47064
rect 86592 42560 86644 42566
rect 86592 42502 86644 42508
rect 86868 42560 86920 42566
rect 86868 42502 86920 42508
rect 86880 41750 86908 42502
rect 86868 41744 86920 41750
rect 86868 41686 86920 41692
rect 86868 40996 86920 41002
rect 86868 40938 86920 40944
rect 86880 40730 86908 40938
rect 86868 40724 86920 40730
rect 86868 40666 86920 40672
rect 87616 38486 87644 47466
rect 87604 38480 87656 38486
rect 87604 38422 87656 38428
rect 87708 37874 87736 64398
rect 87788 46504 87840 46510
rect 87788 46446 87840 46452
rect 87800 46102 87828 46446
rect 87788 46096 87840 46102
rect 87788 46038 87840 46044
rect 87696 37868 87748 37874
rect 87696 37810 87748 37816
rect 87788 37868 87840 37874
rect 87788 37810 87840 37816
rect 87512 37732 87564 37738
rect 87512 37674 87564 37680
rect 87524 37466 87552 37674
rect 87512 37460 87564 37466
rect 87512 37402 87564 37408
rect 87512 29844 87564 29850
rect 87512 29786 87564 29792
rect 87052 26988 87104 26994
rect 87052 26930 87104 26936
rect 87064 26790 87092 26930
rect 87052 26784 87104 26790
rect 87052 26726 87104 26732
rect 87420 26784 87472 26790
rect 87420 26726 87472 26732
rect 87432 26586 87460 26726
rect 87420 26580 87472 26586
rect 87420 26522 87472 26528
rect 87524 22094 87552 29786
rect 87432 22066 87552 22094
rect 86868 19236 86920 19242
rect 86868 19178 86920 19184
rect 86880 17134 86908 19178
rect 87432 17134 87460 22066
rect 86868 17128 86920 17134
rect 86868 17070 86920 17076
rect 87420 17128 87472 17134
rect 87420 17070 87472 17076
rect 87800 14822 87828 37810
rect 87788 14816 87840 14822
rect 87788 14758 87840 14764
rect 86500 12300 86552 12306
rect 86500 12242 86552 12248
rect 86408 12232 86460 12238
rect 86408 12174 86460 12180
rect 86420 9586 86448 12174
rect 86408 9580 86460 9586
rect 86408 9522 86460 9528
rect 86960 5024 87012 5030
rect 86960 4966 87012 4972
rect 86684 4072 86736 4078
rect 86684 4014 86736 4020
rect 86040 3528 86092 3534
rect 86040 3470 86092 3476
rect 85948 2576 86000 2582
rect 85948 2518 86000 2524
rect 85856 2372 85908 2378
rect 85856 2314 85908 2320
rect 85868 800 85896 2314
rect 86052 800 86080 3470
rect 86224 2984 86276 2990
rect 86224 2926 86276 2932
rect 86236 800 86264 2926
rect 86408 2440 86460 2446
rect 86408 2382 86460 2388
rect 86420 800 86448 2382
rect 86696 800 86724 4014
rect 86868 2984 86920 2990
rect 86868 2926 86920 2932
rect 86880 800 86908 2926
rect 86972 2582 87000 4966
rect 87236 4072 87288 4078
rect 87236 4014 87288 4020
rect 87052 2848 87104 2854
rect 87052 2790 87104 2796
rect 86960 2576 87012 2582
rect 86960 2518 87012 2524
rect 87064 800 87092 2790
rect 87248 800 87276 4014
rect 87512 2984 87564 2990
rect 87512 2926 87564 2932
rect 87524 800 87552 2926
rect 87892 2582 87920 75210
rect 87984 47598 88012 89558
rect 88248 89480 88300 89486
rect 88248 89422 88300 89428
rect 88616 89480 88668 89486
rect 88616 89422 88668 89428
rect 87972 47592 88024 47598
rect 87972 47534 88024 47540
rect 88156 47456 88208 47462
rect 88156 47398 88208 47404
rect 88168 47258 88196 47398
rect 88156 47252 88208 47258
rect 88156 47194 88208 47200
rect 88156 46572 88208 46578
rect 88156 46514 88208 46520
rect 87972 37460 88024 37466
rect 87972 37402 88024 37408
rect 87984 7206 88012 37402
rect 88064 29844 88116 29850
rect 88064 29786 88116 29792
rect 88076 29646 88104 29786
rect 88064 29640 88116 29646
rect 88064 29582 88116 29588
rect 88168 22030 88196 46514
rect 88156 22024 88208 22030
rect 88156 21966 88208 21972
rect 88260 13258 88288 89422
rect 88524 84040 88576 84046
rect 88524 83982 88576 83988
rect 88536 83706 88564 83982
rect 88524 83700 88576 83706
rect 88524 83642 88576 83648
rect 88340 65136 88392 65142
rect 88340 65078 88392 65084
rect 88248 13252 88300 13258
rect 88248 13194 88300 13200
rect 87972 7200 88024 7206
rect 87972 7142 88024 7148
rect 87972 3596 88024 3602
rect 87972 3538 88024 3544
rect 87880 2576 87932 2582
rect 87880 2518 87932 2524
rect 87788 2372 87840 2378
rect 87708 2332 87788 2360
rect 87708 800 87736 2332
rect 87788 2314 87840 2320
rect 87984 1306 88012 3538
rect 88156 2984 88208 2990
rect 87892 1278 88012 1306
rect 88076 2944 88156 2972
rect 87892 800 87920 1278
rect 88076 800 88104 2944
rect 88156 2926 88208 2932
rect 88352 2650 88380 65078
rect 88628 54738 88656 89422
rect 88708 69216 88760 69222
rect 88708 69158 88760 69164
rect 88616 54732 88668 54738
rect 88616 54674 88668 54680
rect 88432 40928 88484 40934
rect 88432 40870 88484 40876
rect 88444 36718 88472 40870
rect 88432 36712 88484 36718
rect 88432 36654 88484 36660
rect 88432 36576 88484 36582
rect 88432 36518 88484 36524
rect 88444 20466 88472 36518
rect 88432 20460 88484 20466
rect 88432 20402 88484 20408
rect 88524 4072 88576 4078
rect 88524 4014 88576 4020
rect 88340 2644 88392 2650
rect 88340 2586 88392 2592
rect 88248 2304 88300 2310
rect 88248 2246 88300 2252
rect 88260 800 88288 2246
rect 88536 800 88564 4014
rect 88720 3466 88748 69158
rect 88996 35894 89024 95610
rect 89628 87916 89680 87922
rect 89628 87858 89680 87864
rect 89640 87514 89668 87858
rect 89628 87508 89680 87514
rect 89628 87450 89680 87456
rect 89732 81734 89760 96902
rect 90652 96626 90680 96970
rect 90836 96626 90864 99200
rect 90640 96620 90692 96626
rect 90640 96562 90692 96568
rect 90824 96620 90876 96626
rect 90824 96562 90876 96568
rect 91664 96558 91692 99200
rect 92492 97238 92520 99200
rect 92480 97232 92532 97238
rect 92480 97174 92532 97180
rect 93308 97164 93360 97170
rect 93308 97106 93360 97112
rect 92756 97028 92808 97034
rect 92756 96970 92808 96976
rect 92296 96960 92348 96966
rect 92296 96902 92348 96908
rect 91652 96552 91704 96558
rect 91652 96494 91704 96500
rect 92204 92132 92256 92138
rect 92204 92074 92256 92080
rect 91744 90432 91796 90438
rect 91744 90374 91796 90380
rect 90272 88052 90324 88058
rect 90272 87994 90324 88000
rect 89812 87508 89864 87514
rect 89812 87450 89864 87456
rect 89824 87242 89852 87450
rect 90284 87378 90312 87994
rect 89904 87372 89956 87378
rect 89904 87314 89956 87320
rect 90272 87372 90324 87378
rect 90272 87314 90324 87320
rect 89812 87236 89864 87242
rect 89812 87178 89864 87184
rect 89916 81802 89944 87314
rect 90088 87304 90140 87310
rect 90088 87246 90140 87252
rect 89904 81796 89956 81802
rect 89904 81738 89956 81744
rect 89720 81728 89772 81734
rect 89720 81670 89772 81676
rect 89168 79756 89220 79762
rect 89168 79698 89220 79704
rect 89628 79756 89680 79762
rect 89628 79698 89680 79704
rect 89180 79558 89208 79698
rect 89352 79688 89404 79694
rect 89352 79630 89404 79636
rect 89364 79558 89392 79630
rect 89168 79552 89220 79558
rect 89168 79494 89220 79500
rect 89352 79552 89404 79558
rect 89352 79494 89404 79500
rect 89180 67318 89208 79494
rect 89260 71936 89312 71942
rect 89260 71878 89312 71884
rect 89272 69834 89300 71878
rect 89260 69828 89312 69834
rect 89260 69770 89312 69776
rect 89168 67312 89220 67318
rect 89168 67254 89220 67260
rect 89076 61056 89128 61062
rect 89076 60998 89128 61004
rect 88904 35866 89024 35894
rect 88904 31754 88932 35866
rect 88984 32224 89036 32230
rect 88984 32166 89036 32172
rect 88996 31890 89024 32166
rect 88984 31884 89036 31890
rect 88984 31826 89036 31832
rect 88904 31726 89024 31754
rect 88800 27668 88852 27674
rect 88800 27610 88852 27616
rect 88812 19990 88840 27610
rect 88800 19984 88852 19990
rect 88800 19926 88852 19932
rect 88996 5846 89024 31726
rect 89088 16114 89116 60998
rect 89260 36780 89312 36786
rect 89260 36722 89312 36728
rect 89272 29646 89300 36722
rect 89260 29640 89312 29646
rect 89260 29582 89312 29588
rect 89272 29306 89300 29582
rect 89260 29300 89312 29306
rect 89260 29242 89312 29248
rect 89076 16108 89128 16114
rect 89076 16050 89128 16056
rect 89364 11354 89392 79494
rect 89444 66836 89496 66842
rect 89444 66778 89496 66784
rect 89352 11348 89404 11354
rect 89352 11290 89404 11296
rect 88984 5840 89036 5846
rect 88984 5782 89036 5788
rect 89076 4072 89128 4078
rect 89076 4014 89128 4020
rect 88708 3460 88760 3466
rect 88708 3402 88760 3408
rect 88800 2984 88852 2990
rect 88720 2944 88800 2972
rect 88720 800 88748 2944
rect 88800 2926 88852 2932
rect 88892 2100 88944 2106
rect 88892 2042 88944 2048
rect 88904 800 88932 2042
rect 89088 800 89116 4014
rect 89260 3596 89312 3602
rect 89260 3538 89312 3544
rect 89272 800 89300 3538
rect 89456 2650 89484 66778
rect 89640 37738 89668 79698
rect 89812 79620 89864 79626
rect 89812 79562 89864 79568
rect 89824 38010 89852 79562
rect 90100 68406 90128 87246
rect 91008 87236 91060 87242
rect 91008 87178 91060 87184
rect 90548 86624 90600 86630
rect 90548 86566 90600 86572
rect 90272 86080 90324 86086
rect 90272 86022 90324 86028
rect 90180 68672 90232 68678
rect 90180 68614 90232 68620
rect 90088 68400 90140 68406
rect 90088 68342 90140 68348
rect 89904 60852 89956 60858
rect 89904 60794 89956 60800
rect 89916 60178 89944 60794
rect 89996 60716 90048 60722
rect 89996 60658 90048 60664
rect 89904 60172 89956 60178
rect 89904 60114 89956 60120
rect 90008 60110 90036 60658
rect 89996 60104 90048 60110
rect 89996 60046 90048 60052
rect 89812 38004 89864 38010
rect 89812 37946 89864 37952
rect 89628 37732 89680 37738
rect 89628 37674 89680 37680
rect 90192 27606 90220 68614
rect 90180 27600 90232 27606
rect 90180 27542 90232 27548
rect 89628 27532 89680 27538
rect 89628 27474 89680 27480
rect 89640 19718 89668 27474
rect 90180 23180 90232 23186
rect 90180 23122 90232 23128
rect 90192 21010 90220 23122
rect 90180 21004 90232 21010
rect 90180 20946 90232 20952
rect 90192 19854 90220 20946
rect 90180 19848 90232 19854
rect 90180 19790 90232 19796
rect 89628 19712 89680 19718
rect 89628 19654 89680 19660
rect 90284 12434 90312 86022
rect 90364 78464 90416 78470
rect 90364 78406 90416 78412
rect 90192 12406 90312 12434
rect 89720 4684 89772 4690
rect 89720 4626 89772 4632
rect 89628 2848 89680 2854
rect 89628 2790 89680 2796
rect 89444 2644 89496 2650
rect 89444 2586 89496 2592
rect 89640 2582 89668 2790
rect 89628 2576 89680 2582
rect 89628 2518 89680 2524
rect 89536 1216 89588 1222
rect 89536 1158 89588 1164
rect 89548 800 89576 1158
rect 89732 800 89760 4626
rect 90192 3942 90220 12406
rect 90272 4072 90324 4078
rect 90272 4014 90324 4020
rect 90180 3936 90232 3942
rect 90180 3878 90232 3884
rect 89904 3596 89956 3602
rect 89904 3538 89956 3544
rect 89916 800 89944 3538
rect 90088 2916 90140 2922
rect 90088 2858 90140 2864
rect 90100 800 90128 2858
rect 90284 800 90312 4014
rect 90376 2854 90404 78406
rect 90560 65210 90588 86566
rect 90916 67652 90968 67658
rect 90916 67594 90968 67600
rect 90548 65204 90600 65210
rect 90548 65146 90600 65152
rect 90824 61736 90876 61742
rect 90824 61678 90876 61684
rect 90836 60858 90864 61678
rect 90824 60852 90876 60858
rect 90824 60794 90876 60800
rect 90456 50380 90508 50386
rect 90456 50322 90508 50328
rect 90468 45558 90496 50322
rect 90548 46028 90600 46034
rect 90548 45970 90600 45976
rect 90456 45552 90508 45558
rect 90456 45494 90508 45500
rect 90468 23066 90496 45494
rect 90560 40730 90588 45970
rect 90548 40724 90600 40730
rect 90548 40666 90600 40672
rect 90732 34128 90784 34134
rect 90732 34070 90784 34076
rect 90640 29300 90692 29306
rect 90640 29242 90692 29248
rect 90468 23038 90588 23066
rect 90560 19922 90588 23038
rect 90548 19916 90600 19922
rect 90548 19858 90600 19864
rect 90456 19848 90508 19854
rect 90456 19790 90508 19796
rect 90468 6254 90496 19790
rect 90652 19174 90680 29242
rect 90640 19168 90692 19174
rect 90640 19110 90692 19116
rect 90456 6248 90508 6254
rect 90456 6190 90508 6196
rect 90468 5574 90496 6190
rect 90456 5568 90508 5574
rect 90456 5510 90508 5516
rect 90548 3596 90600 3602
rect 90548 3538 90600 3544
rect 90364 2848 90416 2854
rect 90364 2790 90416 2796
rect 90560 800 90588 3538
rect 90744 2650 90772 34070
rect 90824 33652 90876 33658
rect 90824 33594 90876 33600
rect 90836 3194 90864 33594
rect 90928 4162 90956 67594
rect 91020 9722 91048 87178
rect 91756 82074 91784 90374
rect 91744 82068 91796 82074
rect 91744 82010 91796 82016
rect 91100 75200 91152 75206
rect 91100 75142 91152 75148
rect 91112 22094 91140 75142
rect 91192 68468 91244 68474
rect 91192 68410 91244 68416
rect 91204 66162 91232 68410
rect 91836 68400 91888 68406
rect 91836 68342 91888 68348
rect 91744 68264 91796 68270
rect 91744 68206 91796 68212
rect 91192 66156 91244 66162
rect 91192 66098 91244 66104
rect 91192 65204 91244 65210
rect 91192 65146 91244 65152
rect 91204 64938 91232 65146
rect 91192 64932 91244 64938
rect 91192 64874 91244 64880
rect 91756 64530 91784 68206
rect 91848 64530 91876 68342
rect 91940 68338 92152 68354
rect 91928 68332 92164 68338
rect 91980 68326 92112 68332
rect 91928 68274 91980 68280
rect 92112 68274 92164 68280
rect 91744 64524 91796 64530
rect 91744 64466 91796 64472
rect 91836 64524 91888 64530
rect 91836 64466 91888 64472
rect 91756 55214 91784 64466
rect 91744 55208 91796 55214
rect 91744 55150 91796 55156
rect 91744 48272 91796 48278
rect 91744 48214 91796 48220
rect 91756 47802 91784 48214
rect 91744 47796 91796 47802
rect 91744 47738 91796 47744
rect 91756 47598 91784 47738
rect 91744 47592 91796 47598
rect 91744 47534 91796 47540
rect 91848 38282 91876 64466
rect 91928 61260 91980 61266
rect 91928 61202 91980 61208
rect 91940 60654 91968 61202
rect 92020 61124 92072 61130
rect 92020 61066 92072 61072
rect 91928 60648 91980 60654
rect 91928 60590 91980 60596
rect 91928 55208 91980 55214
rect 91928 55150 91980 55156
rect 91940 42634 91968 55150
rect 91928 42628 91980 42634
rect 91928 42570 91980 42576
rect 92032 40526 92060 61066
rect 92216 45554 92244 92074
rect 92124 45526 92244 45554
rect 92124 41002 92152 45526
rect 92112 40996 92164 41002
rect 92112 40938 92164 40944
rect 92020 40520 92072 40526
rect 92020 40462 92072 40468
rect 91836 38276 91888 38282
rect 91836 38218 91888 38224
rect 92032 31754 92060 40462
rect 92032 31726 92244 31754
rect 91928 28688 91980 28694
rect 91928 28630 91980 28636
rect 91652 28212 91704 28218
rect 91652 28154 91704 28160
rect 91112 22066 91232 22094
rect 91204 12434 91232 22066
rect 91204 12406 91416 12434
rect 91008 9716 91060 9722
rect 91008 9658 91060 9664
rect 91284 9376 91336 9382
rect 91284 9318 91336 9324
rect 90928 4134 91048 4162
rect 90916 4072 90968 4078
rect 90916 4014 90968 4020
rect 90824 3188 90876 3194
rect 90824 3130 90876 3136
rect 90836 2990 90864 3130
rect 90824 2984 90876 2990
rect 90824 2926 90876 2932
rect 90732 2644 90784 2650
rect 90732 2586 90784 2592
rect 90732 2304 90784 2310
rect 90732 2246 90784 2252
rect 90744 800 90772 2246
rect 90928 800 90956 4014
rect 91020 2922 91048 4134
rect 91100 3596 91152 3602
rect 91100 3538 91152 3544
rect 91008 2916 91060 2922
rect 91008 2858 91060 2864
rect 91008 2372 91060 2378
rect 91008 2314 91060 2320
rect 91020 2106 91048 2314
rect 91008 2100 91060 2106
rect 91008 2042 91060 2048
rect 91112 800 91140 3538
rect 91296 3194 91324 9318
rect 91284 3188 91336 3194
rect 91284 3130 91336 3136
rect 91284 2984 91336 2990
rect 91284 2926 91336 2932
rect 91296 800 91324 2926
rect 91388 2650 91416 12406
rect 91468 9172 91520 9178
rect 91468 9114 91520 9120
rect 91376 2644 91428 2650
rect 91376 2586 91428 2592
rect 91480 2582 91508 9114
rect 91664 5778 91692 28154
rect 91940 5778 91968 28630
rect 92112 14544 92164 14550
rect 92112 14486 92164 14492
rect 92124 6458 92152 14486
rect 92216 13802 92244 31726
rect 92308 15366 92336 96902
rect 92768 96490 92796 96970
rect 92756 96484 92808 96490
rect 92756 96426 92808 96432
rect 93216 96416 93268 96422
rect 93216 96358 93268 96364
rect 92664 92268 92716 92274
rect 92664 92210 92716 92216
rect 92480 92200 92532 92206
rect 92480 92142 92532 92148
rect 92492 69170 92520 92142
rect 92572 81864 92624 81870
rect 92572 81806 92624 81812
rect 92584 77994 92612 81806
rect 92572 77988 92624 77994
rect 92572 77930 92624 77936
rect 92584 76430 92612 77930
rect 92572 76424 92624 76430
rect 92572 76366 92624 76372
rect 92400 69142 92520 69170
rect 92400 69018 92428 69142
rect 92388 69012 92440 69018
rect 92388 68954 92440 68960
rect 92584 68898 92612 76366
rect 92400 68882 92612 68898
rect 92388 68876 92612 68882
rect 92440 68870 92612 68876
rect 92388 68818 92440 68824
rect 92676 56234 92704 92210
rect 93032 69896 93084 69902
rect 93032 69838 93084 69844
rect 92756 64388 92808 64394
rect 92756 64330 92808 64336
rect 92768 63850 92796 64330
rect 92756 63844 92808 63850
rect 92756 63786 92808 63792
rect 92940 63776 92992 63782
rect 92940 63718 92992 63724
rect 92664 56228 92716 56234
rect 92664 56170 92716 56176
rect 92848 49292 92900 49298
rect 92848 49234 92900 49240
rect 92480 48000 92532 48006
rect 92480 47942 92532 47948
rect 92492 47666 92520 47942
rect 92480 47660 92532 47666
rect 92480 47602 92532 47608
rect 92860 47598 92888 49234
rect 92848 47592 92900 47598
rect 92848 47534 92900 47540
rect 92860 42226 92888 47534
rect 92848 42220 92900 42226
rect 92848 42162 92900 42168
rect 92572 42152 92624 42158
rect 92572 42094 92624 42100
rect 92388 40520 92440 40526
rect 92388 40462 92440 40468
rect 92400 37942 92428 40462
rect 92388 37936 92440 37942
rect 92388 37878 92440 37884
rect 92388 32496 92440 32502
rect 92388 32438 92440 32444
rect 92400 30734 92428 32438
rect 92480 32428 92532 32434
rect 92480 32370 92532 32376
rect 92388 30728 92440 30734
rect 92388 30670 92440 30676
rect 92492 25702 92520 32370
rect 92480 25696 92532 25702
rect 92480 25638 92532 25644
rect 92296 15360 92348 15366
rect 92296 15302 92348 15308
rect 92204 13796 92256 13802
rect 92204 13738 92256 13744
rect 92216 13190 92244 13738
rect 92204 13184 92256 13190
rect 92204 13126 92256 13132
rect 92584 9654 92612 42094
rect 92664 37664 92716 37670
rect 92664 37606 92716 37612
rect 92676 31822 92704 37606
rect 92952 33998 92980 63718
rect 93044 37194 93072 69838
rect 93032 37188 93084 37194
rect 93032 37130 93084 37136
rect 92940 33992 92992 33998
rect 92940 33934 92992 33940
rect 92756 32224 92808 32230
rect 92756 32166 92808 32172
rect 92664 31816 92716 31822
rect 92664 31758 92716 31764
rect 92768 10062 92796 32166
rect 93228 10674 93256 96358
rect 93320 89714 93348 97106
rect 93412 96626 93440 99200
rect 93400 96620 93452 96626
rect 93400 96562 93452 96568
rect 94240 96558 94268 99200
rect 95160 97238 95188 99200
rect 95148 97232 95200 97238
rect 95148 97174 95200 97180
rect 95884 97028 95936 97034
rect 95884 96970 95936 96976
rect 94964 96960 95016 96966
rect 94964 96902 95016 96908
rect 94228 96552 94280 96558
rect 94228 96494 94280 96500
rect 93768 92336 93820 92342
rect 93768 92278 93820 92284
rect 93676 92200 93728 92206
rect 93676 92142 93728 92148
rect 93492 92132 93544 92138
rect 93492 92074 93544 92080
rect 93320 89686 93440 89714
rect 93412 70394 93440 89686
rect 93320 70366 93440 70394
rect 93320 55214 93348 70366
rect 93504 62830 93532 92074
rect 93584 76492 93636 76498
rect 93584 76434 93636 76440
rect 93596 76294 93624 76434
rect 93584 76288 93636 76294
rect 93584 76230 93636 76236
rect 93492 62824 93544 62830
rect 93492 62766 93544 62772
rect 93400 61600 93452 61606
rect 93400 61542 93452 61548
rect 93412 61402 93440 61542
rect 93400 61396 93452 61402
rect 93400 61338 93452 61344
rect 93320 55186 93440 55214
rect 93216 10668 93268 10674
rect 93216 10610 93268 10616
rect 93412 10130 93440 55186
rect 93596 10470 93624 76230
rect 93688 72010 93716 92142
rect 93780 77586 93808 92278
rect 93860 92268 93912 92274
rect 93860 92210 93912 92216
rect 93768 77580 93820 77586
rect 93768 77522 93820 77528
rect 93676 72004 93728 72010
rect 93676 71946 93728 71952
rect 93676 59220 93728 59226
rect 93676 59162 93728 59168
rect 93688 59022 93716 59162
rect 93676 59016 93728 59022
rect 93676 58958 93728 58964
rect 93676 57792 93728 57798
rect 93676 57734 93728 57740
rect 93584 10464 93636 10470
rect 93584 10406 93636 10412
rect 93400 10124 93452 10130
rect 93400 10066 93452 10072
rect 92756 10056 92808 10062
rect 92756 9998 92808 10004
rect 92572 9648 92624 9654
rect 92572 9590 92624 9596
rect 92848 9512 92900 9518
rect 92848 9454 92900 9460
rect 92112 6452 92164 6458
rect 92112 6394 92164 6400
rect 91652 5772 91704 5778
rect 91652 5714 91704 5720
rect 91928 5772 91980 5778
rect 91928 5714 91980 5720
rect 91560 4072 91612 4078
rect 91560 4014 91612 4020
rect 92112 4072 92164 4078
rect 92112 4014 92164 4020
rect 92756 4072 92808 4078
rect 92756 4014 92808 4020
rect 91468 2576 91520 2582
rect 91468 2518 91520 2524
rect 91572 800 91600 4014
rect 91744 2984 91796 2990
rect 91744 2926 91796 2932
rect 91756 800 91784 2926
rect 91928 2440 91980 2446
rect 91928 2382 91980 2388
rect 91940 800 91968 2382
rect 92124 800 92152 4014
rect 92388 3596 92440 3602
rect 92388 3538 92440 3544
rect 92400 800 92428 3538
rect 92572 1420 92624 1426
rect 92572 1362 92624 1368
rect 92584 800 92612 1362
rect 92768 800 92796 4014
rect 92860 2650 92888 9454
rect 93400 4684 93452 4690
rect 93400 4626 93452 4632
rect 92940 3596 92992 3602
rect 92940 3538 92992 3544
rect 92848 2644 92900 2650
rect 92848 2586 92900 2592
rect 92952 800 92980 3538
rect 93124 2916 93176 2922
rect 93124 2858 93176 2864
rect 93032 2372 93084 2378
rect 93032 2314 93084 2320
rect 93044 1222 93072 2314
rect 93032 1216 93084 1222
rect 93032 1158 93084 1164
rect 93136 800 93164 2858
rect 93412 800 93440 4626
rect 93584 3596 93636 3602
rect 93584 3538 93636 3544
rect 93596 800 93624 3538
rect 93688 3194 93716 57734
rect 93872 37806 93900 92210
rect 94136 92064 94188 92070
rect 94136 92006 94188 92012
rect 93952 75200 94004 75206
rect 93952 75142 94004 75148
rect 93860 37800 93912 37806
rect 93860 37742 93912 37748
rect 93860 15904 93912 15910
rect 93860 15846 93912 15852
rect 93872 7954 93900 15846
rect 93860 7948 93912 7954
rect 93860 7890 93912 7896
rect 93964 7562 93992 75142
rect 94044 56976 94096 56982
rect 94044 56918 94096 56924
rect 94056 55146 94084 56918
rect 94044 55140 94096 55146
rect 94044 55082 94096 55088
rect 94044 43308 94096 43314
rect 94044 43250 94096 43256
rect 94056 31958 94084 43250
rect 94044 31952 94096 31958
rect 94044 31894 94096 31900
rect 94044 13796 94096 13802
rect 94044 13738 94096 13744
rect 94056 9450 94084 13738
rect 94148 9994 94176 92006
rect 94504 75404 94556 75410
rect 94504 75346 94556 75352
rect 94320 57384 94372 57390
rect 94320 57326 94372 57332
rect 94228 38548 94280 38554
rect 94228 38490 94280 38496
rect 94240 37330 94268 38490
rect 94228 37324 94280 37330
rect 94228 37266 94280 37272
rect 94136 9988 94188 9994
rect 94136 9930 94188 9936
rect 94044 9444 94096 9450
rect 94044 9386 94096 9392
rect 93872 7534 93992 7562
rect 93676 3188 93728 3194
rect 93676 3130 93728 3136
rect 93688 2990 93716 3130
rect 93676 2984 93728 2990
rect 93676 2926 93728 2932
rect 93768 2916 93820 2922
rect 93768 2858 93820 2864
rect 93780 800 93808 2858
rect 93872 2582 93900 7534
rect 93952 4684 94004 4690
rect 93952 4626 94004 4632
rect 93860 2576 93912 2582
rect 93860 2518 93912 2524
rect 93964 800 93992 4626
rect 94136 4072 94188 4078
rect 94136 4014 94188 4020
rect 94148 800 94176 4014
rect 94332 2650 94360 57326
rect 94412 9444 94464 9450
rect 94412 9386 94464 9392
rect 94424 7954 94452 9386
rect 94412 7948 94464 7954
rect 94412 7890 94464 7896
rect 94412 7744 94464 7750
rect 94412 7686 94464 7692
rect 94424 7002 94452 7686
rect 94412 6996 94464 7002
rect 94412 6938 94464 6944
rect 94516 3534 94544 75346
rect 94780 70916 94832 70922
rect 94780 70858 94832 70864
rect 94792 22094 94820 70858
rect 94976 56710 95004 96902
rect 95896 96626 95924 96970
rect 95988 96626 96016 99200
rect 96380 96860 96676 96880
rect 96436 96858 96460 96860
rect 96516 96858 96540 96860
rect 96596 96858 96620 96860
rect 96458 96806 96460 96858
rect 96522 96806 96534 96858
rect 96596 96806 96598 96858
rect 96436 96804 96460 96806
rect 96516 96804 96540 96806
rect 96596 96804 96620 96806
rect 96380 96784 96676 96804
rect 95884 96620 95936 96626
rect 95884 96562 95936 96568
rect 95976 96620 96028 96626
rect 95976 96562 96028 96568
rect 96068 96484 96120 96490
rect 96068 96426 96120 96432
rect 95884 96416 95936 96422
rect 95884 96358 95936 96364
rect 95608 93968 95660 93974
rect 95608 93910 95660 93916
rect 95620 93702 95648 93910
rect 95608 93696 95660 93702
rect 95608 93638 95660 93644
rect 95700 85264 95752 85270
rect 95700 85206 95752 85212
rect 95240 81728 95292 81734
rect 95240 81670 95292 81676
rect 95252 81530 95280 81670
rect 95240 81524 95292 81530
rect 95240 81466 95292 81472
rect 95148 76288 95200 76294
rect 95148 76230 95200 76236
rect 95160 76090 95188 76230
rect 95148 76084 95200 76090
rect 95148 76026 95200 76032
rect 95608 70984 95660 70990
rect 95608 70926 95660 70932
rect 95056 64524 95108 64530
rect 95056 64466 95108 64472
rect 94964 56704 95016 56710
rect 94964 56646 95016 56652
rect 95068 55894 95096 64466
rect 95240 64456 95292 64462
rect 95240 64398 95292 64404
rect 95056 55888 95108 55894
rect 95056 55830 95108 55836
rect 95056 32360 95108 32366
rect 95056 32302 95108 32308
rect 95068 32026 95096 32302
rect 95056 32020 95108 32026
rect 95056 31962 95108 31968
rect 95252 27334 95280 64398
rect 95424 54868 95476 54874
rect 95424 54810 95476 54816
rect 95240 27328 95292 27334
rect 95240 27270 95292 27276
rect 95436 22094 95464 54810
rect 95516 41676 95568 41682
rect 95516 41618 95568 41624
rect 95528 40730 95556 41618
rect 95516 40724 95568 40730
rect 95516 40666 95568 40672
rect 95620 22094 95648 70926
rect 95712 42294 95740 85206
rect 95792 64524 95844 64530
rect 95792 64466 95844 64472
rect 95804 53038 95832 64466
rect 95792 53032 95844 53038
rect 95792 52974 95844 52980
rect 95700 42288 95752 42294
rect 95700 42230 95752 42236
rect 95792 33856 95844 33862
rect 95792 33798 95844 33804
rect 95804 22094 95832 33798
rect 95896 22982 95924 96358
rect 95976 93900 96028 93906
rect 95976 93842 96028 93848
rect 95988 28218 96016 93842
rect 96080 74254 96108 96426
rect 96908 96082 96936 99200
rect 97736 97238 97764 99200
rect 97724 97232 97776 97238
rect 97724 97174 97776 97180
rect 97540 96960 97592 96966
rect 97540 96902 97592 96908
rect 96896 96076 96948 96082
rect 96896 96018 96948 96024
rect 96380 95772 96676 95792
rect 96436 95770 96460 95772
rect 96516 95770 96540 95772
rect 96596 95770 96620 95772
rect 96458 95718 96460 95770
rect 96522 95718 96534 95770
rect 96596 95718 96598 95770
rect 96436 95716 96460 95718
rect 96516 95716 96540 95718
rect 96596 95716 96620 95718
rect 96380 95696 96676 95716
rect 96160 95328 96212 95334
rect 96160 95270 96212 95276
rect 96068 74248 96120 74254
rect 96068 74190 96120 74196
rect 96068 56908 96120 56914
rect 96068 56850 96120 56856
rect 95976 28212 96028 28218
rect 95976 28154 96028 28160
rect 95976 26308 96028 26314
rect 95976 26250 96028 26256
rect 95884 22976 95936 22982
rect 95884 22918 95936 22924
rect 94792 22066 94912 22094
rect 95436 22066 95556 22094
rect 95620 22066 95740 22094
rect 95804 22066 95924 22094
rect 94596 4684 94648 4690
rect 94596 4626 94648 4632
rect 94504 3528 94556 3534
rect 94504 3470 94556 3476
rect 94412 2984 94464 2990
rect 94412 2926 94464 2932
rect 94320 2644 94372 2650
rect 94320 2586 94372 2592
rect 94228 2372 94280 2378
rect 94228 2314 94280 2320
rect 94240 1426 94268 2314
rect 94228 1420 94280 1426
rect 94228 1362 94280 1368
rect 94424 800 94452 2926
rect 94608 800 94636 4626
rect 94780 4072 94832 4078
rect 94780 4014 94832 4020
rect 94792 800 94820 4014
rect 94884 3738 94912 22066
rect 95240 20800 95292 20806
rect 95240 20742 95292 20748
rect 95252 20058 95280 20742
rect 95240 20052 95292 20058
rect 95240 19994 95292 20000
rect 95240 19236 95292 19242
rect 95240 19178 95292 19184
rect 95252 12306 95280 19178
rect 95240 12300 95292 12306
rect 95240 12242 95292 12248
rect 95240 4684 95292 4690
rect 95240 4626 95292 4632
rect 94872 3732 94924 3738
rect 94872 3674 94924 3680
rect 94964 3460 95016 3466
rect 94964 3402 95016 3408
rect 94976 800 95004 3402
rect 95252 2774 95280 4626
rect 95424 3596 95476 3602
rect 95424 3538 95476 3544
rect 95160 2746 95280 2774
rect 95160 800 95188 2746
rect 95436 800 95464 3538
rect 95528 2650 95556 22066
rect 95608 2848 95660 2854
rect 95608 2790 95660 2796
rect 95516 2644 95568 2650
rect 95516 2586 95568 2592
rect 95620 800 95648 2790
rect 95712 2514 95740 22066
rect 95792 4684 95844 4690
rect 95792 4626 95844 4632
rect 95700 2508 95752 2514
rect 95700 2450 95752 2456
rect 95804 800 95832 4626
rect 95896 3194 95924 22066
rect 95988 16250 96016 26250
rect 95976 16244 96028 16250
rect 95976 16186 96028 16192
rect 96080 14890 96108 56850
rect 96172 41614 96200 95270
rect 96380 94684 96676 94704
rect 96436 94682 96460 94684
rect 96516 94682 96540 94684
rect 96596 94682 96620 94684
rect 96458 94630 96460 94682
rect 96522 94630 96534 94682
rect 96596 94630 96598 94682
rect 96436 94628 96460 94630
rect 96516 94628 96540 94630
rect 96596 94628 96620 94630
rect 96380 94608 96676 94628
rect 96380 93596 96676 93616
rect 96436 93594 96460 93596
rect 96516 93594 96540 93596
rect 96596 93594 96620 93596
rect 96458 93542 96460 93594
rect 96522 93542 96534 93594
rect 96596 93542 96598 93594
rect 96436 93540 96460 93542
rect 96516 93540 96540 93542
rect 96596 93540 96620 93542
rect 96380 93520 96676 93540
rect 96380 92508 96676 92528
rect 96436 92506 96460 92508
rect 96516 92506 96540 92508
rect 96596 92506 96620 92508
rect 96458 92454 96460 92506
rect 96522 92454 96534 92506
rect 96596 92454 96598 92506
rect 96436 92452 96460 92454
rect 96516 92452 96540 92454
rect 96596 92452 96620 92454
rect 96380 92432 96676 92452
rect 96380 91420 96676 91440
rect 96436 91418 96460 91420
rect 96516 91418 96540 91420
rect 96596 91418 96620 91420
rect 96458 91366 96460 91418
rect 96522 91366 96534 91418
rect 96596 91366 96598 91418
rect 96436 91364 96460 91366
rect 96516 91364 96540 91366
rect 96596 91364 96620 91366
rect 96380 91344 96676 91364
rect 96380 90332 96676 90352
rect 96436 90330 96460 90332
rect 96516 90330 96540 90332
rect 96596 90330 96620 90332
rect 96458 90278 96460 90330
rect 96522 90278 96534 90330
rect 96596 90278 96598 90330
rect 96436 90276 96460 90278
rect 96516 90276 96540 90278
rect 96596 90276 96620 90278
rect 96380 90256 96676 90276
rect 96380 89244 96676 89264
rect 96436 89242 96460 89244
rect 96516 89242 96540 89244
rect 96596 89242 96620 89244
rect 96458 89190 96460 89242
rect 96522 89190 96534 89242
rect 96596 89190 96598 89242
rect 96436 89188 96460 89190
rect 96516 89188 96540 89190
rect 96596 89188 96620 89190
rect 96380 89168 96676 89188
rect 96380 88156 96676 88176
rect 96436 88154 96460 88156
rect 96516 88154 96540 88156
rect 96596 88154 96620 88156
rect 96458 88102 96460 88154
rect 96522 88102 96534 88154
rect 96596 88102 96598 88154
rect 96436 88100 96460 88102
rect 96516 88100 96540 88102
rect 96596 88100 96620 88102
rect 96380 88080 96676 88100
rect 96380 87068 96676 87088
rect 96436 87066 96460 87068
rect 96516 87066 96540 87068
rect 96596 87066 96620 87068
rect 96458 87014 96460 87066
rect 96522 87014 96534 87066
rect 96596 87014 96598 87066
rect 96436 87012 96460 87014
rect 96516 87012 96540 87014
rect 96596 87012 96620 87014
rect 96380 86992 96676 87012
rect 96380 85980 96676 86000
rect 96436 85978 96460 85980
rect 96516 85978 96540 85980
rect 96596 85978 96620 85980
rect 96458 85926 96460 85978
rect 96522 85926 96534 85978
rect 96596 85926 96598 85978
rect 96436 85924 96460 85926
rect 96516 85924 96540 85926
rect 96596 85924 96620 85926
rect 96380 85904 96676 85924
rect 96380 84892 96676 84912
rect 96436 84890 96460 84892
rect 96516 84890 96540 84892
rect 96596 84890 96620 84892
rect 96458 84838 96460 84890
rect 96522 84838 96534 84890
rect 96596 84838 96598 84890
rect 96436 84836 96460 84838
rect 96516 84836 96540 84838
rect 96596 84836 96620 84838
rect 96380 84816 96676 84836
rect 96896 83904 96948 83910
rect 96896 83846 96948 83852
rect 96380 83804 96676 83824
rect 96436 83802 96460 83804
rect 96516 83802 96540 83804
rect 96596 83802 96620 83804
rect 96458 83750 96460 83802
rect 96522 83750 96534 83802
rect 96596 83750 96598 83802
rect 96436 83748 96460 83750
rect 96516 83748 96540 83750
rect 96596 83748 96620 83750
rect 96380 83728 96676 83748
rect 96380 82716 96676 82736
rect 96436 82714 96460 82716
rect 96516 82714 96540 82716
rect 96596 82714 96620 82716
rect 96458 82662 96460 82714
rect 96522 82662 96534 82714
rect 96596 82662 96598 82714
rect 96436 82660 96460 82662
rect 96516 82660 96540 82662
rect 96596 82660 96620 82662
rect 96380 82640 96676 82660
rect 96380 81628 96676 81648
rect 96436 81626 96460 81628
rect 96516 81626 96540 81628
rect 96596 81626 96620 81628
rect 96458 81574 96460 81626
rect 96522 81574 96534 81626
rect 96596 81574 96598 81626
rect 96436 81572 96460 81574
rect 96516 81572 96540 81574
rect 96596 81572 96620 81574
rect 96380 81552 96676 81572
rect 96380 80540 96676 80560
rect 96436 80538 96460 80540
rect 96516 80538 96540 80540
rect 96596 80538 96620 80540
rect 96458 80486 96460 80538
rect 96522 80486 96534 80538
rect 96596 80486 96598 80538
rect 96436 80484 96460 80486
rect 96516 80484 96540 80486
rect 96596 80484 96620 80486
rect 96380 80464 96676 80484
rect 96380 79452 96676 79472
rect 96436 79450 96460 79452
rect 96516 79450 96540 79452
rect 96596 79450 96620 79452
rect 96458 79398 96460 79450
rect 96522 79398 96534 79450
rect 96596 79398 96598 79450
rect 96436 79396 96460 79398
rect 96516 79396 96540 79398
rect 96596 79396 96620 79398
rect 96380 79376 96676 79396
rect 96908 79234 96936 83846
rect 97172 83428 97224 83434
rect 97172 83370 97224 83376
rect 96816 79206 96936 79234
rect 96380 78364 96676 78384
rect 96436 78362 96460 78364
rect 96516 78362 96540 78364
rect 96596 78362 96620 78364
rect 96458 78310 96460 78362
rect 96522 78310 96534 78362
rect 96596 78310 96598 78362
rect 96436 78308 96460 78310
rect 96516 78308 96540 78310
rect 96596 78308 96620 78310
rect 96380 78288 96676 78308
rect 96816 77654 96844 79206
rect 96896 79144 96948 79150
rect 96896 79086 96948 79092
rect 97080 79144 97132 79150
rect 97080 79086 97132 79092
rect 96804 77648 96856 77654
rect 96804 77590 96856 77596
rect 96380 77276 96676 77296
rect 96436 77274 96460 77276
rect 96516 77274 96540 77276
rect 96596 77274 96620 77276
rect 96458 77222 96460 77274
rect 96522 77222 96534 77274
rect 96596 77222 96598 77274
rect 96436 77220 96460 77222
rect 96516 77220 96540 77222
rect 96596 77220 96620 77222
rect 96380 77200 96676 77220
rect 96380 76188 96676 76208
rect 96436 76186 96460 76188
rect 96516 76186 96540 76188
rect 96596 76186 96620 76188
rect 96458 76134 96460 76186
rect 96522 76134 96534 76186
rect 96596 76134 96598 76186
rect 96436 76132 96460 76134
rect 96516 76132 96540 76134
rect 96596 76132 96620 76134
rect 96380 76112 96676 76132
rect 96380 75100 96676 75120
rect 96436 75098 96460 75100
rect 96516 75098 96540 75100
rect 96596 75098 96620 75100
rect 96458 75046 96460 75098
rect 96522 75046 96534 75098
rect 96596 75046 96598 75098
rect 96436 75044 96460 75046
rect 96516 75044 96540 75046
rect 96596 75044 96620 75046
rect 96380 75024 96676 75044
rect 96380 74012 96676 74032
rect 96436 74010 96460 74012
rect 96516 74010 96540 74012
rect 96596 74010 96620 74012
rect 96458 73958 96460 74010
rect 96522 73958 96534 74010
rect 96596 73958 96598 74010
rect 96436 73956 96460 73958
rect 96516 73956 96540 73958
rect 96596 73956 96620 73958
rect 96380 73936 96676 73956
rect 96380 72924 96676 72944
rect 96436 72922 96460 72924
rect 96516 72922 96540 72924
rect 96596 72922 96620 72924
rect 96458 72870 96460 72922
rect 96522 72870 96534 72922
rect 96596 72870 96598 72922
rect 96436 72868 96460 72870
rect 96516 72868 96540 72870
rect 96596 72868 96620 72870
rect 96380 72848 96676 72868
rect 96380 71836 96676 71856
rect 96436 71834 96460 71836
rect 96516 71834 96540 71836
rect 96596 71834 96620 71836
rect 96458 71782 96460 71834
rect 96522 71782 96534 71834
rect 96596 71782 96598 71834
rect 96436 71780 96460 71782
rect 96516 71780 96540 71782
rect 96596 71780 96620 71782
rect 96380 71760 96676 71780
rect 96380 70748 96676 70768
rect 96436 70746 96460 70748
rect 96516 70746 96540 70748
rect 96596 70746 96620 70748
rect 96458 70694 96460 70746
rect 96522 70694 96534 70746
rect 96596 70694 96598 70746
rect 96436 70692 96460 70694
rect 96516 70692 96540 70694
rect 96596 70692 96620 70694
rect 96380 70672 96676 70692
rect 96380 69660 96676 69680
rect 96436 69658 96460 69660
rect 96516 69658 96540 69660
rect 96596 69658 96620 69660
rect 96458 69606 96460 69658
rect 96522 69606 96534 69658
rect 96596 69606 96598 69658
rect 96436 69604 96460 69606
rect 96516 69604 96540 69606
rect 96596 69604 96620 69606
rect 96380 69584 96676 69604
rect 96380 68572 96676 68592
rect 96436 68570 96460 68572
rect 96516 68570 96540 68572
rect 96596 68570 96620 68572
rect 96458 68518 96460 68570
rect 96522 68518 96534 68570
rect 96596 68518 96598 68570
rect 96436 68516 96460 68518
rect 96516 68516 96540 68518
rect 96596 68516 96620 68518
rect 96380 68496 96676 68516
rect 96380 67484 96676 67504
rect 96436 67482 96460 67484
rect 96516 67482 96540 67484
rect 96596 67482 96620 67484
rect 96458 67430 96460 67482
rect 96522 67430 96534 67482
rect 96596 67430 96598 67482
rect 96436 67428 96460 67430
rect 96516 67428 96540 67430
rect 96596 67428 96620 67430
rect 96380 67408 96676 67428
rect 96380 66396 96676 66416
rect 96436 66394 96460 66396
rect 96516 66394 96540 66396
rect 96596 66394 96620 66396
rect 96458 66342 96460 66394
rect 96522 66342 96534 66394
rect 96596 66342 96598 66394
rect 96436 66340 96460 66342
rect 96516 66340 96540 66342
rect 96596 66340 96620 66342
rect 96380 66320 96676 66340
rect 96380 65308 96676 65328
rect 96436 65306 96460 65308
rect 96516 65306 96540 65308
rect 96596 65306 96620 65308
rect 96458 65254 96460 65306
rect 96522 65254 96534 65306
rect 96596 65254 96598 65306
rect 96436 65252 96460 65254
rect 96516 65252 96540 65254
rect 96596 65252 96620 65254
rect 96380 65232 96676 65252
rect 96380 64220 96676 64240
rect 96436 64218 96460 64220
rect 96516 64218 96540 64220
rect 96596 64218 96620 64220
rect 96458 64166 96460 64218
rect 96522 64166 96534 64218
rect 96596 64166 96598 64218
rect 96436 64164 96460 64166
rect 96516 64164 96540 64166
rect 96596 64164 96620 64166
rect 96380 64144 96676 64164
rect 96380 63132 96676 63152
rect 96436 63130 96460 63132
rect 96516 63130 96540 63132
rect 96596 63130 96620 63132
rect 96458 63078 96460 63130
rect 96522 63078 96534 63130
rect 96596 63078 96598 63130
rect 96436 63076 96460 63078
rect 96516 63076 96540 63078
rect 96596 63076 96620 63078
rect 96380 63056 96676 63076
rect 96380 62044 96676 62064
rect 96436 62042 96460 62044
rect 96516 62042 96540 62044
rect 96596 62042 96620 62044
rect 96458 61990 96460 62042
rect 96522 61990 96534 62042
rect 96596 61990 96598 62042
rect 96436 61988 96460 61990
rect 96516 61988 96540 61990
rect 96596 61988 96620 61990
rect 96380 61968 96676 61988
rect 96380 60956 96676 60976
rect 96436 60954 96460 60956
rect 96516 60954 96540 60956
rect 96596 60954 96620 60956
rect 96458 60902 96460 60954
rect 96522 60902 96534 60954
rect 96596 60902 96598 60954
rect 96436 60900 96460 60902
rect 96516 60900 96540 60902
rect 96596 60900 96620 60902
rect 96380 60880 96676 60900
rect 96380 59868 96676 59888
rect 96436 59866 96460 59868
rect 96516 59866 96540 59868
rect 96596 59866 96620 59868
rect 96458 59814 96460 59866
rect 96522 59814 96534 59866
rect 96596 59814 96598 59866
rect 96436 59812 96460 59814
rect 96516 59812 96540 59814
rect 96596 59812 96620 59814
rect 96380 59792 96676 59812
rect 96380 58780 96676 58800
rect 96436 58778 96460 58780
rect 96516 58778 96540 58780
rect 96596 58778 96620 58780
rect 96458 58726 96460 58778
rect 96522 58726 96534 58778
rect 96596 58726 96598 58778
rect 96436 58724 96460 58726
rect 96516 58724 96540 58726
rect 96596 58724 96620 58726
rect 96380 58704 96676 58724
rect 96380 57692 96676 57712
rect 96436 57690 96460 57692
rect 96516 57690 96540 57692
rect 96596 57690 96620 57692
rect 96458 57638 96460 57690
rect 96522 57638 96534 57690
rect 96596 57638 96598 57690
rect 96436 57636 96460 57638
rect 96516 57636 96540 57638
rect 96596 57636 96620 57638
rect 96380 57616 96676 57636
rect 96380 56604 96676 56624
rect 96436 56602 96460 56604
rect 96516 56602 96540 56604
rect 96596 56602 96620 56604
rect 96458 56550 96460 56602
rect 96522 56550 96534 56602
rect 96596 56550 96598 56602
rect 96436 56548 96460 56550
rect 96516 56548 96540 56550
rect 96596 56548 96620 56550
rect 96380 56528 96676 56548
rect 96252 56500 96304 56506
rect 96252 56442 96304 56448
rect 96160 41608 96212 41614
rect 96160 41550 96212 41556
rect 96160 29640 96212 29646
rect 96160 29582 96212 29588
rect 96172 18970 96200 29582
rect 96160 18964 96212 18970
rect 96160 18906 96212 18912
rect 96068 14884 96120 14890
rect 96068 14826 96120 14832
rect 96264 12434 96292 56442
rect 96380 55516 96676 55536
rect 96436 55514 96460 55516
rect 96516 55514 96540 55516
rect 96596 55514 96620 55516
rect 96458 55462 96460 55514
rect 96522 55462 96534 55514
rect 96596 55462 96598 55514
rect 96436 55460 96460 55462
rect 96516 55460 96540 55462
rect 96596 55460 96620 55462
rect 96380 55440 96676 55460
rect 96380 54428 96676 54448
rect 96436 54426 96460 54428
rect 96516 54426 96540 54428
rect 96596 54426 96620 54428
rect 96458 54374 96460 54426
rect 96522 54374 96534 54426
rect 96596 54374 96598 54426
rect 96436 54372 96460 54374
rect 96516 54372 96540 54374
rect 96596 54372 96620 54374
rect 96380 54352 96676 54372
rect 96380 53340 96676 53360
rect 96436 53338 96460 53340
rect 96516 53338 96540 53340
rect 96596 53338 96620 53340
rect 96458 53286 96460 53338
rect 96522 53286 96534 53338
rect 96596 53286 96598 53338
rect 96436 53284 96460 53286
rect 96516 53284 96540 53286
rect 96596 53284 96620 53286
rect 96380 53264 96676 53284
rect 96380 52252 96676 52272
rect 96436 52250 96460 52252
rect 96516 52250 96540 52252
rect 96596 52250 96620 52252
rect 96458 52198 96460 52250
rect 96522 52198 96534 52250
rect 96596 52198 96598 52250
rect 96436 52196 96460 52198
rect 96516 52196 96540 52198
rect 96596 52196 96620 52198
rect 96380 52176 96676 52196
rect 96380 51164 96676 51184
rect 96436 51162 96460 51164
rect 96516 51162 96540 51164
rect 96596 51162 96620 51164
rect 96458 51110 96460 51162
rect 96522 51110 96534 51162
rect 96596 51110 96598 51162
rect 96436 51108 96460 51110
rect 96516 51108 96540 51110
rect 96596 51108 96620 51110
rect 96380 51088 96676 51108
rect 96380 50076 96676 50096
rect 96436 50074 96460 50076
rect 96516 50074 96540 50076
rect 96596 50074 96620 50076
rect 96458 50022 96460 50074
rect 96522 50022 96534 50074
rect 96596 50022 96598 50074
rect 96436 50020 96460 50022
rect 96516 50020 96540 50022
rect 96596 50020 96620 50022
rect 96380 50000 96676 50020
rect 96380 48988 96676 49008
rect 96436 48986 96460 48988
rect 96516 48986 96540 48988
rect 96596 48986 96620 48988
rect 96458 48934 96460 48986
rect 96522 48934 96534 48986
rect 96596 48934 96598 48986
rect 96436 48932 96460 48934
rect 96516 48932 96540 48934
rect 96596 48932 96620 48934
rect 96380 48912 96676 48932
rect 96380 47900 96676 47920
rect 96436 47898 96460 47900
rect 96516 47898 96540 47900
rect 96596 47898 96620 47900
rect 96458 47846 96460 47898
rect 96522 47846 96534 47898
rect 96596 47846 96598 47898
rect 96436 47844 96460 47846
rect 96516 47844 96540 47846
rect 96596 47844 96620 47846
rect 96380 47824 96676 47844
rect 96380 46812 96676 46832
rect 96436 46810 96460 46812
rect 96516 46810 96540 46812
rect 96596 46810 96620 46812
rect 96458 46758 96460 46810
rect 96522 46758 96534 46810
rect 96596 46758 96598 46810
rect 96436 46756 96460 46758
rect 96516 46756 96540 46758
rect 96596 46756 96620 46758
rect 96380 46736 96676 46756
rect 96908 46646 96936 79086
rect 97092 74662 97120 79086
rect 97080 74656 97132 74662
rect 97080 74598 97132 74604
rect 97184 56914 97212 83370
rect 97448 79144 97500 79150
rect 97448 79086 97500 79092
rect 97172 56908 97224 56914
rect 97172 56850 97224 56856
rect 96896 46640 96948 46646
rect 96896 46582 96948 46588
rect 96380 45724 96676 45744
rect 96436 45722 96460 45724
rect 96516 45722 96540 45724
rect 96596 45722 96620 45724
rect 96458 45670 96460 45722
rect 96522 45670 96534 45722
rect 96596 45670 96598 45722
rect 96436 45668 96460 45670
rect 96516 45668 96540 45670
rect 96596 45668 96620 45670
rect 96380 45648 96676 45668
rect 96380 44636 96676 44656
rect 96436 44634 96460 44636
rect 96516 44634 96540 44636
rect 96596 44634 96620 44636
rect 96458 44582 96460 44634
rect 96522 44582 96534 44634
rect 96596 44582 96598 44634
rect 96436 44580 96460 44582
rect 96516 44580 96540 44582
rect 96596 44580 96620 44582
rect 96380 44560 96676 44580
rect 96380 43548 96676 43568
rect 96436 43546 96460 43548
rect 96516 43546 96540 43548
rect 96596 43546 96620 43548
rect 96458 43494 96460 43546
rect 96522 43494 96534 43546
rect 96596 43494 96598 43546
rect 96436 43492 96460 43494
rect 96516 43492 96540 43494
rect 96596 43492 96620 43494
rect 96380 43472 96676 43492
rect 96380 42460 96676 42480
rect 96436 42458 96460 42460
rect 96516 42458 96540 42460
rect 96596 42458 96620 42460
rect 96458 42406 96460 42458
rect 96522 42406 96534 42458
rect 96596 42406 96598 42458
rect 96436 42404 96460 42406
rect 96516 42404 96540 42406
rect 96596 42404 96620 42406
rect 96380 42384 96676 42404
rect 96528 42288 96580 42294
rect 96528 42230 96580 42236
rect 96540 41614 96568 42230
rect 96528 41608 96580 41614
rect 96528 41550 96580 41556
rect 96380 41372 96676 41392
rect 96436 41370 96460 41372
rect 96516 41370 96540 41372
rect 96596 41370 96620 41372
rect 96458 41318 96460 41370
rect 96522 41318 96534 41370
rect 96596 41318 96598 41370
rect 96436 41316 96460 41318
rect 96516 41316 96540 41318
rect 96596 41316 96620 41318
rect 96380 41296 96676 41316
rect 96380 40284 96676 40304
rect 96436 40282 96460 40284
rect 96516 40282 96540 40284
rect 96596 40282 96620 40284
rect 96458 40230 96460 40282
rect 96522 40230 96534 40282
rect 96596 40230 96598 40282
rect 96436 40228 96460 40230
rect 96516 40228 96540 40230
rect 96596 40228 96620 40230
rect 96380 40208 96676 40228
rect 96380 39196 96676 39216
rect 96436 39194 96460 39196
rect 96516 39194 96540 39196
rect 96596 39194 96620 39196
rect 96458 39142 96460 39194
rect 96522 39142 96534 39194
rect 96596 39142 96598 39194
rect 96436 39140 96460 39142
rect 96516 39140 96540 39142
rect 96596 39140 96620 39142
rect 96380 39120 96676 39140
rect 96380 38108 96676 38128
rect 96436 38106 96460 38108
rect 96516 38106 96540 38108
rect 96596 38106 96620 38108
rect 96458 38054 96460 38106
rect 96522 38054 96534 38106
rect 96596 38054 96598 38106
rect 96436 38052 96460 38054
rect 96516 38052 96540 38054
rect 96596 38052 96620 38054
rect 96380 38032 96676 38052
rect 96380 37020 96676 37040
rect 96436 37018 96460 37020
rect 96516 37018 96540 37020
rect 96596 37018 96620 37020
rect 96458 36966 96460 37018
rect 96522 36966 96534 37018
rect 96596 36966 96598 37018
rect 96436 36964 96460 36966
rect 96516 36964 96540 36966
rect 96596 36964 96620 36966
rect 96380 36944 96676 36964
rect 96380 35932 96676 35952
rect 96436 35930 96460 35932
rect 96516 35930 96540 35932
rect 96596 35930 96620 35932
rect 96458 35878 96460 35930
rect 96522 35878 96534 35930
rect 96596 35878 96598 35930
rect 96436 35876 96460 35878
rect 96516 35876 96540 35878
rect 96596 35876 96620 35878
rect 96380 35856 96676 35876
rect 96380 34844 96676 34864
rect 96436 34842 96460 34844
rect 96516 34842 96540 34844
rect 96596 34842 96620 34844
rect 96458 34790 96460 34842
rect 96522 34790 96534 34842
rect 96596 34790 96598 34842
rect 96436 34788 96460 34790
rect 96516 34788 96540 34790
rect 96596 34788 96620 34790
rect 96380 34768 96676 34788
rect 96380 33756 96676 33776
rect 96436 33754 96460 33756
rect 96516 33754 96540 33756
rect 96596 33754 96620 33756
rect 96458 33702 96460 33754
rect 96522 33702 96534 33754
rect 96596 33702 96598 33754
rect 96436 33700 96460 33702
rect 96516 33700 96540 33702
rect 96596 33700 96620 33702
rect 96380 33680 96676 33700
rect 96380 32668 96676 32688
rect 96436 32666 96460 32668
rect 96516 32666 96540 32668
rect 96596 32666 96620 32668
rect 96458 32614 96460 32666
rect 96522 32614 96534 32666
rect 96596 32614 96598 32666
rect 96436 32612 96460 32614
rect 96516 32612 96540 32614
rect 96596 32612 96620 32614
rect 96380 32592 96676 32612
rect 96380 31580 96676 31600
rect 96436 31578 96460 31580
rect 96516 31578 96540 31580
rect 96596 31578 96620 31580
rect 96458 31526 96460 31578
rect 96522 31526 96534 31578
rect 96596 31526 96598 31578
rect 96436 31524 96460 31526
rect 96516 31524 96540 31526
rect 96596 31524 96620 31526
rect 96380 31504 96676 31524
rect 96380 30492 96676 30512
rect 96436 30490 96460 30492
rect 96516 30490 96540 30492
rect 96596 30490 96620 30492
rect 96458 30438 96460 30490
rect 96522 30438 96534 30490
rect 96596 30438 96598 30490
rect 96436 30436 96460 30438
rect 96516 30436 96540 30438
rect 96596 30436 96620 30438
rect 96380 30416 96676 30436
rect 96380 29404 96676 29424
rect 96436 29402 96460 29404
rect 96516 29402 96540 29404
rect 96596 29402 96620 29404
rect 96458 29350 96460 29402
rect 96522 29350 96534 29402
rect 96596 29350 96598 29402
rect 96436 29348 96460 29350
rect 96516 29348 96540 29350
rect 96596 29348 96620 29350
rect 96380 29328 96676 29348
rect 96380 28316 96676 28336
rect 96436 28314 96460 28316
rect 96516 28314 96540 28316
rect 96596 28314 96620 28316
rect 96458 28262 96460 28314
rect 96522 28262 96534 28314
rect 96596 28262 96598 28314
rect 96436 28260 96460 28262
rect 96516 28260 96540 28262
rect 96596 28260 96620 28262
rect 96380 28240 96676 28260
rect 96380 27228 96676 27248
rect 96436 27226 96460 27228
rect 96516 27226 96540 27228
rect 96596 27226 96620 27228
rect 96458 27174 96460 27226
rect 96522 27174 96534 27226
rect 96596 27174 96598 27226
rect 96436 27172 96460 27174
rect 96516 27172 96540 27174
rect 96596 27172 96620 27174
rect 96380 27152 96676 27172
rect 96380 26140 96676 26160
rect 96436 26138 96460 26140
rect 96516 26138 96540 26140
rect 96596 26138 96620 26140
rect 96458 26086 96460 26138
rect 96522 26086 96534 26138
rect 96596 26086 96598 26138
rect 96436 26084 96460 26086
rect 96516 26084 96540 26086
rect 96596 26084 96620 26086
rect 96380 26064 96676 26084
rect 96380 25052 96676 25072
rect 96436 25050 96460 25052
rect 96516 25050 96540 25052
rect 96596 25050 96620 25052
rect 96458 24998 96460 25050
rect 96522 24998 96534 25050
rect 96596 24998 96598 25050
rect 96436 24996 96460 24998
rect 96516 24996 96540 24998
rect 96596 24996 96620 24998
rect 96380 24976 96676 24996
rect 96380 23964 96676 23984
rect 96436 23962 96460 23964
rect 96516 23962 96540 23964
rect 96596 23962 96620 23964
rect 96458 23910 96460 23962
rect 96522 23910 96534 23962
rect 96596 23910 96598 23962
rect 96436 23908 96460 23910
rect 96516 23908 96540 23910
rect 96596 23908 96620 23910
rect 96380 23888 96676 23908
rect 96380 22876 96676 22896
rect 96436 22874 96460 22876
rect 96516 22874 96540 22876
rect 96596 22874 96620 22876
rect 96458 22822 96460 22874
rect 96522 22822 96534 22874
rect 96596 22822 96598 22874
rect 96436 22820 96460 22822
rect 96516 22820 96540 22822
rect 96596 22820 96620 22822
rect 96380 22800 96676 22820
rect 96380 21788 96676 21808
rect 96436 21786 96460 21788
rect 96516 21786 96540 21788
rect 96596 21786 96620 21788
rect 96458 21734 96460 21786
rect 96522 21734 96534 21786
rect 96596 21734 96598 21786
rect 96436 21732 96460 21734
rect 96516 21732 96540 21734
rect 96596 21732 96620 21734
rect 96380 21712 96676 21732
rect 97184 21146 97212 56850
rect 97460 39438 97488 79086
rect 97448 39432 97500 39438
rect 97448 39374 97500 39380
rect 97552 33454 97580 96902
rect 98656 96626 98684 99200
rect 98644 96620 98696 96626
rect 98644 96562 98696 96568
rect 99484 96558 99512 99200
rect 99472 96552 99524 96558
rect 99472 96494 99524 96500
rect 97908 96484 97960 96490
rect 97908 96426 97960 96432
rect 97632 86080 97684 86086
rect 97632 86022 97684 86028
rect 97540 33448 97592 33454
rect 97540 33390 97592 33396
rect 97644 22094 97672 86022
rect 97644 22066 97764 22094
rect 97172 21140 97224 21146
rect 97172 21082 97224 21088
rect 96380 20700 96676 20720
rect 96436 20698 96460 20700
rect 96516 20698 96540 20700
rect 96596 20698 96620 20700
rect 96458 20646 96460 20698
rect 96522 20646 96534 20698
rect 96596 20646 96598 20698
rect 96436 20644 96460 20646
rect 96516 20644 96540 20646
rect 96596 20644 96620 20646
rect 96380 20624 96676 20644
rect 96380 19612 96676 19632
rect 96436 19610 96460 19612
rect 96516 19610 96540 19612
rect 96596 19610 96620 19612
rect 96458 19558 96460 19610
rect 96522 19558 96534 19610
rect 96596 19558 96598 19610
rect 96436 19556 96460 19558
rect 96516 19556 96540 19558
rect 96596 19556 96620 19558
rect 96380 19536 96676 19556
rect 97264 19168 97316 19174
rect 97264 19110 97316 19116
rect 97276 18834 97304 19110
rect 96988 18828 97040 18834
rect 96988 18770 97040 18776
rect 97264 18828 97316 18834
rect 97264 18770 97316 18776
rect 96380 18524 96676 18544
rect 96436 18522 96460 18524
rect 96516 18522 96540 18524
rect 96596 18522 96620 18524
rect 96458 18470 96460 18522
rect 96522 18470 96534 18522
rect 96596 18470 96598 18522
rect 96436 18468 96460 18470
rect 96516 18468 96540 18470
rect 96596 18468 96620 18470
rect 96380 18448 96676 18468
rect 97000 18154 97028 18770
rect 96712 18148 96764 18154
rect 96712 18090 96764 18096
rect 96988 18148 97040 18154
rect 96988 18090 97040 18096
rect 96380 17436 96676 17456
rect 96436 17434 96460 17436
rect 96516 17434 96540 17436
rect 96596 17434 96620 17436
rect 96458 17382 96460 17434
rect 96522 17382 96534 17434
rect 96596 17382 96598 17434
rect 96436 17380 96460 17382
rect 96516 17380 96540 17382
rect 96596 17380 96620 17382
rect 96380 17360 96676 17380
rect 96380 16348 96676 16368
rect 96436 16346 96460 16348
rect 96516 16346 96540 16348
rect 96596 16346 96620 16348
rect 96458 16294 96460 16346
rect 96522 16294 96534 16346
rect 96596 16294 96598 16346
rect 96436 16292 96460 16294
rect 96516 16292 96540 16294
rect 96596 16292 96620 16294
rect 96380 16272 96676 16292
rect 96380 15260 96676 15280
rect 96436 15258 96460 15260
rect 96516 15258 96540 15260
rect 96596 15258 96620 15260
rect 96458 15206 96460 15258
rect 96522 15206 96534 15258
rect 96596 15206 96598 15258
rect 96436 15204 96460 15206
rect 96516 15204 96540 15206
rect 96596 15204 96620 15206
rect 96380 15184 96676 15204
rect 96380 14172 96676 14192
rect 96436 14170 96460 14172
rect 96516 14170 96540 14172
rect 96596 14170 96620 14172
rect 96458 14118 96460 14170
rect 96522 14118 96534 14170
rect 96596 14118 96598 14170
rect 96436 14116 96460 14118
rect 96516 14116 96540 14118
rect 96596 14116 96620 14118
rect 96380 14096 96676 14116
rect 96380 13084 96676 13104
rect 96436 13082 96460 13084
rect 96516 13082 96540 13084
rect 96596 13082 96620 13084
rect 96458 13030 96460 13082
rect 96522 13030 96534 13082
rect 96596 13030 96598 13082
rect 96436 13028 96460 13030
rect 96516 13028 96540 13030
rect 96596 13028 96620 13030
rect 96380 13008 96676 13028
rect 96724 12782 96752 18090
rect 97172 17128 97224 17134
rect 97172 17070 97224 17076
rect 97184 16794 97212 17070
rect 97172 16788 97224 16794
rect 97172 16730 97224 16736
rect 96712 12776 96764 12782
rect 96712 12718 96764 12724
rect 96172 12406 96292 12434
rect 96068 8968 96120 8974
rect 96068 8910 96120 8916
rect 95976 4072 96028 4078
rect 95976 4014 96028 4020
rect 95884 3188 95936 3194
rect 95884 3130 95936 3136
rect 95988 800 96016 4014
rect 96080 2990 96108 8910
rect 96068 2984 96120 2990
rect 96068 2926 96120 2932
rect 96172 2650 96200 12406
rect 96804 12232 96856 12238
rect 96804 12174 96856 12180
rect 96988 12232 97040 12238
rect 96988 12174 97040 12180
rect 96380 11996 96676 12016
rect 96436 11994 96460 11996
rect 96516 11994 96540 11996
rect 96596 11994 96620 11996
rect 96458 11942 96460 11994
rect 96522 11942 96534 11994
rect 96596 11942 96598 11994
rect 96436 11940 96460 11942
rect 96516 11940 96540 11942
rect 96596 11940 96620 11942
rect 96380 11920 96676 11940
rect 96380 10908 96676 10928
rect 96436 10906 96460 10908
rect 96516 10906 96540 10908
rect 96596 10906 96620 10908
rect 96458 10854 96460 10906
rect 96522 10854 96534 10906
rect 96596 10854 96598 10906
rect 96436 10852 96460 10854
rect 96516 10852 96540 10854
rect 96596 10852 96620 10854
rect 96380 10832 96676 10852
rect 96380 9820 96676 9840
rect 96436 9818 96460 9820
rect 96516 9818 96540 9820
rect 96596 9818 96620 9820
rect 96458 9766 96460 9818
rect 96522 9766 96534 9818
rect 96596 9766 96598 9818
rect 96436 9764 96460 9766
rect 96516 9764 96540 9766
rect 96596 9764 96620 9766
rect 96380 9744 96676 9764
rect 96380 8732 96676 8752
rect 96436 8730 96460 8732
rect 96516 8730 96540 8732
rect 96596 8730 96620 8732
rect 96458 8678 96460 8730
rect 96522 8678 96534 8730
rect 96596 8678 96598 8730
rect 96436 8676 96460 8678
rect 96516 8676 96540 8678
rect 96596 8676 96620 8678
rect 96380 8656 96676 8676
rect 96816 8090 96844 12174
rect 97000 11558 97028 12174
rect 97540 12096 97592 12102
rect 97540 12038 97592 12044
rect 97552 11898 97580 12038
rect 97540 11892 97592 11898
rect 97540 11834 97592 11840
rect 96988 11552 97040 11558
rect 96988 11494 97040 11500
rect 97448 9104 97500 9110
rect 97448 9046 97500 9052
rect 96896 9036 96948 9042
rect 96896 8978 96948 8984
rect 96804 8084 96856 8090
rect 96804 8026 96856 8032
rect 96380 7644 96676 7664
rect 96436 7642 96460 7644
rect 96516 7642 96540 7644
rect 96596 7642 96620 7644
rect 96458 7590 96460 7642
rect 96522 7590 96534 7642
rect 96596 7590 96598 7642
rect 96436 7588 96460 7590
rect 96516 7588 96540 7590
rect 96596 7588 96620 7590
rect 96380 7568 96676 7588
rect 96380 6556 96676 6576
rect 96436 6554 96460 6556
rect 96516 6554 96540 6556
rect 96596 6554 96620 6556
rect 96458 6502 96460 6554
rect 96522 6502 96534 6554
rect 96596 6502 96598 6554
rect 96436 6500 96460 6502
rect 96516 6500 96540 6502
rect 96596 6500 96620 6502
rect 96380 6480 96676 6500
rect 96380 5468 96676 5488
rect 96436 5466 96460 5468
rect 96516 5466 96540 5468
rect 96596 5466 96620 5468
rect 96458 5414 96460 5466
rect 96522 5414 96534 5466
rect 96596 5414 96598 5466
rect 96436 5412 96460 5414
rect 96516 5412 96540 5414
rect 96596 5412 96620 5414
rect 96380 5392 96676 5412
rect 96252 5160 96304 5166
rect 96252 5102 96304 5108
rect 96264 3074 96292 5102
rect 96712 4684 96764 4690
rect 96712 4626 96764 4632
rect 96380 4380 96676 4400
rect 96436 4378 96460 4380
rect 96516 4378 96540 4380
rect 96596 4378 96620 4380
rect 96458 4326 96460 4378
rect 96522 4326 96534 4378
rect 96596 4326 96598 4378
rect 96436 4324 96460 4326
rect 96516 4324 96540 4326
rect 96596 4324 96620 4326
rect 96380 4304 96676 4324
rect 96380 3292 96676 3312
rect 96436 3290 96460 3292
rect 96516 3290 96540 3292
rect 96596 3290 96620 3292
rect 96458 3238 96460 3290
rect 96522 3238 96534 3290
rect 96596 3238 96598 3290
rect 96436 3236 96460 3238
rect 96516 3236 96540 3238
rect 96596 3236 96620 3238
rect 96380 3216 96676 3236
rect 96264 3046 96476 3074
rect 96252 2916 96304 2922
rect 96252 2858 96304 2864
rect 96160 2644 96212 2650
rect 96160 2586 96212 2592
rect 96264 2530 96292 2858
rect 96172 2502 96292 2530
rect 96172 1306 96200 2502
rect 96448 2394 96476 3046
rect 96264 2366 96476 2394
rect 96264 1442 96292 2366
rect 96380 2204 96676 2224
rect 96436 2202 96460 2204
rect 96516 2202 96540 2204
rect 96596 2202 96620 2204
rect 96458 2150 96460 2202
rect 96522 2150 96534 2202
rect 96596 2150 96598 2202
rect 96436 2148 96460 2150
rect 96516 2148 96540 2150
rect 96596 2148 96620 2150
rect 96380 2128 96676 2148
rect 96724 1442 96752 4626
rect 96908 4146 96936 8978
rect 96988 5772 97040 5778
rect 96988 5714 97040 5720
rect 96896 4140 96948 4146
rect 96896 4082 96948 4088
rect 96804 2984 96856 2990
rect 96804 2926 96856 2932
rect 96264 1414 96476 1442
rect 96172 1278 96292 1306
rect 96264 800 96292 1278
rect 96448 800 96476 1414
rect 96632 1414 96752 1442
rect 96632 800 96660 1414
rect 96816 800 96844 2926
rect 97000 800 97028 5714
rect 97264 4684 97316 4690
rect 97264 4626 97316 4632
rect 97276 800 97304 4626
rect 97460 4010 97488 9046
rect 97540 6656 97592 6662
rect 97540 6598 97592 6604
rect 97448 4004 97500 4010
rect 97448 3946 97500 3952
rect 97448 3460 97500 3466
rect 97448 3402 97500 3408
rect 97460 800 97488 3402
rect 97552 2922 97580 6598
rect 97632 6248 97684 6254
rect 97632 6190 97684 6196
rect 97540 2916 97592 2922
rect 97540 2858 97592 2864
rect 97644 800 97672 6190
rect 97736 3670 97764 22066
rect 97816 15088 97868 15094
rect 97816 15030 97868 15036
rect 97828 12918 97856 15030
rect 97920 14958 97948 96426
rect 98000 83360 98052 83366
rect 98000 83302 98052 83308
rect 98012 78674 98040 83302
rect 98000 78668 98052 78674
rect 98000 78610 98052 78616
rect 97908 14952 97960 14958
rect 97908 14894 97960 14900
rect 97816 12912 97868 12918
rect 97816 12854 97868 12860
rect 98276 6860 98328 6866
rect 98276 6802 98328 6808
rect 97816 5160 97868 5166
rect 97816 5102 97868 5108
rect 97724 3664 97776 3670
rect 97724 3606 97776 3612
rect 97724 2848 97776 2854
rect 97724 2790 97776 2796
rect 97736 2582 97764 2790
rect 97724 2576 97776 2582
rect 97724 2518 97776 2524
rect 97828 800 97856 5102
rect 98000 3936 98052 3942
rect 98000 3878 98052 3884
rect 98012 800 98040 3878
rect 98288 800 98316 6802
rect 98828 6180 98880 6186
rect 98828 6122 98880 6128
rect 98460 5092 98512 5098
rect 98460 5034 98512 5040
rect 98472 800 98500 5034
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 98656 800 98684 3470
rect 98840 800 98868 6122
rect 99012 5772 99064 5778
rect 99012 5714 99064 5720
rect 99024 800 99052 5714
rect 99472 5704 99524 5710
rect 99472 5646 99524 5652
rect 99288 4072 99340 4078
rect 99288 4014 99340 4020
rect 99300 800 99328 4014
rect 99484 800 99512 5646
rect 99840 2848 99892 2854
rect 99840 2790 99892 2796
rect 99656 2372 99708 2378
rect 99656 2314 99708 2320
rect 99668 800 99696 2314
rect 99852 800 99880 2790
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 13910 0 13966 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19338 0 19394 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36450 0 36506 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38658 0 38714 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40130 0 40186 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62026 0 62082 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63498 0 63554 800
rect 63682 0 63738 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65338 0 65394 800
rect 65522 0 65578 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67546 0 67602 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70766 0 70822 800
rect 71042 0 71098 800
rect 71226 0 71282 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73250 0 73306 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73802 0 73858 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74906 0 74962 800
rect 75090 0 75146 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76286 0 76342 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78770 0 78826 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81346 0 81402 800
rect 81530 0 81586 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83002 0 83058 800
rect 83186 0 83242 800
rect 83370 0 83426 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85026 0 85082 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88522 0 88578 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89258 0 89314 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 92938 0 92994 800
rect 93122 0 93178 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95146 0 95202 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< via2 >>
rect 1398 49952 1454 50008
rect 4220 96858 4276 96860
rect 4300 96858 4356 96860
rect 4380 96858 4436 96860
rect 4460 96858 4516 96860
rect 4220 96806 4246 96858
rect 4246 96806 4276 96858
rect 4300 96806 4310 96858
rect 4310 96806 4356 96858
rect 4380 96806 4426 96858
rect 4426 96806 4436 96858
rect 4460 96806 4490 96858
rect 4490 96806 4516 96858
rect 4220 96804 4276 96806
rect 4300 96804 4356 96806
rect 4380 96804 4436 96806
rect 4460 96804 4516 96806
rect 4220 95770 4276 95772
rect 4300 95770 4356 95772
rect 4380 95770 4436 95772
rect 4460 95770 4516 95772
rect 4220 95718 4246 95770
rect 4246 95718 4276 95770
rect 4300 95718 4310 95770
rect 4310 95718 4356 95770
rect 4380 95718 4426 95770
rect 4426 95718 4436 95770
rect 4460 95718 4490 95770
rect 4490 95718 4516 95770
rect 4220 95716 4276 95718
rect 4300 95716 4356 95718
rect 4380 95716 4436 95718
rect 4460 95716 4516 95718
rect 4220 94682 4276 94684
rect 4300 94682 4356 94684
rect 4380 94682 4436 94684
rect 4460 94682 4516 94684
rect 4220 94630 4246 94682
rect 4246 94630 4276 94682
rect 4300 94630 4310 94682
rect 4310 94630 4356 94682
rect 4380 94630 4426 94682
rect 4426 94630 4436 94682
rect 4460 94630 4490 94682
rect 4490 94630 4516 94682
rect 4220 94628 4276 94630
rect 4300 94628 4356 94630
rect 4380 94628 4436 94630
rect 4460 94628 4516 94630
rect 4220 93594 4276 93596
rect 4300 93594 4356 93596
rect 4380 93594 4436 93596
rect 4460 93594 4516 93596
rect 4220 93542 4246 93594
rect 4246 93542 4276 93594
rect 4300 93542 4310 93594
rect 4310 93542 4356 93594
rect 4380 93542 4426 93594
rect 4426 93542 4436 93594
rect 4460 93542 4490 93594
rect 4490 93542 4516 93594
rect 4220 93540 4276 93542
rect 4300 93540 4356 93542
rect 4380 93540 4436 93542
rect 4460 93540 4516 93542
rect 4220 92506 4276 92508
rect 4300 92506 4356 92508
rect 4380 92506 4436 92508
rect 4460 92506 4516 92508
rect 4220 92454 4246 92506
rect 4246 92454 4276 92506
rect 4300 92454 4310 92506
rect 4310 92454 4356 92506
rect 4380 92454 4426 92506
rect 4426 92454 4436 92506
rect 4460 92454 4490 92506
rect 4490 92454 4516 92506
rect 4220 92452 4276 92454
rect 4300 92452 4356 92454
rect 4380 92452 4436 92454
rect 4460 92452 4516 92454
rect 4220 91418 4276 91420
rect 4300 91418 4356 91420
rect 4380 91418 4436 91420
rect 4460 91418 4516 91420
rect 4220 91366 4246 91418
rect 4246 91366 4276 91418
rect 4300 91366 4310 91418
rect 4310 91366 4356 91418
rect 4380 91366 4426 91418
rect 4426 91366 4436 91418
rect 4460 91366 4490 91418
rect 4490 91366 4516 91418
rect 4220 91364 4276 91366
rect 4300 91364 4356 91366
rect 4380 91364 4436 91366
rect 4460 91364 4516 91366
rect 4220 90330 4276 90332
rect 4300 90330 4356 90332
rect 4380 90330 4436 90332
rect 4460 90330 4516 90332
rect 4220 90278 4246 90330
rect 4246 90278 4276 90330
rect 4300 90278 4310 90330
rect 4310 90278 4356 90330
rect 4380 90278 4426 90330
rect 4426 90278 4436 90330
rect 4460 90278 4490 90330
rect 4490 90278 4516 90330
rect 4220 90276 4276 90278
rect 4300 90276 4356 90278
rect 4380 90276 4436 90278
rect 4460 90276 4516 90278
rect 4220 89242 4276 89244
rect 4300 89242 4356 89244
rect 4380 89242 4436 89244
rect 4460 89242 4516 89244
rect 4220 89190 4246 89242
rect 4246 89190 4276 89242
rect 4300 89190 4310 89242
rect 4310 89190 4356 89242
rect 4380 89190 4426 89242
rect 4426 89190 4436 89242
rect 4460 89190 4490 89242
rect 4490 89190 4516 89242
rect 4220 89188 4276 89190
rect 4300 89188 4356 89190
rect 4380 89188 4436 89190
rect 4460 89188 4516 89190
rect 4220 88154 4276 88156
rect 4300 88154 4356 88156
rect 4380 88154 4436 88156
rect 4460 88154 4516 88156
rect 4220 88102 4246 88154
rect 4246 88102 4276 88154
rect 4300 88102 4310 88154
rect 4310 88102 4356 88154
rect 4380 88102 4426 88154
rect 4426 88102 4436 88154
rect 4460 88102 4490 88154
rect 4490 88102 4516 88154
rect 4220 88100 4276 88102
rect 4300 88100 4356 88102
rect 4380 88100 4436 88102
rect 4460 88100 4516 88102
rect 4220 87066 4276 87068
rect 4300 87066 4356 87068
rect 4380 87066 4436 87068
rect 4460 87066 4516 87068
rect 4220 87014 4246 87066
rect 4246 87014 4276 87066
rect 4300 87014 4310 87066
rect 4310 87014 4356 87066
rect 4380 87014 4426 87066
rect 4426 87014 4436 87066
rect 4460 87014 4490 87066
rect 4490 87014 4516 87066
rect 4220 87012 4276 87014
rect 4300 87012 4356 87014
rect 4380 87012 4436 87014
rect 4460 87012 4516 87014
rect 4220 85978 4276 85980
rect 4300 85978 4356 85980
rect 4380 85978 4436 85980
rect 4460 85978 4516 85980
rect 4220 85926 4246 85978
rect 4246 85926 4276 85978
rect 4300 85926 4310 85978
rect 4310 85926 4356 85978
rect 4380 85926 4426 85978
rect 4426 85926 4436 85978
rect 4460 85926 4490 85978
rect 4490 85926 4516 85978
rect 4220 85924 4276 85926
rect 4300 85924 4356 85926
rect 4380 85924 4436 85926
rect 4460 85924 4516 85926
rect 4220 84890 4276 84892
rect 4300 84890 4356 84892
rect 4380 84890 4436 84892
rect 4460 84890 4516 84892
rect 4220 84838 4246 84890
rect 4246 84838 4276 84890
rect 4300 84838 4310 84890
rect 4310 84838 4356 84890
rect 4380 84838 4426 84890
rect 4426 84838 4436 84890
rect 4460 84838 4490 84890
rect 4490 84838 4516 84890
rect 4220 84836 4276 84838
rect 4300 84836 4356 84838
rect 4380 84836 4436 84838
rect 4460 84836 4516 84838
rect 4220 83802 4276 83804
rect 4300 83802 4356 83804
rect 4380 83802 4436 83804
rect 4460 83802 4516 83804
rect 4220 83750 4246 83802
rect 4246 83750 4276 83802
rect 4300 83750 4310 83802
rect 4310 83750 4356 83802
rect 4380 83750 4426 83802
rect 4426 83750 4436 83802
rect 4460 83750 4490 83802
rect 4490 83750 4516 83802
rect 4220 83748 4276 83750
rect 4300 83748 4356 83750
rect 4380 83748 4436 83750
rect 4460 83748 4516 83750
rect 4220 82714 4276 82716
rect 4300 82714 4356 82716
rect 4380 82714 4436 82716
rect 4460 82714 4516 82716
rect 4220 82662 4246 82714
rect 4246 82662 4276 82714
rect 4300 82662 4310 82714
rect 4310 82662 4356 82714
rect 4380 82662 4426 82714
rect 4426 82662 4436 82714
rect 4460 82662 4490 82714
rect 4490 82662 4516 82714
rect 4220 82660 4276 82662
rect 4300 82660 4356 82662
rect 4380 82660 4436 82662
rect 4460 82660 4516 82662
rect 4220 81626 4276 81628
rect 4300 81626 4356 81628
rect 4380 81626 4436 81628
rect 4460 81626 4516 81628
rect 4220 81574 4246 81626
rect 4246 81574 4276 81626
rect 4300 81574 4310 81626
rect 4310 81574 4356 81626
rect 4380 81574 4426 81626
rect 4426 81574 4436 81626
rect 4460 81574 4490 81626
rect 4490 81574 4516 81626
rect 4220 81572 4276 81574
rect 4300 81572 4356 81574
rect 4380 81572 4436 81574
rect 4460 81572 4516 81574
rect 4220 80538 4276 80540
rect 4300 80538 4356 80540
rect 4380 80538 4436 80540
rect 4460 80538 4516 80540
rect 4220 80486 4246 80538
rect 4246 80486 4276 80538
rect 4300 80486 4310 80538
rect 4310 80486 4356 80538
rect 4380 80486 4426 80538
rect 4426 80486 4436 80538
rect 4460 80486 4490 80538
rect 4490 80486 4516 80538
rect 4220 80484 4276 80486
rect 4300 80484 4356 80486
rect 4380 80484 4436 80486
rect 4460 80484 4516 80486
rect 4220 79450 4276 79452
rect 4300 79450 4356 79452
rect 4380 79450 4436 79452
rect 4460 79450 4516 79452
rect 4220 79398 4246 79450
rect 4246 79398 4276 79450
rect 4300 79398 4310 79450
rect 4310 79398 4356 79450
rect 4380 79398 4426 79450
rect 4426 79398 4436 79450
rect 4460 79398 4490 79450
rect 4490 79398 4516 79450
rect 4220 79396 4276 79398
rect 4300 79396 4356 79398
rect 4380 79396 4436 79398
rect 4460 79396 4516 79398
rect 4220 78362 4276 78364
rect 4300 78362 4356 78364
rect 4380 78362 4436 78364
rect 4460 78362 4516 78364
rect 4220 78310 4246 78362
rect 4246 78310 4276 78362
rect 4300 78310 4310 78362
rect 4310 78310 4356 78362
rect 4380 78310 4426 78362
rect 4426 78310 4436 78362
rect 4460 78310 4490 78362
rect 4490 78310 4516 78362
rect 4220 78308 4276 78310
rect 4300 78308 4356 78310
rect 4380 78308 4436 78310
rect 4460 78308 4516 78310
rect 4220 77274 4276 77276
rect 4300 77274 4356 77276
rect 4380 77274 4436 77276
rect 4460 77274 4516 77276
rect 4220 77222 4246 77274
rect 4246 77222 4276 77274
rect 4300 77222 4310 77274
rect 4310 77222 4356 77274
rect 4380 77222 4426 77274
rect 4426 77222 4436 77274
rect 4460 77222 4490 77274
rect 4490 77222 4516 77274
rect 4220 77220 4276 77222
rect 4300 77220 4356 77222
rect 4380 77220 4436 77222
rect 4460 77220 4516 77222
rect 4220 76186 4276 76188
rect 4300 76186 4356 76188
rect 4380 76186 4436 76188
rect 4460 76186 4516 76188
rect 4220 76134 4246 76186
rect 4246 76134 4276 76186
rect 4300 76134 4310 76186
rect 4310 76134 4356 76186
rect 4380 76134 4426 76186
rect 4426 76134 4436 76186
rect 4460 76134 4490 76186
rect 4490 76134 4516 76186
rect 4220 76132 4276 76134
rect 4300 76132 4356 76134
rect 4380 76132 4436 76134
rect 4460 76132 4516 76134
rect 4220 75098 4276 75100
rect 4300 75098 4356 75100
rect 4380 75098 4436 75100
rect 4460 75098 4516 75100
rect 4220 75046 4246 75098
rect 4246 75046 4276 75098
rect 4300 75046 4310 75098
rect 4310 75046 4356 75098
rect 4380 75046 4426 75098
rect 4426 75046 4436 75098
rect 4460 75046 4490 75098
rect 4490 75046 4516 75098
rect 4220 75044 4276 75046
rect 4300 75044 4356 75046
rect 4380 75044 4436 75046
rect 4460 75044 4516 75046
rect 4220 74010 4276 74012
rect 4300 74010 4356 74012
rect 4380 74010 4436 74012
rect 4460 74010 4516 74012
rect 4220 73958 4246 74010
rect 4246 73958 4276 74010
rect 4300 73958 4310 74010
rect 4310 73958 4356 74010
rect 4380 73958 4426 74010
rect 4426 73958 4436 74010
rect 4460 73958 4490 74010
rect 4490 73958 4516 74010
rect 4220 73956 4276 73958
rect 4300 73956 4356 73958
rect 4380 73956 4436 73958
rect 4460 73956 4516 73958
rect 4220 72922 4276 72924
rect 4300 72922 4356 72924
rect 4380 72922 4436 72924
rect 4460 72922 4516 72924
rect 4220 72870 4246 72922
rect 4246 72870 4276 72922
rect 4300 72870 4310 72922
rect 4310 72870 4356 72922
rect 4380 72870 4426 72922
rect 4426 72870 4436 72922
rect 4460 72870 4490 72922
rect 4490 72870 4516 72922
rect 4220 72868 4276 72870
rect 4300 72868 4356 72870
rect 4380 72868 4436 72870
rect 4460 72868 4516 72870
rect 4220 71834 4276 71836
rect 4300 71834 4356 71836
rect 4380 71834 4436 71836
rect 4460 71834 4516 71836
rect 4220 71782 4246 71834
rect 4246 71782 4276 71834
rect 4300 71782 4310 71834
rect 4310 71782 4356 71834
rect 4380 71782 4426 71834
rect 4426 71782 4436 71834
rect 4460 71782 4490 71834
rect 4490 71782 4516 71834
rect 4220 71780 4276 71782
rect 4300 71780 4356 71782
rect 4380 71780 4436 71782
rect 4460 71780 4516 71782
rect 4220 70746 4276 70748
rect 4300 70746 4356 70748
rect 4380 70746 4436 70748
rect 4460 70746 4516 70748
rect 4220 70694 4246 70746
rect 4246 70694 4276 70746
rect 4300 70694 4310 70746
rect 4310 70694 4356 70746
rect 4380 70694 4426 70746
rect 4426 70694 4436 70746
rect 4460 70694 4490 70746
rect 4490 70694 4516 70746
rect 4220 70692 4276 70694
rect 4300 70692 4356 70694
rect 4380 70692 4436 70694
rect 4460 70692 4516 70694
rect 4220 69658 4276 69660
rect 4300 69658 4356 69660
rect 4380 69658 4436 69660
rect 4460 69658 4516 69660
rect 4220 69606 4246 69658
rect 4246 69606 4276 69658
rect 4300 69606 4310 69658
rect 4310 69606 4356 69658
rect 4380 69606 4426 69658
rect 4426 69606 4436 69658
rect 4460 69606 4490 69658
rect 4490 69606 4516 69658
rect 4220 69604 4276 69606
rect 4300 69604 4356 69606
rect 4380 69604 4436 69606
rect 4460 69604 4516 69606
rect 4220 68570 4276 68572
rect 4300 68570 4356 68572
rect 4380 68570 4436 68572
rect 4460 68570 4516 68572
rect 4220 68518 4246 68570
rect 4246 68518 4276 68570
rect 4300 68518 4310 68570
rect 4310 68518 4356 68570
rect 4380 68518 4426 68570
rect 4426 68518 4436 68570
rect 4460 68518 4490 68570
rect 4490 68518 4516 68570
rect 4220 68516 4276 68518
rect 4300 68516 4356 68518
rect 4380 68516 4436 68518
rect 4460 68516 4516 68518
rect 4220 67482 4276 67484
rect 4300 67482 4356 67484
rect 4380 67482 4436 67484
rect 4460 67482 4516 67484
rect 4220 67430 4246 67482
rect 4246 67430 4276 67482
rect 4300 67430 4310 67482
rect 4310 67430 4356 67482
rect 4380 67430 4426 67482
rect 4426 67430 4436 67482
rect 4460 67430 4490 67482
rect 4490 67430 4516 67482
rect 4220 67428 4276 67430
rect 4300 67428 4356 67430
rect 4380 67428 4436 67430
rect 4460 67428 4516 67430
rect 3974 67124 3976 67144
rect 3976 67124 4028 67144
rect 4028 67124 4030 67144
rect 3974 67088 4030 67124
rect 4220 66394 4276 66396
rect 4300 66394 4356 66396
rect 4380 66394 4436 66396
rect 4460 66394 4516 66396
rect 4220 66342 4246 66394
rect 4246 66342 4276 66394
rect 4300 66342 4310 66394
rect 4310 66342 4356 66394
rect 4380 66342 4426 66394
rect 4426 66342 4436 66394
rect 4460 66342 4490 66394
rect 4490 66342 4516 66394
rect 4220 66340 4276 66342
rect 4300 66340 4356 66342
rect 4380 66340 4436 66342
rect 4460 66340 4516 66342
rect 4220 65306 4276 65308
rect 4300 65306 4356 65308
rect 4380 65306 4436 65308
rect 4460 65306 4516 65308
rect 4220 65254 4246 65306
rect 4246 65254 4276 65306
rect 4300 65254 4310 65306
rect 4310 65254 4356 65306
rect 4380 65254 4426 65306
rect 4426 65254 4436 65306
rect 4460 65254 4490 65306
rect 4490 65254 4516 65306
rect 4220 65252 4276 65254
rect 4300 65252 4356 65254
rect 4380 65252 4436 65254
rect 4460 65252 4516 65254
rect 4220 64218 4276 64220
rect 4300 64218 4356 64220
rect 4380 64218 4436 64220
rect 4460 64218 4516 64220
rect 4220 64166 4246 64218
rect 4246 64166 4276 64218
rect 4300 64166 4310 64218
rect 4310 64166 4356 64218
rect 4380 64166 4426 64218
rect 4426 64166 4436 64218
rect 4460 64166 4490 64218
rect 4490 64166 4516 64218
rect 4220 64164 4276 64166
rect 4300 64164 4356 64166
rect 4380 64164 4436 64166
rect 4460 64164 4516 64166
rect 4220 63130 4276 63132
rect 4300 63130 4356 63132
rect 4380 63130 4436 63132
rect 4460 63130 4516 63132
rect 4220 63078 4246 63130
rect 4246 63078 4276 63130
rect 4300 63078 4310 63130
rect 4310 63078 4356 63130
rect 4380 63078 4426 63130
rect 4426 63078 4436 63130
rect 4460 63078 4490 63130
rect 4490 63078 4516 63130
rect 4220 63076 4276 63078
rect 4300 63076 4356 63078
rect 4380 63076 4436 63078
rect 4460 63076 4516 63078
rect 4220 62042 4276 62044
rect 4300 62042 4356 62044
rect 4380 62042 4436 62044
rect 4460 62042 4516 62044
rect 4220 61990 4246 62042
rect 4246 61990 4276 62042
rect 4300 61990 4310 62042
rect 4310 61990 4356 62042
rect 4380 61990 4426 62042
rect 4426 61990 4436 62042
rect 4460 61990 4490 62042
rect 4490 61990 4516 62042
rect 4220 61988 4276 61990
rect 4300 61988 4356 61990
rect 4380 61988 4436 61990
rect 4460 61988 4516 61990
rect 4220 60954 4276 60956
rect 4300 60954 4356 60956
rect 4380 60954 4436 60956
rect 4460 60954 4516 60956
rect 4220 60902 4246 60954
rect 4246 60902 4276 60954
rect 4300 60902 4310 60954
rect 4310 60902 4356 60954
rect 4380 60902 4426 60954
rect 4426 60902 4436 60954
rect 4460 60902 4490 60954
rect 4490 60902 4516 60954
rect 4220 60900 4276 60902
rect 4300 60900 4356 60902
rect 4380 60900 4436 60902
rect 4460 60900 4516 60902
rect 4220 59866 4276 59868
rect 4300 59866 4356 59868
rect 4380 59866 4436 59868
rect 4460 59866 4516 59868
rect 4220 59814 4246 59866
rect 4246 59814 4276 59866
rect 4300 59814 4310 59866
rect 4310 59814 4356 59866
rect 4380 59814 4426 59866
rect 4426 59814 4436 59866
rect 4460 59814 4490 59866
rect 4490 59814 4516 59866
rect 4220 59812 4276 59814
rect 4300 59812 4356 59814
rect 4380 59812 4436 59814
rect 4460 59812 4516 59814
rect 4220 58778 4276 58780
rect 4300 58778 4356 58780
rect 4380 58778 4436 58780
rect 4460 58778 4516 58780
rect 4220 58726 4246 58778
rect 4246 58726 4276 58778
rect 4300 58726 4310 58778
rect 4310 58726 4356 58778
rect 4380 58726 4426 58778
rect 4426 58726 4436 58778
rect 4460 58726 4490 58778
rect 4490 58726 4516 58778
rect 4220 58724 4276 58726
rect 4300 58724 4356 58726
rect 4380 58724 4436 58726
rect 4460 58724 4516 58726
rect 4220 57690 4276 57692
rect 4300 57690 4356 57692
rect 4380 57690 4436 57692
rect 4460 57690 4516 57692
rect 4220 57638 4246 57690
rect 4246 57638 4276 57690
rect 4300 57638 4310 57690
rect 4310 57638 4356 57690
rect 4380 57638 4426 57690
rect 4426 57638 4436 57690
rect 4460 57638 4490 57690
rect 4490 57638 4516 57690
rect 4220 57636 4276 57638
rect 4300 57636 4356 57638
rect 4380 57636 4436 57638
rect 4460 57636 4516 57638
rect 4220 56602 4276 56604
rect 4300 56602 4356 56604
rect 4380 56602 4436 56604
rect 4460 56602 4516 56604
rect 4220 56550 4246 56602
rect 4246 56550 4276 56602
rect 4300 56550 4310 56602
rect 4310 56550 4356 56602
rect 4380 56550 4426 56602
rect 4426 56550 4436 56602
rect 4460 56550 4490 56602
rect 4490 56550 4516 56602
rect 4220 56548 4276 56550
rect 4300 56548 4356 56550
rect 4380 56548 4436 56550
rect 4460 56548 4516 56550
rect 4220 55514 4276 55516
rect 4300 55514 4356 55516
rect 4380 55514 4436 55516
rect 4460 55514 4516 55516
rect 4220 55462 4246 55514
rect 4246 55462 4276 55514
rect 4300 55462 4310 55514
rect 4310 55462 4356 55514
rect 4380 55462 4426 55514
rect 4426 55462 4436 55514
rect 4460 55462 4490 55514
rect 4490 55462 4516 55514
rect 4220 55460 4276 55462
rect 4300 55460 4356 55462
rect 4380 55460 4436 55462
rect 4460 55460 4516 55462
rect 4220 54426 4276 54428
rect 4300 54426 4356 54428
rect 4380 54426 4436 54428
rect 4460 54426 4516 54428
rect 4220 54374 4246 54426
rect 4246 54374 4276 54426
rect 4300 54374 4310 54426
rect 4310 54374 4356 54426
rect 4380 54374 4426 54426
rect 4426 54374 4436 54426
rect 4460 54374 4490 54426
rect 4490 54374 4516 54426
rect 4220 54372 4276 54374
rect 4300 54372 4356 54374
rect 4380 54372 4436 54374
rect 4460 54372 4516 54374
rect 4220 53338 4276 53340
rect 4300 53338 4356 53340
rect 4380 53338 4436 53340
rect 4460 53338 4516 53340
rect 4220 53286 4246 53338
rect 4246 53286 4276 53338
rect 4300 53286 4310 53338
rect 4310 53286 4356 53338
rect 4380 53286 4426 53338
rect 4426 53286 4436 53338
rect 4460 53286 4490 53338
rect 4490 53286 4516 53338
rect 4220 53284 4276 53286
rect 4300 53284 4356 53286
rect 4380 53284 4436 53286
rect 4460 53284 4516 53286
rect 4220 52250 4276 52252
rect 4300 52250 4356 52252
rect 4380 52250 4436 52252
rect 4460 52250 4516 52252
rect 4220 52198 4246 52250
rect 4246 52198 4276 52250
rect 4300 52198 4310 52250
rect 4310 52198 4356 52250
rect 4380 52198 4426 52250
rect 4426 52198 4436 52250
rect 4460 52198 4490 52250
rect 4490 52198 4516 52250
rect 4220 52196 4276 52198
rect 4300 52196 4356 52198
rect 4380 52196 4436 52198
rect 4460 52196 4516 52198
rect 4220 51162 4276 51164
rect 4300 51162 4356 51164
rect 4380 51162 4436 51164
rect 4460 51162 4516 51164
rect 4220 51110 4246 51162
rect 4246 51110 4276 51162
rect 4300 51110 4310 51162
rect 4310 51110 4356 51162
rect 4380 51110 4426 51162
rect 4426 51110 4436 51162
rect 4460 51110 4490 51162
rect 4490 51110 4516 51162
rect 4220 51108 4276 51110
rect 4300 51108 4356 51110
rect 4380 51108 4436 51110
rect 4460 51108 4516 51110
rect 4220 50074 4276 50076
rect 4300 50074 4356 50076
rect 4380 50074 4436 50076
rect 4460 50074 4516 50076
rect 4220 50022 4246 50074
rect 4246 50022 4276 50074
rect 4300 50022 4310 50074
rect 4310 50022 4356 50074
rect 4380 50022 4426 50074
rect 4426 50022 4436 50074
rect 4460 50022 4490 50074
rect 4490 50022 4516 50074
rect 4220 50020 4276 50022
rect 4300 50020 4356 50022
rect 4380 50020 4436 50022
rect 4460 50020 4516 50022
rect 4220 48986 4276 48988
rect 4300 48986 4356 48988
rect 4380 48986 4436 48988
rect 4460 48986 4516 48988
rect 4220 48934 4246 48986
rect 4246 48934 4276 48986
rect 4300 48934 4310 48986
rect 4310 48934 4356 48986
rect 4380 48934 4426 48986
rect 4426 48934 4436 48986
rect 4460 48934 4490 48986
rect 4490 48934 4516 48986
rect 4220 48932 4276 48934
rect 4300 48932 4356 48934
rect 4380 48932 4436 48934
rect 4460 48932 4516 48934
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4246 47898
rect 4246 47846 4276 47898
rect 4300 47846 4310 47898
rect 4310 47846 4356 47898
rect 4380 47846 4426 47898
rect 4426 47846 4436 47898
rect 4460 47846 4490 47898
rect 4490 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 5170 67088 5226 67144
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 10046 85196 10102 85232
rect 10046 85176 10048 85196
rect 10048 85176 10100 85196
rect 10100 85176 10102 85196
rect 14646 85176 14702 85232
rect 19580 97402 19636 97404
rect 19660 97402 19716 97404
rect 19740 97402 19796 97404
rect 19820 97402 19876 97404
rect 19580 97350 19606 97402
rect 19606 97350 19636 97402
rect 19660 97350 19670 97402
rect 19670 97350 19716 97402
rect 19740 97350 19786 97402
rect 19786 97350 19796 97402
rect 19820 97350 19850 97402
rect 19850 97350 19876 97402
rect 19580 97348 19636 97350
rect 19660 97348 19716 97350
rect 19740 97348 19796 97350
rect 19820 97348 19876 97350
rect 19580 96314 19636 96316
rect 19660 96314 19716 96316
rect 19740 96314 19796 96316
rect 19820 96314 19876 96316
rect 19580 96262 19606 96314
rect 19606 96262 19636 96314
rect 19660 96262 19670 96314
rect 19670 96262 19716 96314
rect 19740 96262 19786 96314
rect 19786 96262 19796 96314
rect 19820 96262 19850 96314
rect 19850 96262 19876 96314
rect 19580 96260 19636 96262
rect 19660 96260 19716 96262
rect 19740 96260 19796 96262
rect 19820 96260 19876 96262
rect 19580 95226 19636 95228
rect 19660 95226 19716 95228
rect 19740 95226 19796 95228
rect 19820 95226 19876 95228
rect 19580 95174 19606 95226
rect 19606 95174 19636 95226
rect 19660 95174 19670 95226
rect 19670 95174 19716 95226
rect 19740 95174 19786 95226
rect 19786 95174 19796 95226
rect 19820 95174 19850 95226
rect 19850 95174 19876 95226
rect 19580 95172 19636 95174
rect 19660 95172 19716 95174
rect 19740 95172 19796 95174
rect 19820 95172 19876 95174
rect 19580 94138 19636 94140
rect 19660 94138 19716 94140
rect 19740 94138 19796 94140
rect 19820 94138 19876 94140
rect 19580 94086 19606 94138
rect 19606 94086 19636 94138
rect 19660 94086 19670 94138
rect 19670 94086 19716 94138
rect 19740 94086 19786 94138
rect 19786 94086 19796 94138
rect 19820 94086 19850 94138
rect 19850 94086 19876 94138
rect 19580 94084 19636 94086
rect 19660 94084 19716 94086
rect 19740 94084 19796 94086
rect 19820 94084 19876 94086
rect 19580 93050 19636 93052
rect 19660 93050 19716 93052
rect 19740 93050 19796 93052
rect 19820 93050 19876 93052
rect 19580 92998 19606 93050
rect 19606 92998 19636 93050
rect 19660 92998 19670 93050
rect 19670 92998 19716 93050
rect 19740 92998 19786 93050
rect 19786 92998 19796 93050
rect 19820 92998 19850 93050
rect 19850 92998 19876 93050
rect 19580 92996 19636 92998
rect 19660 92996 19716 92998
rect 19740 92996 19796 92998
rect 19820 92996 19876 92998
rect 19580 91962 19636 91964
rect 19660 91962 19716 91964
rect 19740 91962 19796 91964
rect 19820 91962 19876 91964
rect 19580 91910 19606 91962
rect 19606 91910 19636 91962
rect 19660 91910 19670 91962
rect 19670 91910 19716 91962
rect 19740 91910 19786 91962
rect 19786 91910 19796 91962
rect 19820 91910 19850 91962
rect 19850 91910 19876 91962
rect 19580 91908 19636 91910
rect 19660 91908 19716 91910
rect 19740 91908 19796 91910
rect 19820 91908 19876 91910
rect 19580 90874 19636 90876
rect 19660 90874 19716 90876
rect 19740 90874 19796 90876
rect 19820 90874 19876 90876
rect 19580 90822 19606 90874
rect 19606 90822 19636 90874
rect 19660 90822 19670 90874
rect 19670 90822 19716 90874
rect 19740 90822 19786 90874
rect 19786 90822 19796 90874
rect 19820 90822 19850 90874
rect 19850 90822 19876 90874
rect 19580 90820 19636 90822
rect 19660 90820 19716 90822
rect 19740 90820 19796 90822
rect 19820 90820 19876 90822
rect 19580 89786 19636 89788
rect 19660 89786 19716 89788
rect 19740 89786 19796 89788
rect 19820 89786 19876 89788
rect 19580 89734 19606 89786
rect 19606 89734 19636 89786
rect 19660 89734 19670 89786
rect 19670 89734 19716 89786
rect 19740 89734 19786 89786
rect 19786 89734 19796 89786
rect 19820 89734 19850 89786
rect 19850 89734 19876 89786
rect 19580 89732 19636 89734
rect 19660 89732 19716 89734
rect 19740 89732 19796 89734
rect 19820 89732 19876 89734
rect 19580 88698 19636 88700
rect 19660 88698 19716 88700
rect 19740 88698 19796 88700
rect 19820 88698 19876 88700
rect 19580 88646 19606 88698
rect 19606 88646 19636 88698
rect 19660 88646 19670 88698
rect 19670 88646 19716 88698
rect 19740 88646 19786 88698
rect 19786 88646 19796 88698
rect 19820 88646 19850 88698
rect 19850 88646 19876 88698
rect 19580 88644 19636 88646
rect 19660 88644 19716 88646
rect 19740 88644 19796 88646
rect 19820 88644 19876 88646
rect 19580 87610 19636 87612
rect 19660 87610 19716 87612
rect 19740 87610 19796 87612
rect 19820 87610 19876 87612
rect 19580 87558 19606 87610
rect 19606 87558 19636 87610
rect 19660 87558 19670 87610
rect 19670 87558 19716 87610
rect 19740 87558 19786 87610
rect 19786 87558 19796 87610
rect 19820 87558 19850 87610
rect 19850 87558 19876 87610
rect 19580 87556 19636 87558
rect 19660 87556 19716 87558
rect 19740 87556 19796 87558
rect 19820 87556 19876 87558
rect 19580 86522 19636 86524
rect 19660 86522 19716 86524
rect 19740 86522 19796 86524
rect 19820 86522 19876 86524
rect 19580 86470 19606 86522
rect 19606 86470 19636 86522
rect 19660 86470 19670 86522
rect 19670 86470 19716 86522
rect 19740 86470 19786 86522
rect 19786 86470 19796 86522
rect 19820 86470 19850 86522
rect 19850 86470 19876 86522
rect 19580 86468 19636 86470
rect 19660 86468 19716 86470
rect 19740 86468 19796 86470
rect 19820 86468 19876 86470
rect 19580 85434 19636 85436
rect 19660 85434 19716 85436
rect 19740 85434 19796 85436
rect 19820 85434 19876 85436
rect 19580 85382 19606 85434
rect 19606 85382 19636 85434
rect 19660 85382 19670 85434
rect 19670 85382 19716 85434
rect 19740 85382 19786 85434
rect 19786 85382 19796 85434
rect 19820 85382 19850 85434
rect 19850 85382 19876 85434
rect 19580 85380 19636 85382
rect 19660 85380 19716 85382
rect 19740 85380 19796 85382
rect 19820 85380 19876 85382
rect 19580 84346 19636 84348
rect 19660 84346 19716 84348
rect 19740 84346 19796 84348
rect 19820 84346 19876 84348
rect 19580 84294 19606 84346
rect 19606 84294 19636 84346
rect 19660 84294 19670 84346
rect 19670 84294 19716 84346
rect 19740 84294 19786 84346
rect 19786 84294 19796 84346
rect 19820 84294 19850 84346
rect 19850 84294 19876 84346
rect 19580 84292 19636 84294
rect 19660 84292 19716 84294
rect 19740 84292 19796 84294
rect 19820 84292 19876 84294
rect 19580 83258 19636 83260
rect 19660 83258 19716 83260
rect 19740 83258 19796 83260
rect 19820 83258 19876 83260
rect 19580 83206 19606 83258
rect 19606 83206 19636 83258
rect 19660 83206 19670 83258
rect 19670 83206 19716 83258
rect 19740 83206 19786 83258
rect 19786 83206 19796 83258
rect 19820 83206 19850 83258
rect 19850 83206 19876 83258
rect 19580 83204 19636 83206
rect 19660 83204 19716 83206
rect 19740 83204 19796 83206
rect 19820 83204 19876 83206
rect 19580 82170 19636 82172
rect 19660 82170 19716 82172
rect 19740 82170 19796 82172
rect 19820 82170 19876 82172
rect 19580 82118 19606 82170
rect 19606 82118 19636 82170
rect 19660 82118 19670 82170
rect 19670 82118 19716 82170
rect 19740 82118 19786 82170
rect 19786 82118 19796 82170
rect 19820 82118 19850 82170
rect 19850 82118 19876 82170
rect 19580 82116 19636 82118
rect 19660 82116 19716 82118
rect 19740 82116 19796 82118
rect 19820 82116 19876 82118
rect 19580 81082 19636 81084
rect 19660 81082 19716 81084
rect 19740 81082 19796 81084
rect 19820 81082 19876 81084
rect 19580 81030 19606 81082
rect 19606 81030 19636 81082
rect 19660 81030 19670 81082
rect 19670 81030 19716 81082
rect 19740 81030 19786 81082
rect 19786 81030 19796 81082
rect 19820 81030 19850 81082
rect 19850 81030 19876 81082
rect 19580 81028 19636 81030
rect 19660 81028 19716 81030
rect 19740 81028 19796 81030
rect 19820 81028 19876 81030
rect 19580 79994 19636 79996
rect 19660 79994 19716 79996
rect 19740 79994 19796 79996
rect 19820 79994 19876 79996
rect 19580 79942 19606 79994
rect 19606 79942 19636 79994
rect 19660 79942 19670 79994
rect 19670 79942 19716 79994
rect 19740 79942 19786 79994
rect 19786 79942 19796 79994
rect 19820 79942 19850 79994
rect 19850 79942 19876 79994
rect 19580 79940 19636 79942
rect 19660 79940 19716 79942
rect 19740 79940 19796 79942
rect 19820 79940 19876 79942
rect 19580 78906 19636 78908
rect 19660 78906 19716 78908
rect 19740 78906 19796 78908
rect 19820 78906 19876 78908
rect 19580 78854 19606 78906
rect 19606 78854 19636 78906
rect 19660 78854 19670 78906
rect 19670 78854 19716 78906
rect 19740 78854 19786 78906
rect 19786 78854 19796 78906
rect 19820 78854 19850 78906
rect 19850 78854 19876 78906
rect 19580 78852 19636 78854
rect 19660 78852 19716 78854
rect 19740 78852 19796 78854
rect 19820 78852 19876 78854
rect 19580 77818 19636 77820
rect 19660 77818 19716 77820
rect 19740 77818 19796 77820
rect 19820 77818 19876 77820
rect 19580 77766 19606 77818
rect 19606 77766 19636 77818
rect 19660 77766 19670 77818
rect 19670 77766 19716 77818
rect 19740 77766 19786 77818
rect 19786 77766 19796 77818
rect 19820 77766 19850 77818
rect 19850 77766 19876 77818
rect 19580 77764 19636 77766
rect 19660 77764 19716 77766
rect 19740 77764 19796 77766
rect 19820 77764 19876 77766
rect 19580 76730 19636 76732
rect 19660 76730 19716 76732
rect 19740 76730 19796 76732
rect 19820 76730 19876 76732
rect 19580 76678 19606 76730
rect 19606 76678 19636 76730
rect 19660 76678 19670 76730
rect 19670 76678 19716 76730
rect 19740 76678 19786 76730
rect 19786 76678 19796 76730
rect 19820 76678 19850 76730
rect 19850 76678 19876 76730
rect 19580 76676 19636 76678
rect 19660 76676 19716 76678
rect 19740 76676 19796 76678
rect 19820 76676 19876 76678
rect 19580 75642 19636 75644
rect 19660 75642 19716 75644
rect 19740 75642 19796 75644
rect 19820 75642 19876 75644
rect 19580 75590 19606 75642
rect 19606 75590 19636 75642
rect 19660 75590 19670 75642
rect 19670 75590 19716 75642
rect 19740 75590 19786 75642
rect 19786 75590 19796 75642
rect 19820 75590 19850 75642
rect 19850 75590 19876 75642
rect 19580 75588 19636 75590
rect 19660 75588 19716 75590
rect 19740 75588 19796 75590
rect 19820 75588 19876 75590
rect 19580 74554 19636 74556
rect 19660 74554 19716 74556
rect 19740 74554 19796 74556
rect 19820 74554 19876 74556
rect 19580 74502 19606 74554
rect 19606 74502 19636 74554
rect 19660 74502 19670 74554
rect 19670 74502 19716 74554
rect 19740 74502 19786 74554
rect 19786 74502 19796 74554
rect 19820 74502 19850 74554
rect 19850 74502 19876 74554
rect 19580 74500 19636 74502
rect 19660 74500 19716 74502
rect 19740 74500 19796 74502
rect 19820 74500 19876 74502
rect 19580 73466 19636 73468
rect 19660 73466 19716 73468
rect 19740 73466 19796 73468
rect 19820 73466 19876 73468
rect 19580 73414 19606 73466
rect 19606 73414 19636 73466
rect 19660 73414 19670 73466
rect 19670 73414 19716 73466
rect 19740 73414 19786 73466
rect 19786 73414 19796 73466
rect 19820 73414 19850 73466
rect 19850 73414 19876 73466
rect 19580 73412 19636 73414
rect 19660 73412 19716 73414
rect 19740 73412 19796 73414
rect 19820 73412 19876 73414
rect 19580 72378 19636 72380
rect 19660 72378 19716 72380
rect 19740 72378 19796 72380
rect 19820 72378 19876 72380
rect 19580 72326 19606 72378
rect 19606 72326 19636 72378
rect 19660 72326 19670 72378
rect 19670 72326 19716 72378
rect 19740 72326 19786 72378
rect 19786 72326 19796 72378
rect 19820 72326 19850 72378
rect 19850 72326 19876 72378
rect 19580 72324 19636 72326
rect 19660 72324 19716 72326
rect 19740 72324 19796 72326
rect 19820 72324 19876 72326
rect 19580 71290 19636 71292
rect 19660 71290 19716 71292
rect 19740 71290 19796 71292
rect 19820 71290 19876 71292
rect 19580 71238 19606 71290
rect 19606 71238 19636 71290
rect 19660 71238 19670 71290
rect 19670 71238 19716 71290
rect 19740 71238 19786 71290
rect 19786 71238 19796 71290
rect 19820 71238 19850 71290
rect 19850 71238 19876 71290
rect 19580 71236 19636 71238
rect 19660 71236 19716 71238
rect 19740 71236 19796 71238
rect 19820 71236 19876 71238
rect 19580 70202 19636 70204
rect 19660 70202 19716 70204
rect 19740 70202 19796 70204
rect 19820 70202 19876 70204
rect 19580 70150 19606 70202
rect 19606 70150 19636 70202
rect 19660 70150 19670 70202
rect 19670 70150 19716 70202
rect 19740 70150 19786 70202
rect 19786 70150 19796 70202
rect 19820 70150 19850 70202
rect 19850 70150 19876 70202
rect 19580 70148 19636 70150
rect 19660 70148 19716 70150
rect 19740 70148 19796 70150
rect 19820 70148 19876 70150
rect 19580 69114 19636 69116
rect 19660 69114 19716 69116
rect 19740 69114 19796 69116
rect 19820 69114 19876 69116
rect 19580 69062 19606 69114
rect 19606 69062 19636 69114
rect 19660 69062 19670 69114
rect 19670 69062 19716 69114
rect 19740 69062 19786 69114
rect 19786 69062 19796 69114
rect 19820 69062 19850 69114
rect 19850 69062 19876 69114
rect 19580 69060 19636 69062
rect 19660 69060 19716 69062
rect 19740 69060 19796 69062
rect 19820 69060 19876 69062
rect 19580 68026 19636 68028
rect 19660 68026 19716 68028
rect 19740 68026 19796 68028
rect 19820 68026 19876 68028
rect 19580 67974 19606 68026
rect 19606 67974 19636 68026
rect 19660 67974 19670 68026
rect 19670 67974 19716 68026
rect 19740 67974 19786 68026
rect 19786 67974 19796 68026
rect 19820 67974 19850 68026
rect 19850 67974 19876 68026
rect 19580 67972 19636 67974
rect 19660 67972 19716 67974
rect 19740 67972 19796 67974
rect 19820 67972 19876 67974
rect 19580 66938 19636 66940
rect 19660 66938 19716 66940
rect 19740 66938 19796 66940
rect 19820 66938 19876 66940
rect 19580 66886 19606 66938
rect 19606 66886 19636 66938
rect 19660 66886 19670 66938
rect 19670 66886 19716 66938
rect 19740 66886 19786 66938
rect 19786 66886 19796 66938
rect 19820 66886 19850 66938
rect 19850 66886 19876 66938
rect 19580 66884 19636 66886
rect 19660 66884 19716 66886
rect 19740 66884 19796 66886
rect 19820 66884 19876 66886
rect 19580 65850 19636 65852
rect 19660 65850 19716 65852
rect 19740 65850 19796 65852
rect 19820 65850 19876 65852
rect 19580 65798 19606 65850
rect 19606 65798 19636 65850
rect 19660 65798 19670 65850
rect 19670 65798 19716 65850
rect 19740 65798 19786 65850
rect 19786 65798 19796 65850
rect 19820 65798 19850 65850
rect 19850 65798 19876 65850
rect 19580 65796 19636 65798
rect 19660 65796 19716 65798
rect 19740 65796 19796 65798
rect 19820 65796 19876 65798
rect 19580 64762 19636 64764
rect 19660 64762 19716 64764
rect 19740 64762 19796 64764
rect 19820 64762 19876 64764
rect 19580 64710 19606 64762
rect 19606 64710 19636 64762
rect 19660 64710 19670 64762
rect 19670 64710 19716 64762
rect 19740 64710 19786 64762
rect 19786 64710 19796 64762
rect 19820 64710 19850 64762
rect 19850 64710 19876 64762
rect 19580 64708 19636 64710
rect 19660 64708 19716 64710
rect 19740 64708 19796 64710
rect 19820 64708 19876 64710
rect 19580 63674 19636 63676
rect 19660 63674 19716 63676
rect 19740 63674 19796 63676
rect 19820 63674 19876 63676
rect 19580 63622 19606 63674
rect 19606 63622 19636 63674
rect 19660 63622 19670 63674
rect 19670 63622 19716 63674
rect 19740 63622 19786 63674
rect 19786 63622 19796 63674
rect 19820 63622 19850 63674
rect 19850 63622 19876 63674
rect 19580 63620 19636 63622
rect 19660 63620 19716 63622
rect 19740 63620 19796 63622
rect 19820 63620 19876 63622
rect 19580 62586 19636 62588
rect 19660 62586 19716 62588
rect 19740 62586 19796 62588
rect 19820 62586 19876 62588
rect 19580 62534 19606 62586
rect 19606 62534 19636 62586
rect 19660 62534 19670 62586
rect 19670 62534 19716 62586
rect 19740 62534 19786 62586
rect 19786 62534 19796 62586
rect 19820 62534 19850 62586
rect 19850 62534 19876 62586
rect 19580 62532 19636 62534
rect 19660 62532 19716 62534
rect 19740 62532 19796 62534
rect 19820 62532 19876 62534
rect 19580 61498 19636 61500
rect 19660 61498 19716 61500
rect 19740 61498 19796 61500
rect 19820 61498 19876 61500
rect 19580 61446 19606 61498
rect 19606 61446 19636 61498
rect 19660 61446 19670 61498
rect 19670 61446 19716 61498
rect 19740 61446 19786 61498
rect 19786 61446 19796 61498
rect 19820 61446 19850 61498
rect 19850 61446 19876 61498
rect 19580 61444 19636 61446
rect 19660 61444 19716 61446
rect 19740 61444 19796 61446
rect 19820 61444 19876 61446
rect 19580 60410 19636 60412
rect 19660 60410 19716 60412
rect 19740 60410 19796 60412
rect 19820 60410 19876 60412
rect 19580 60358 19606 60410
rect 19606 60358 19636 60410
rect 19660 60358 19670 60410
rect 19670 60358 19716 60410
rect 19740 60358 19786 60410
rect 19786 60358 19796 60410
rect 19820 60358 19850 60410
rect 19850 60358 19876 60410
rect 19580 60356 19636 60358
rect 19660 60356 19716 60358
rect 19740 60356 19796 60358
rect 19820 60356 19876 60358
rect 19580 59322 19636 59324
rect 19660 59322 19716 59324
rect 19740 59322 19796 59324
rect 19820 59322 19876 59324
rect 19580 59270 19606 59322
rect 19606 59270 19636 59322
rect 19660 59270 19670 59322
rect 19670 59270 19716 59322
rect 19740 59270 19786 59322
rect 19786 59270 19796 59322
rect 19820 59270 19850 59322
rect 19850 59270 19876 59322
rect 19580 59268 19636 59270
rect 19660 59268 19716 59270
rect 19740 59268 19796 59270
rect 19820 59268 19876 59270
rect 19580 58234 19636 58236
rect 19660 58234 19716 58236
rect 19740 58234 19796 58236
rect 19820 58234 19876 58236
rect 19580 58182 19606 58234
rect 19606 58182 19636 58234
rect 19660 58182 19670 58234
rect 19670 58182 19716 58234
rect 19740 58182 19786 58234
rect 19786 58182 19796 58234
rect 19820 58182 19850 58234
rect 19850 58182 19876 58234
rect 19580 58180 19636 58182
rect 19660 58180 19716 58182
rect 19740 58180 19796 58182
rect 19820 58180 19876 58182
rect 19580 57146 19636 57148
rect 19660 57146 19716 57148
rect 19740 57146 19796 57148
rect 19820 57146 19876 57148
rect 19580 57094 19606 57146
rect 19606 57094 19636 57146
rect 19660 57094 19670 57146
rect 19670 57094 19716 57146
rect 19740 57094 19786 57146
rect 19786 57094 19796 57146
rect 19820 57094 19850 57146
rect 19850 57094 19876 57146
rect 19580 57092 19636 57094
rect 19660 57092 19716 57094
rect 19740 57092 19796 57094
rect 19820 57092 19876 57094
rect 19580 56058 19636 56060
rect 19660 56058 19716 56060
rect 19740 56058 19796 56060
rect 19820 56058 19876 56060
rect 19580 56006 19606 56058
rect 19606 56006 19636 56058
rect 19660 56006 19670 56058
rect 19670 56006 19716 56058
rect 19740 56006 19786 56058
rect 19786 56006 19796 56058
rect 19820 56006 19850 56058
rect 19850 56006 19876 56058
rect 19580 56004 19636 56006
rect 19660 56004 19716 56006
rect 19740 56004 19796 56006
rect 19820 56004 19876 56006
rect 19580 54970 19636 54972
rect 19660 54970 19716 54972
rect 19740 54970 19796 54972
rect 19820 54970 19876 54972
rect 19580 54918 19606 54970
rect 19606 54918 19636 54970
rect 19660 54918 19670 54970
rect 19670 54918 19716 54970
rect 19740 54918 19786 54970
rect 19786 54918 19796 54970
rect 19820 54918 19850 54970
rect 19850 54918 19876 54970
rect 19580 54916 19636 54918
rect 19660 54916 19716 54918
rect 19740 54916 19796 54918
rect 19820 54916 19876 54918
rect 19580 53882 19636 53884
rect 19660 53882 19716 53884
rect 19740 53882 19796 53884
rect 19820 53882 19876 53884
rect 19580 53830 19606 53882
rect 19606 53830 19636 53882
rect 19660 53830 19670 53882
rect 19670 53830 19716 53882
rect 19740 53830 19786 53882
rect 19786 53830 19796 53882
rect 19820 53830 19850 53882
rect 19850 53830 19876 53882
rect 19580 53828 19636 53830
rect 19660 53828 19716 53830
rect 19740 53828 19796 53830
rect 19820 53828 19876 53830
rect 19580 52794 19636 52796
rect 19660 52794 19716 52796
rect 19740 52794 19796 52796
rect 19820 52794 19876 52796
rect 19580 52742 19606 52794
rect 19606 52742 19636 52794
rect 19660 52742 19670 52794
rect 19670 52742 19716 52794
rect 19740 52742 19786 52794
rect 19786 52742 19796 52794
rect 19820 52742 19850 52794
rect 19850 52742 19876 52794
rect 19580 52740 19636 52742
rect 19660 52740 19716 52742
rect 19740 52740 19796 52742
rect 19820 52740 19876 52742
rect 19580 51706 19636 51708
rect 19660 51706 19716 51708
rect 19740 51706 19796 51708
rect 19820 51706 19876 51708
rect 19580 51654 19606 51706
rect 19606 51654 19636 51706
rect 19660 51654 19670 51706
rect 19670 51654 19716 51706
rect 19740 51654 19786 51706
rect 19786 51654 19796 51706
rect 19820 51654 19850 51706
rect 19850 51654 19876 51706
rect 19580 51652 19636 51654
rect 19660 51652 19716 51654
rect 19740 51652 19796 51654
rect 19820 51652 19876 51654
rect 19580 50618 19636 50620
rect 19660 50618 19716 50620
rect 19740 50618 19796 50620
rect 19820 50618 19876 50620
rect 19580 50566 19606 50618
rect 19606 50566 19636 50618
rect 19660 50566 19670 50618
rect 19670 50566 19716 50618
rect 19740 50566 19786 50618
rect 19786 50566 19796 50618
rect 19820 50566 19850 50618
rect 19850 50566 19876 50618
rect 19580 50564 19636 50566
rect 19660 50564 19716 50566
rect 19740 50564 19796 50566
rect 19820 50564 19876 50566
rect 19580 49530 19636 49532
rect 19660 49530 19716 49532
rect 19740 49530 19796 49532
rect 19820 49530 19876 49532
rect 19580 49478 19606 49530
rect 19606 49478 19636 49530
rect 19660 49478 19670 49530
rect 19670 49478 19716 49530
rect 19740 49478 19786 49530
rect 19786 49478 19796 49530
rect 19820 49478 19850 49530
rect 19850 49478 19876 49530
rect 19580 49476 19636 49478
rect 19660 49476 19716 49478
rect 19740 49476 19796 49478
rect 19820 49476 19876 49478
rect 19580 48442 19636 48444
rect 19660 48442 19716 48444
rect 19740 48442 19796 48444
rect 19820 48442 19876 48444
rect 19580 48390 19606 48442
rect 19606 48390 19636 48442
rect 19660 48390 19670 48442
rect 19670 48390 19716 48442
rect 19740 48390 19786 48442
rect 19786 48390 19796 48442
rect 19820 48390 19850 48442
rect 19850 48390 19876 48442
rect 19580 48388 19636 48390
rect 19660 48388 19716 48390
rect 19740 48388 19796 48390
rect 19820 48388 19876 48390
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 25686 29028 25742 29064
rect 25686 29008 25688 29028
rect 25688 29008 25740 29028
rect 25740 29008 25742 29028
rect 26422 71032 26478 71088
rect 26698 71052 26754 71088
rect 26698 71032 26700 71052
rect 26700 71032 26752 71052
rect 26752 71032 26754 71052
rect 26514 29044 26516 29064
rect 26516 29044 26568 29064
rect 26568 29044 26570 29064
rect 26514 29008 26570 29044
rect 34940 96858 34996 96860
rect 35020 96858 35076 96860
rect 35100 96858 35156 96860
rect 35180 96858 35236 96860
rect 34940 96806 34966 96858
rect 34966 96806 34996 96858
rect 35020 96806 35030 96858
rect 35030 96806 35076 96858
rect 35100 96806 35146 96858
rect 35146 96806 35156 96858
rect 35180 96806 35210 96858
rect 35210 96806 35236 96858
rect 34940 96804 34996 96806
rect 35020 96804 35076 96806
rect 35100 96804 35156 96806
rect 35180 96804 35236 96806
rect 34940 95770 34996 95772
rect 35020 95770 35076 95772
rect 35100 95770 35156 95772
rect 35180 95770 35236 95772
rect 34940 95718 34966 95770
rect 34966 95718 34996 95770
rect 35020 95718 35030 95770
rect 35030 95718 35076 95770
rect 35100 95718 35146 95770
rect 35146 95718 35156 95770
rect 35180 95718 35210 95770
rect 35210 95718 35236 95770
rect 34940 95716 34996 95718
rect 35020 95716 35076 95718
rect 35100 95716 35156 95718
rect 35180 95716 35236 95718
rect 34940 94682 34996 94684
rect 35020 94682 35076 94684
rect 35100 94682 35156 94684
rect 35180 94682 35236 94684
rect 34940 94630 34966 94682
rect 34966 94630 34996 94682
rect 35020 94630 35030 94682
rect 35030 94630 35076 94682
rect 35100 94630 35146 94682
rect 35146 94630 35156 94682
rect 35180 94630 35210 94682
rect 35210 94630 35236 94682
rect 34940 94628 34996 94630
rect 35020 94628 35076 94630
rect 35100 94628 35156 94630
rect 35180 94628 35236 94630
rect 34940 93594 34996 93596
rect 35020 93594 35076 93596
rect 35100 93594 35156 93596
rect 35180 93594 35236 93596
rect 34940 93542 34966 93594
rect 34966 93542 34996 93594
rect 35020 93542 35030 93594
rect 35030 93542 35076 93594
rect 35100 93542 35146 93594
rect 35146 93542 35156 93594
rect 35180 93542 35210 93594
rect 35210 93542 35236 93594
rect 34940 93540 34996 93542
rect 35020 93540 35076 93542
rect 35100 93540 35156 93542
rect 35180 93540 35236 93542
rect 34940 92506 34996 92508
rect 35020 92506 35076 92508
rect 35100 92506 35156 92508
rect 35180 92506 35236 92508
rect 34940 92454 34966 92506
rect 34966 92454 34996 92506
rect 35020 92454 35030 92506
rect 35030 92454 35076 92506
rect 35100 92454 35146 92506
rect 35146 92454 35156 92506
rect 35180 92454 35210 92506
rect 35210 92454 35236 92506
rect 34940 92452 34996 92454
rect 35020 92452 35076 92454
rect 35100 92452 35156 92454
rect 35180 92452 35236 92454
rect 34940 91418 34996 91420
rect 35020 91418 35076 91420
rect 35100 91418 35156 91420
rect 35180 91418 35236 91420
rect 34940 91366 34966 91418
rect 34966 91366 34996 91418
rect 35020 91366 35030 91418
rect 35030 91366 35076 91418
rect 35100 91366 35146 91418
rect 35146 91366 35156 91418
rect 35180 91366 35210 91418
rect 35210 91366 35236 91418
rect 34940 91364 34996 91366
rect 35020 91364 35076 91366
rect 35100 91364 35156 91366
rect 35180 91364 35236 91366
rect 34940 90330 34996 90332
rect 35020 90330 35076 90332
rect 35100 90330 35156 90332
rect 35180 90330 35236 90332
rect 34940 90278 34966 90330
rect 34966 90278 34996 90330
rect 35020 90278 35030 90330
rect 35030 90278 35076 90330
rect 35100 90278 35146 90330
rect 35146 90278 35156 90330
rect 35180 90278 35210 90330
rect 35210 90278 35236 90330
rect 34940 90276 34996 90278
rect 35020 90276 35076 90278
rect 35100 90276 35156 90278
rect 35180 90276 35236 90278
rect 34940 89242 34996 89244
rect 35020 89242 35076 89244
rect 35100 89242 35156 89244
rect 35180 89242 35236 89244
rect 34940 89190 34966 89242
rect 34966 89190 34996 89242
rect 35020 89190 35030 89242
rect 35030 89190 35076 89242
rect 35100 89190 35146 89242
rect 35146 89190 35156 89242
rect 35180 89190 35210 89242
rect 35210 89190 35236 89242
rect 34940 89188 34996 89190
rect 35020 89188 35076 89190
rect 35100 89188 35156 89190
rect 35180 89188 35236 89190
rect 34940 88154 34996 88156
rect 35020 88154 35076 88156
rect 35100 88154 35156 88156
rect 35180 88154 35236 88156
rect 34940 88102 34966 88154
rect 34966 88102 34996 88154
rect 35020 88102 35030 88154
rect 35030 88102 35076 88154
rect 35100 88102 35146 88154
rect 35146 88102 35156 88154
rect 35180 88102 35210 88154
rect 35210 88102 35236 88154
rect 34940 88100 34996 88102
rect 35020 88100 35076 88102
rect 35100 88100 35156 88102
rect 35180 88100 35236 88102
rect 34940 87066 34996 87068
rect 35020 87066 35076 87068
rect 35100 87066 35156 87068
rect 35180 87066 35236 87068
rect 34940 87014 34966 87066
rect 34966 87014 34996 87066
rect 35020 87014 35030 87066
rect 35030 87014 35076 87066
rect 35100 87014 35146 87066
rect 35146 87014 35156 87066
rect 35180 87014 35210 87066
rect 35210 87014 35236 87066
rect 34940 87012 34996 87014
rect 35020 87012 35076 87014
rect 35100 87012 35156 87014
rect 35180 87012 35236 87014
rect 34940 85978 34996 85980
rect 35020 85978 35076 85980
rect 35100 85978 35156 85980
rect 35180 85978 35236 85980
rect 34940 85926 34966 85978
rect 34966 85926 34996 85978
rect 35020 85926 35030 85978
rect 35030 85926 35076 85978
rect 35100 85926 35146 85978
rect 35146 85926 35156 85978
rect 35180 85926 35210 85978
rect 35210 85926 35236 85978
rect 34940 85924 34996 85926
rect 35020 85924 35076 85926
rect 35100 85924 35156 85926
rect 35180 85924 35236 85926
rect 34940 84890 34996 84892
rect 35020 84890 35076 84892
rect 35100 84890 35156 84892
rect 35180 84890 35236 84892
rect 34940 84838 34966 84890
rect 34966 84838 34996 84890
rect 35020 84838 35030 84890
rect 35030 84838 35076 84890
rect 35100 84838 35146 84890
rect 35146 84838 35156 84890
rect 35180 84838 35210 84890
rect 35210 84838 35236 84890
rect 34940 84836 34996 84838
rect 35020 84836 35076 84838
rect 35100 84836 35156 84838
rect 35180 84836 35236 84838
rect 34940 83802 34996 83804
rect 35020 83802 35076 83804
rect 35100 83802 35156 83804
rect 35180 83802 35236 83804
rect 34940 83750 34966 83802
rect 34966 83750 34996 83802
rect 35020 83750 35030 83802
rect 35030 83750 35076 83802
rect 35100 83750 35146 83802
rect 35146 83750 35156 83802
rect 35180 83750 35210 83802
rect 35210 83750 35236 83802
rect 34940 83748 34996 83750
rect 35020 83748 35076 83750
rect 35100 83748 35156 83750
rect 35180 83748 35236 83750
rect 34940 82714 34996 82716
rect 35020 82714 35076 82716
rect 35100 82714 35156 82716
rect 35180 82714 35236 82716
rect 34940 82662 34966 82714
rect 34966 82662 34996 82714
rect 35020 82662 35030 82714
rect 35030 82662 35076 82714
rect 35100 82662 35146 82714
rect 35146 82662 35156 82714
rect 35180 82662 35210 82714
rect 35210 82662 35236 82714
rect 34940 82660 34996 82662
rect 35020 82660 35076 82662
rect 35100 82660 35156 82662
rect 35180 82660 35236 82662
rect 34940 81626 34996 81628
rect 35020 81626 35076 81628
rect 35100 81626 35156 81628
rect 35180 81626 35236 81628
rect 34940 81574 34966 81626
rect 34966 81574 34996 81626
rect 35020 81574 35030 81626
rect 35030 81574 35076 81626
rect 35100 81574 35146 81626
rect 35146 81574 35156 81626
rect 35180 81574 35210 81626
rect 35210 81574 35236 81626
rect 34940 81572 34996 81574
rect 35020 81572 35076 81574
rect 35100 81572 35156 81574
rect 35180 81572 35236 81574
rect 34940 80538 34996 80540
rect 35020 80538 35076 80540
rect 35100 80538 35156 80540
rect 35180 80538 35236 80540
rect 34940 80486 34966 80538
rect 34966 80486 34996 80538
rect 35020 80486 35030 80538
rect 35030 80486 35076 80538
rect 35100 80486 35146 80538
rect 35146 80486 35156 80538
rect 35180 80486 35210 80538
rect 35210 80486 35236 80538
rect 34940 80484 34996 80486
rect 35020 80484 35076 80486
rect 35100 80484 35156 80486
rect 35180 80484 35236 80486
rect 34940 79450 34996 79452
rect 35020 79450 35076 79452
rect 35100 79450 35156 79452
rect 35180 79450 35236 79452
rect 34940 79398 34966 79450
rect 34966 79398 34996 79450
rect 35020 79398 35030 79450
rect 35030 79398 35076 79450
rect 35100 79398 35146 79450
rect 35146 79398 35156 79450
rect 35180 79398 35210 79450
rect 35210 79398 35236 79450
rect 34940 79396 34996 79398
rect 35020 79396 35076 79398
rect 35100 79396 35156 79398
rect 35180 79396 35236 79398
rect 34940 78362 34996 78364
rect 35020 78362 35076 78364
rect 35100 78362 35156 78364
rect 35180 78362 35236 78364
rect 34940 78310 34966 78362
rect 34966 78310 34996 78362
rect 35020 78310 35030 78362
rect 35030 78310 35076 78362
rect 35100 78310 35146 78362
rect 35146 78310 35156 78362
rect 35180 78310 35210 78362
rect 35210 78310 35236 78362
rect 34940 78308 34996 78310
rect 35020 78308 35076 78310
rect 35100 78308 35156 78310
rect 35180 78308 35236 78310
rect 34940 77274 34996 77276
rect 35020 77274 35076 77276
rect 35100 77274 35156 77276
rect 35180 77274 35236 77276
rect 34940 77222 34966 77274
rect 34966 77222 34996 77274
rect 35020 77222 35030 77274
rect 35030 77222 35076 77274
rect 35100 77222 35146 77274
rect 35146 77222 35156 77274
rect 35180 77222 35210 77274
rect 35210 77222 35236 77274
rect 34940 77220 34996 77222
rect 35020 77220 35076 77222
rect 35100 77220 35156 77222
rect 35180 77220 35236 77222
rect 34940 76186 34996 76188
rect 35020 76186 35076 76188
rect 35100 76186 35156 76188
rect 35180 76186 35236 76188
rect 34940 76134 34966 76186
rect 34966 76134 34996 76186
rect 35020 76134 35030 76186
rect 35030 76134 35076 76186
rect 35100 76134 35146 76186
rect 35146 76134 35156 76186
rect 35180 76134 35210 76186
rect 35210 76134 35236 76186
rect 34940 76132 34996 76134
rect 35020 76132 35076 76134
rect 35100 76132 35156 76134
rect 35180 76132 35236 76134
rect 34940 75098 34996 75100
rect 35020 75098 35076 75100
rect 35100 75098 35156 75100
rect 35180 75098 35236 75100
rect 34940 75046 34966 75098
rect 34966 75046 34996 75098
rect 35020 75046 35030 75098
rect 35030 75046 35076 75098
rect 35100 75046 35146 75098
rect 35146 75046 35156 75098
rect 35180 75046 35210 75098
rect 35210 75046 35236 75098
rect 34940 75044 34996 75046
rect 35020 75044 35076 75046
rect 35100 75044 35156 75046
rect 35180 75044 35236 75046
rect 34940 74010 34996 74012
rect 35020 74010 35076 74012
rect 35100 74010 35156 74012
rect 35180 74010 35236 74012
rect 34940 73958 34966 74010
rect 34966 73958 34996 74010
rect 35020 73958 35030 74010
rect 35030 73958 35076 74010
rect 35100 73958 35146 74010
rect 35146 73958 35156 74010
rect 35180 73958 35210 74010
rect 35210 73958 35236 74010
rect 34940 73956 34996 73958
rect 35020 73956 35076 73958
rect 35100 73956 35156 73958
rect 35180 73956 35236 73958
rect 34940 72922 34996 72924
rect 35020 72922 35076 72924
rect 35100 72922 35156 72924
rect 35180 72922 35236 72924
rect 34940 72870 34966 72922
rect 34966 72870 34996 72922
rect 35020 72870 35030 72922
rect 35030 72870 35076 72922
rect 35100 72870 35146 72922
rect 35146 72870 35156 72922
rect 35180 72870 35210 72922
rect 35210 72870 35236 72922
rect 34940 72868 34996 72870
rect 35020 72868 35076 72870
rect 35100 72868 35156 72870
rect 35180 72868 35236 72870
rect 34940 71834 34996 71836
rect 35020 71834 35076 71836
rect 35100 71834 35156 71836
rect 35180 71834 35236 71836
rect 34940 71782 34966 71834
rect 34966 71782 34996 71834
rect 35020 71782 35030 71834
rect 35030 71782 35076 71834
rect 35100 71782 35146 71834
rect 35146 71782 35156 71834
rect 35180 71782 35210 71834
rect 35210 71782 35236 71834
rect 34940 71780 34996 71782
rect 35020 71780 35076 71782
rect 35100 71780 35156 71782
rect 35180 71780 35236 71782
rect 34940 70746 34996 70748
rect 35020 70746 35076 70748
rect 35100 70746 35156 70748
rect 35180 70746 35236 70748
rect 34940 70694 34966 70746
rect 34966 70694 34996 70746
rect 35020 70694 35030 70746
rect 35030 70694 35076 70746
rect 35100 70694 35146 70746
rect 35146 70694 35156 70746
rect 35180 70694 35210 70746
rect 35210 70694 35236 70746
rect 34940 70692 34996 70694
rect 35020 70692 35076 70694
rect 35100 70692 35156 70694
rect 35180 70692 35236 70694
rect 34940 69658 34996 69660
rect 35020 69658 35076 69660
rect 35100 69658 35156 69660
rect 35180 69658 35236 69660
rect 34940 69606 34966 69658
rect 34966 69606 34996 69658
rect 35020 69606 35030 69658
rect 35030 69606 35076 69658
rect 35100 69606 35146 69658
rect 35146 69606 35156 69658
rect 35180 69606 35210 69658
rect 35210 69606 35236 69658
rect 34940 69604 34996 69606
rect 35020 69604 35076 69606
rect 35100 69604 35156 69606
rect 35180 69604 35236 69606
rect 34940 68570 34996 68572
rect 35020 68570 35076 68572
rect 35100 68570 35156 68572
rect 35180 68570 35236 68572
rect 34940 68518 34966 68570
rect 34966 68518 34996 68570
rect 35020 68518 35030 68570
rect 35030 68518 35076 68570
rect 35100 68518 35146 68570
rect 35146 68518 35156 68570
rect 35180 68518 35210 68570
rect 35210 68518 35236 68570
rect 34940 68516 34996 68518
rect 35020 68516 35076 68518
rect 35100 68516 35156 68518
rect 35180 68516 35236 68518
rect 34940 67482 34996 67484
rect 35020 67482 35076 67484
rect 35100 67482 35156 67484
rect 35180 67482 35236 67484
rect 34940 67430 34966 67482
rect 34966 67430 34996 67482
rect 35020 67430 35030 67482
rect 35030 67430 35076 67482
rect 35100 67430 35146 67482
rect 35146 67430 35156 67482
rect 35180 67430 35210 67482
rect 35210 67430 35236 67482
rect 34940 67428 34996 67430
rect 35020 67428 35076 67430
rect 35100 67428 35156 67430
rect 35180 67428 35236 67430
rect 34940 66394 34996 66396
rect 35020 66394 35076 66396
rect 35100 66394 35156 66396
rect 35180 66394 35236 66396
rect 34940 66342 34966 66394
rect 34966 66342 34996 66394
rect 35020 66342 35030 66394
rect 35030 66342 35076 66394
rect 35100 66342 35146 66394
rect 35146 66342 35156 66394
rect 35180 66342 35210 66394
rect 35210 66342 35236 66394
rect 34940 66340 34996 66342
rect 35020 66340 35076 66342
rect 35100 66340 35156 66342
rect 35180 66340 35236 66342
rect 34940 65306 34996 65308
rect 35020 65306 35076 65308
rect 35100 65306 35156 65308
rect 35180 65306 35236 65308
rect 34940 65254 34966 65306
rect 34966 65254 34996 65306
rect 35020 65254 35030 65306
rect 35030 65254 35076 65306
rect 35100 65254 35146 65306
rect 35146 65254 35156 65306
rect 35180 65254 35210 65306
rect 35210 65254 35236 65306
rect 34940 65252 34996 65254
rect 35020 65252 35076 65254
rect 35100 65252 35156 65254
rect 35180 65252 35236 65254
rect 34940 64218 34996 64220
rect 35020 64218 35076 64220
rect 35100 64218 35156 64220
rect 35180 64218 35236 64220
rect 34940 64166 34966 64218
rect 34966 64166 34996 64218
rect 35020 64166 35030 64218
rect 35030 64166 35076 64218
rect 35100 64166 35146 64218
rect 35146 64166 35156 64218
rect 35180 64166 35210 64218
rect 35210 64166 35236 64218
rect 34940 64164 34996 64166
rect 35020 64164 35076 64166
rect 35100 64164 35156 64166
rect 35180 64164 35236 64166
rect 34940 63130 34996 63132
rect 35020 63130 35076 63132
rect 35100 63130 35156 63132
rect 35180 63130 35236 63132
rect 34940 63078 34966 63130
rect 34966 63078 34996 63130
rect 35020 63078 35030 63130
rect 35030 63078 35076 63130
rect 35100 63078 35146 63130
rect 35146 63078 35156 63130
rect 35180 63078 35210 63130
rect 35210 63078 35236 63130
rect 34940 63076 34996 63078
rect 35020 63076 35076 63078
rect 35100 63076 35156 63078
rect 35180 63076 35236 63078
rect 34940 62042 34996 62044
rect 35020 62042 35076 62044
rect 35100 62042 35156 62044
rect 35180 62042 35236 62044
rect 34940 61990 34966 62042
rect 34966 61990 34996 62042
rect 35020 61990 35030 62042
rect 35030 61990 35076 62042
rect 35100 61990 35146 62042
rect 35146 61990 35156 62042
rect 35180 61990 35210 62042
rect 35210 61990 35236 62042
rect 34940 61988 34996 61990
rect 35020 61988 35076 61990
rect 35100 61988 35156 61990
rect 35180 61988 35236 61990
rect 34940 60954 34996 60956
rect 35020 60954 35076 60956
rect 35100 60954 35156 60956
rect 35180 60954 35236 60956
rect 34940 60902 34966 60954
rect 34966 60902 34996 60954
rect 35020 60902 35030 60954
rect 35030 60902 35076 60954
rect 35100 60902 35146 60954
rect 35146 60902 35156 60954
rect 35180 60902 35210 60954
rect 35210 60902 35236 60954
rect 34940 60900 34996 60902
rect 35020 60900 35076 60902
rect 35100 60900 35156 60902
rect 35180 60900 35236 60902
rect 34940 59866 34996 59868
rect 35020 59866 35076 59868
rect 35100 59866 35156 59868
rect 35180 59866 35236 59868
rect 34940 59814 34966 59866
rect 34966 59814 34996 59866
rect 35020 59814 35030 59866
rect 35030 59814 35076 59866
rect 35100 59814 35146 59866
rect 35146 59814 35156 59866
rect 35180 59814 35210 59866
rect 35210 59814 35236 59866
rect 34940 59812 34996 59814
rect 35020 59812 35076 59814
rect 35100 59812 35156 59814
rect 35180 59812 35236 59814
rect 34940 58778 34996 58780
rect 35020 58778 35076 58780
rect 35100 58778 35156 58780
rect 35180 58778 35236 58780
rect 34940 58726 34966 58778
rect 34966 58726 34996 58778
rect 35020 58726 35030 58778
rect 35030 58726 35076 58778
rect 35100 58726 35146 58778
rect 35146 58726 35156 58778
rect 35180 58726 35210 58778
rect 35210 58726 35236 58778
rect 34940 58724 34996 58726
rect 35020 58724 35076 58726
rect 35100 58724 35156 58726
rect 35180 58724 35236 58726
rect 34940 57690 34996 57692
rect 35020 57690 35076 57692
rect 35100 57690 35156 57692
rect 35180 57690 35236 57692
rect 34940 57638 34966 57690
rect 34966 57638 34996 57690
rect 35020 57638 35030 57690
rect 35030 57638 35076 57690
rect 35100 57638 35146 57690
rect 35146 57638 35156 57690
rect 35180 57638 35210 57690
rect 35210 57638 35236 57690
rect 34940 57636 34996 57638
rect 35020 57636 35076 57638
rect 35100 57636 35156 57638
rect 35180 57636 35236 57638
rect 34940 56602 34996 56604
rect 35020 56602 35076 56604
rect 35100 56602 35156 56604
rect 35180 56602 35236 56604
rect 34940 56550 34966 56602
rect 34966 56550 34996 56602
rect 35020 56550 35030 56602
rect 35030 56550 35076 56602
rect 35100 56550 35146 56602
rect 35146 56550 35156 56602
rect 35180 56550 35210 56602
rect 35210 56550 35236 56602
rect 34940 56548 34996 56550
rect 35020 56548 35076 56550
rect 35100 56548 35156 56550
rect 35180 56548 35236 56550
rect 34940 55514 34996 55516
rect 35020 55514 35076 55516
rect 35100 55514 35156 55516
rect 35180 55514 35236 55516
rect 34940 55462 34966 55514
rect 34966 55462 34996 55514
rect 35020 55462 35030 55514
rect 35030 55462 35076 55514
rect 35100 55462 35146 55514
rect 35146 55462 35156 55514
rect 35180 55462 35210 55514
rect 35210 55462 35236 55514
rect 34940 55460 34996 55462
rect 35020 55460 35076 55462
rect 35100 55460 35156 55462
rect 35180 55460 35236 55462
rect 34940 54426 34996 54428
rect 35020 54426 35076 54428
rect 35100 54426 35156 54428
rect 35180 54426 35236 54428
rect 34940 54374 34966 54426
rect 34966 54374 34996 54426
rect 35020 54374 35030 54426
rect 35030 54374 35076 54426
rect 35100 54374 35146 54426
rect 35146 54374 35156 54426
rect 35180 54374 35210 54426
rect 35210 54374 35236 54426
rect 34940 54372 34996 54374
rect 35020 54372 35076 54374
rect 35100 54372 35156 54374
rect 35180 54372 35236 54374
rect 34940 53338 34996 53340
rect 35020 53338 35076 53340
rect 35100 53338 35156 53340
rect 35180 53338 35236 53340
rect 34940 53286 34966 53338
rect 34966 53286 34996 53338
rect 35020 53286 35030 53338
rect 35030 53286 35076 53338
rect 35100 53286 35146 53338
rect 35146 53286 35156 53338
rect 35180 53286 35210 53338
rect 35210 53286 35236 53338
rect 34940 53284 34996 53286
rect 35020 53284 35076 53286
rect 35100 53284 35156 53286
rect 35180 53284 35236 53286
rect 34940 52250 34996 52252
rect 35020 52250 35076 52252
rect 35100 52250 35156 52252
rect 35180 52250 35236 52252
rect 34940 52198 34966 52250
rect 34966 52198 34996 52250
rect 35020 52198 35030 52250
rect 35030 52198 35076 52250
rect 35100 52198 35146 52250
rect 35146 52198 35156 52250
rect 35180 52198 35210 52250
rect 35210 52198 35236 52250
rect 34940 52196 34996 52198
rect 35020 52196 35076 52198
rect 35100 52196 35156 52198
rect 35180 52196 35236 52198
rect 34940 51162 34996 51164
rect 35020 51162 35076 51164
rect 35100 51162 35156 51164
rect 35180 51162 35236 51164
rect 34940 51110 34966 51162
rect 34966 51110 34996 51162
rect 35020 51110 35030 51162
rect 35030 51110 35076 51162
rect 35100 51110 35146 51162
rect 35146 51110 35156 51162
rect 35180 51110 35210 51162
rect 35210 51110 35236 51162
rect 34940 51108 34996 51110
rect 35020 51108 35076 51110
rect 35100 51108 35156 51110
rect 35180 51108 35236 51110
rect 34940 50074 34996 50076
rect 35020 50074 35076 50076
rect 35100 50074 35156 50076
rect 35180 50074 35236 50076
rect 34940 50022 34966 50074
rect 34966 50022 34996 50074
rect 35020 50022 35030 50074
rect 35030 50022 35076 50074
rect 35100 50022 35146 50074
rect 35146 50022 35156 50074
rect 35180 50022 35210 50074
rect 35210 50022 35236 50074
rect 34940 50020 34996 50022
rect 35020 50020 35076 50022
rect 35100 50020 35156 50022
rect 35180 50020 35236 50022
rect 34940 48986 34996 48988
rect 35020 48986 35076 48988
rect 35100 48986 35156 48988
rect 35180 48986 35236 48988
rect 34940 48934 34966 48986
rect 34966 48934 34996 48986
rect 35020 48934 35030 48986
rect 35030 48934 35076 48986
rect 35100 48934 35146 48986
rect 35146 48934 35156 48986
rect 35180 48934 35210 48986
rect 35210 48934 35236 48986
rect 34940 48932 34996 48934
rect 35020 48932 35076 48934
rect 35100 48932 35156 48934
rect 35180 48932 35236 48934
rect 34940 47898 34996 47900
rect 35020 47898 35076 47900
rect 35100 47898 35156 47900
rect 35180 47898 35236 47900
rect 34940 47846 34966 47898
rect 34966 47846 34996 47898
rect 35020 47846 35030 47898
rect 35030 47846 35076 47898
rect 35100 47846 35146 47898
rect 35146 47846 35156 47898
rect 35180 47846 35210 47898
rect 35210 47846 35236 47898
rect 34940 47844 34996 47846
rect 35020 47844 35076 47846
rect 35100 47844 35156 47846
rect 35180 47844 35236 47846
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 42614 79600 42670 79656
rect 43074 21972 43076 21992
rect 43076 21972 43128 21992
rect 43128 21972 43130 21992
rect 43074 21936 43130 21972
rect 43442 79600 43498 79656
rect 44454 19488 44510 19544
rect 44546 19388 44548 19408
rect 44548 19388 44600 19408
rect 44600 19388 44602 19408
rect 44546 19352 44602 19388
rect 45098 19488 45154 19544
rect 44546 14340 44602 14376
rect 44546 14320 44548 14340
rect 44548 14320 44600 14340
rect 44600 14320 44602 14340
rect 45374 19372 45430 19408
rect 45374 19352 45376 19372
rect 45376 19352 45428 19372
rect 45428 19352 45430 19372
rect 45374 14340 45430 14376
rect 45374 14320 45376 14340
rect 45376 14320 45428 14340
rect 45428 14320 45430 14340
rect 47950 21936 48006 21992
rect 50300 97402 50356 97404
rect 50380 97402 50436 97404
rect 50460 97402 50516 97404
rect 50540 97402 50596 97404
rect 50300 97350 50326 97402
rect 50326 97350 50356 97402
rect 50380 97350 50390 97402
rect 50390 97350 50436 97402
rect 50460 97350 50506 97402
rect 50506 97350 50516 97402
rect 50540 97350 50570 97402
rect 50570 97350 50596 97402
rect 50300 97348 50356 97350
rect 50380 97348 50436 97350
rect 50460 97348 50516 97350
rect 50540 97348 50596 97350
rect 50300 96314 50356 96316
rect 50380 96314 50436 96316
rect 50460 96314 50516 96316
rect 50540 96314 50596 96316
rect 50300 96262 50326 96314
rect 50326 96262 50356 96314
rect 50380 96262 50390 96314
rect 50390 96262 50436 96314
rect 50460 96262 50506 96314
rect 50506 96262 50516 96314
rect 50540 96262 50570 96314
rect 50570 96262 50596 96314
rect 50300 96260 50356 96262
rect 50380 96260 50436 96262
rect 50460 96260 50516 96262
rect 50540 96260 50596 96262
rect 50300 95226 50356 95228
rect 50380 95226 50436 95228
rect 50460 95226 50516 95228
rect 50540 95226 50596 95228
rect 50300 95174 50326 95226
rect 50326 95174 50356 95226
rect 50380 95174 50390 95226
rect 50390 95174 50436 95226
rect 50460 95174 50506 95226
rect 50506 95174 50516 95226
rect 50540 95174 50570 95226
rect 50570 95174 50596 95226
rect 50300 95172 50356 95174
rect 50380 95172 50436 95174
rect 50460 95172 50516 95174
rect 50540 95172 50596 95174
rect 50300 94138 50356 94140
rect 50380 94138 50436 94140
rect 50460 94138 50516 94140
rect 50540 94138 50596 94140
rect 50300 94086 50326 94138
rect 50326 94086 50356 94138
rect 50380 94086 50390 94138
rect 50390 94086 50436 94138
rect 50460 94086 50506 94138
rect 50506 94086 50516 94138
rect 50540 94086 50570 94138
rect 50570 94086 50596 94138
rect 50300 94084 50356 94086
rect 50380 94084 50436 94086
rect 50460 94084 50516 94086
rect 50540 94084 50596 94086
rect 49422 64524 49478 64560
rect 49422 64504 49424 64524
rect 49424 64504 49476 64524
rect 49476 64504 49478 64524
rect 50300 93050 50356 93052
rect 50380 93050 50436 93052
rect 50460 93050 50516 93052
rect 50540 93050 50596 93052
rect 50300 92998 50326 93050
rect 50326 92998 50356 93050
rect 50380 92998 50390 93050
rect 50390 92998 50436 93050
rect 50460 92998 50506 93050
rect 50506 92998 50516 93050
rect 50540 92998 50570 93050
rect 50570 92998 50596 93050
rect 50300 92996 50356 92998
rect 50380 92996 50436 92998
rect 50460 92996 50516 92998
rect 50540 92996 50596 92998
rect 50300 91962 50356 91964
rect 50380 91962 50436 91964
rect 50460 91962 50516 91964
rect 50540 91962 50596 91964
rect 50300 91910 50326 91962
rect 50326 91910 50356 91962
rect 50380 91910 50390 91962
rect 50390 91910 50436 91962
rect 50460 91910 50506 91962
rect 50506 91910 50516 91962
rect 50540 91910 50570 91962
rect 50570 91910 50596 91962
rect 50300 91908 50356 91910
rect 50380 91908 50436 91910
rect 50460 91908 50516 91910
rect 50540 91908 50596 91910
rect 50300 90874 50356 90876
rect 50380 90874 50436 90876
rect 50460 90874 50516 90876
rect 50540 90874 50596 90876
rect 50300 90822 50326 90874
rect 50326 90822 50356 90874
rect 50380 90822 50390 90874
rect 50390 90822 50436 90874
rect 50460 90822 50506 90874
rect 50506 90822 50516 90874
rect 50540 90822 50570 90874
rect 50570 90822 50596 90874
rect 50300 90820 50356 90822
rect 50380 90820 50436 90822
rect 50460 90820 50516 90822
rect 50540 90820 50596 90822
rect 50300 89786 50356 89788
rect 50380 89786 50436 89788
rect 50460 89786 50516 89788
rect 50540 89786 50596 89788
rect 50300 89734 50326 89786
rect 50326 89734 50356 89786
rect 50380 89734 50390 89786
rect 50390 89734 50436 89786
rect 50460 89734 50506 89786
rect 50506 89734 50516 89786
rect 50540 89734 50570 89786
rect 50570 89734 50596 89786
rect 50300 89732 50356 89734
rect 50380 89732 50436 89734
rect 50460 89732 50516 89734
rect 50540 89732 50596 89734
rect 50300 88698 50356 88700
rect 50380 88698 50436 88700
rect 50460 88698 50516 88700
rect 50540 88698 50596 88700
rect 50300 88646 50326 88698
rect 50326 88646 50356 88698
rect 50380 88646 50390 88698
rect 50390 88646 50436 88698
rect 50460 88646 50506 88698
rect 50506 88646 50516 88698
rect 50540 88646 50570 88698
rect 50570 88646 50596 88698
rect 50300 88644 50356 88646
rect 50380 88644 50436 88646
rect 50460 88644 50516 88646
rect 50540 88644 50596 88646
rect 50300 87610 50356 87612
rect 50380 87610 50436 87612
rect 50460 87610 50516 87612
rect 50540 87610 50596 87612
rect 50300 87558 50326 87610
rect 50326 87558 50356 87610
rect 50380 87558 50390 87610
rect 50390 87558 50436 87610
rect 50460 87558 50506 87610
rect 50506 87558 50516 87610
rect 50540 87558 50570 87610
rect 50570 87558 50596 87610
rect 50300 87556 50356 87558
rect 50380 87556 50436 87558
rect 50460 87556 50516 87558
rect 50540 87556 50596 87558
rect 50300 86522 50356 86524
rect 50380 86522 50436 86524
rect 50460 86522 50516 86524
rect 50540 86522 50596 86524
rect 50300 86470 50326 86522
rect 50326 86470 50356 86522
rect 50380 86470 50390 86522
rect 50390 86470 50436 86522
rect 50460 86470 50506 86522
rect 50506 86470 50516 86522
rect 50540 86470 50570 86522
rect 50570 86470 50596 86522
rect 50300 86468 50356 86470
rect 50380 86468 50436 86470
rect 50460 86468 50516 86470
rect 50540 86468 50596 86470
rect 50300 85434 50356 85436
rect 50380 85434 50436 85436
rect 50460 85434 50516 85436
rect 50540 85434 50596 85436
rect 50300 85382 50326 85434
rect 50326 85382 50356 85434
rect 50380 85382 50390 85434
rect 50390 85382 50436 85434
rect 50460 85382 50506 85434
rect 50506 85382 50516 85434
rect 50540 85382 50570 85434
rect 50570 85382 50596 85434
rect 50300 85380 50356 85382
rect 50380 85380 50436 85382
rect 50460 85380 50516 85382
rect 50540 85380 50596 85382
rect 50300 84346 50356 84348
rect 50380 84346 50436 84348
rect 50460 84346 50516 84348
rect 50540 84346 50596 84348
rect 50300 84294 50326 84346
rect 50326 84294 50356 84346
rect 50380 84294 50390 84346
rect 50390 84294 50436 84346
rect 50460 84294 50506 84346
rect 50506 84294 50516 84346
rect 50540 84294 50570 84346
rect 50570 84294 50596 84346
rect 50300 84292 50356 84294
rect 50380 84292 50436 84294
rect 50460 84292 50516 84294
rect 50540 84292 50596 84294
rect 50300 83258 50356 83260
rect 50380 83258 50436 83260
rect 50460 83258 50516 83260
rect 50540 83258 50596 83260
rect 50300 83206 50326 83258
rect 50326 83206 50356 83258
rect 50380 83206 50390 83258
rect 50390 83206 50436 83258
rect 50460 83206 50506 83258
rect 50506 83206 50516 83258
rect 50540 83206 50570 83258
rect 50570 83206 50596 83258
rect 50300 83204 50356 83206
rect 50380 83204 50436 83206
rect 50460 83204 50516 83206
rect 50540 83204 50596 83206
rect 50300 82170 50356 82172
rect 50380 82170 50436 82172
rect 50460 82170 50516 82172
rect 50540 82170 50596 82172
rect 50300 82118 50326 82170
rect 50326 82118 50356 82170
rect 50380 82118 50390 82170
rect 50390 82118 50436 82170
rect 50460 82118 50506 82170
rect 50506 82118 50516 82170
rect 50540 82118 50570 82170
rect 50570 82118 50596 82170
rect 50300 82116 50356 82118
rect 50380 82116 50436 82118
rect 50460 82116 50516 82118
rect 50540 82116 50596 82118
rect 50300 81082 50356 81084
rect 50380 81082 50436 81084
rect 50460 81082 50516 81084
rect 50540 81082 50596 81084
rect 50300 81030 50326 81082
rect 50326 81030 50356 81082
rect 50380 81030 50390 81082
rect 50390 81030 50436 81082
rect 50460 81030 50506 81082
rect 50506 81030 50516 81082
rect 50540 81030 50570 81082
rect 50570 81030 50596 81082
rect 50300 81028 50356 81030
rect 50380 81028 50436 81030
rect 50460 81028 50516 81030
rect 50540 81028 50596 81030
rect 50300 79994 50356 79996
rect 50380 79994 50436 79996
rect 50460 79994 50516 79996
rect 50540 79994 50596 79996
rect 50300 79942 50326 79994
rect 50326 79942 50356 79994
rect 50380 79942 50390 79994
rect 50390 79942 50436 79994
rect 50460 79942 50506 79994
rect 50506 79942 50516 79994
rect 50540 79942 50570 79994
rect 50570 79942 50596 79994
rect 50300 79940 50356 79942
rect 50380 79940 50436 79942
rect 50460 79940 50516 79942
rect 50540 79940 50596 79942
rect 50300 78906 50356 78908
rect 50380 78906 50436 78908
rect 50460 78906 50516 78908
rect 50540 78906 50596 78908
rect 50300 78854 50326 78906
rect 50326 78854 50356 78906
rect 50380 78854 50390 78906
rect 50390 78854 50436 78906
rect 50460 78854 50506 78906
rect 50506 78854 50516 78906
rect 50540 78854 50570 78906
rect 50570 78854 50596 78906
rect 50300 78852 50356 78854
rect 50380 78852 50436 78854
rect 50460 78852 50516 78854
rect 50540 78852 50596 78854
rect 50300 77818 50356 77820
rect 50380 77818 50436 77820
rect 50460 77818 50516 77820
rect 50540 77818 50596 77820
rect 50300 77766 50326 77818
rect 50326 77766 50356 77818
rect 50380 77766 50390 77818
rect 50390 77766 50436 77818
rect 50460 77766 50506 77818
rect 50506 77766 50516 77818
rect 50540 77766 50570 77818
rect 50570 77766 50596 77818
rect 50300 77764 50356 77766
rect 50380 77764 50436 77766
rect 50460 77764 50516 77766
rect 50540 77764 50596 77766
rect 50300 76730 50356 76732
rect 50380 76730 50436 76732
rect 50460 76730 50516 76732
rect 50540 76730 50596 76732
rect 50300 76678 50326 76730
rect 50326 76678 50356 76730
rect 50380 76678 50390 76730
rect 50390 76678 50436 76730
rect 50460 76678 50506 76730
rect 50506 76678 50516 76730
rect 50540 76678 50570 76730
rect 50570 76678 50596 76730
rect 50300 76676 50356 76678
rect 50380 76676 50436 76678
rect 50460 76676 50516 76678
rect 50540 76676 50596 76678
rect 50300 75642 50356 75644
rect 50380 75642 50436 75644
rect 50460 75642 50516 75644
rect 50540 75642 50596 75644
rect 50300 75590 50326 75642
rect 50326 75590 50356 75642
rect 50380 75590 50390 75642
rect 50390 75590 50436 75642
rect 50460 75590 50506 75642
rect 50506 75590 50516 75642
rect 50540 75590 50570 75642
rect 50570 75590 50596 75642
rect 50300 75588 50356 75590
rect 50380 75588 50436 75590
rect 50460 75588 50516 75590
rect 50540 75588 50596 75590
rect 50300 74554 50356 74556
rect 50380 74554 50436 74556
rect 50460 74554 50516 74556
rect 50540 74554 50596 74556
rect 50300 74502 50326 74554
rect 50326 74502 50356 74554
rect 50380 74502 50390 74554
rect 50390 74502 50436 74554
rect 50460 74502 50506 74554
rect 50506 74502 50516 74554
rect 50540 74502 50570 74554
rect 50570 74502 50596 74554
rect 50300 74500 50356 74502
rect 50380 74500 50436 74502
rect 50460 74500 50516 74502
rect 50540 74500 50596 74502
rect 50300 73466 50356 73468
rect 50380 73466 50436 73468
rect 50460 73466 50516 73468
rect 50540 73466 50596 73468
rect 50300 73414 50326 73466
rect 50326 73414 50356 73466
rect 50380 73414 50390 73466
rect 50390 73414 50436 73466
rect 50460 73414 50506 73466
rect 50506 73414 50516 73466
rect 50540 73414 50570 73466
rect 50570 73414 50596 73466
rect 50300 73412 50356 73414
rect 50380 73412 50436 73414
rect 50460 73412 50516 73414
rect 50540 73412 50596 73414
rect 50300 72378 50356 72380
rect 50380 72378 50436 72380
rect 50460 72378 50516 72380
rect 50540 72378 50596 72380
rect 50300 72326 50326 72378
rect 50326 72326 50356 72378
rect 50380 72326 50390 72378
rect 50390 72326 50436 72378
rect 50460 72326 50506 72378
rect 50506 72326 50516 72378
rect 50540 72326 50570 72378
rect 50570 72326 50596 72378
rect 50300 72324 50356 72326
rect 50380 72324 50436 72326
rect 50460 72324 50516 72326
rect 50540 72324 50596 72326
rect 50300 71290 50356 71292
rect 50380 71290 50436 71292
rect 50460 71290 50516 71292
rect 50540 71290 50596 71292
rect 50300 71238 50326 71290
rect 50326 71238 50356 71290
rect 50380 71238 50390 71290
rect 50390 71238 50436 71290
rect 50460 71238 50506 71290
rect 50506 71238 50516 71290
rect 50540 71238 50570 71290
rect 50570 71238 50596 71290
rect 50300 71236 50356 71238
rect 50380 71236 50436 71238
rect 50460 71236 50516 71238
rect 50540 71236 50596 71238
rect 50300 70202 50356 70204
rect 50380 70202 50436 70204
rect 50460 70202 50516 70204
rect 50540 70202 50596 70204
rect 50300 70150 50326 70202
rect 50326 70150 50356 70202
rect 50380 70150 50390 70202
rect 50390 70150 50436 70202
rect 50460 70150 50506 70202
rect 50506 70150 50516 70202
rect 50540 70150 50570 70202
rect 50570 70150 50596 70202
rect 50300 70148 50356 70150
rect 50380 70148 50436 70150
rect 50460 70148 50516 70150
rect 50540 70148 50596 70150
rect 49882 64388 49938 64424
rect 49882 64368 49884 64388
rect 49884 64368 49936 64388
rect 49936 64368 49938 64388
rect 50300 69114 50356 69116
rect 50380 69114 50436 69116
rect 50460 69114 50516 69116
rect 50540 69114 50596 69116
rect 50300 69062 50326 69114
rect 50326 69062 50356 69114
rect 50380 69062 50390 69114
rect 50390 69062 50436 69114
rect 50460 69062 50506 69114
rect 50506 69062 50516 69114
rect 50540 69062 50570 69114
rect 50570 69062 50596 69114
rect 50300 69060 50356 69062
rect 50380 69060 50436 69062
rect 50460 69060 50516 69062
rect 50540 69060 50596 69062
rect 50300 68026 50356 68028
rect 50380 68026 50436 68028
rect 50460 68026 50516 68028
rect 50540 68026 50596 68028
rect 50300 67974 50326 68026
rect 50326 67974 50356 68026
rect 50380 67974 50390 68026
rect 50390 67974 50436 68026
rect 50460 67974 50506 68026
rect 50506 67974 50516 68026
rect 50540 67974 50570 68026
rect 50570 67974 50596 68026
rect 50300 67972 50356 67974
rect 50380 67972 50436 67974
rect 50460 67972 50516 67974
rect 50540 67972 50596 67974
rect 50300 66938 50356 66940
rect 50380 66938 50436 66940
rect 50460 66938 50516 66940
rect 50540 66938 50596 66940
rect 50300 66886 50326 66938
rect 50326 66886 50356 66938
rect 50380 66886 50390 66938
rect 50390 66886 50436 66938
rect 50460 66886 50506 66938
rect 50506 66886 50516 66938
rect 50540 66886 50570 66938
rect 50570 66886 50596 66938
rect 50300 66884 50356 66886
rect 50380 66884 50436 66886
rect 50460 66884 50516 66886
rect 50540 66884 50596 66886
rect 50300 65850 50356 65852
rect 50380 65850 50436 65852
rect 50460 65850 50516 65852
rect 50540 65850 50596 65852
rect 50300 65798 50326 65850
rect 50326 65798 50356 65850
rect 50380 65798 50390 65850
rect 50390 65798 50436 65850
rect 50460 65798 50506 65850
rect 50506 65798 50516 65850
rect 50540 65798 50570 65850
rect 50570 65798 50596 65850
rect 50300 65796 50356 65798
rect 50380 65796 50436 65798
rect 50460 65796 50516 65798
rect 50540 65796 50596 65798
rect 50300 64762 50356 64764
rect 50380 64762 50436 64764
rect 50460 64762 50516 64764
rect 50540 64762 50596 64764
rect 50300 64710 50326 64762
rect 50326 64710 50356 64762
rect 50380 64710 50390 64762
rect 50390 64710 50436 64762
rect 50460 64710 50506 64762
rect 50506 64710 50516 64762
rect 50540 64710 50570 64762
rect 50570 64710 50596 64762
rect 50300 64708 50356 64710
rect 50380 64708 50436 64710
rect 50460 64708 50516 64710
rect 50540 64708 50596 64710
rect 50342 64540 50344 64560
rect 50344 64540 50396 64560
rect 50396 64540 50398 64560
rect 50342 64504 50398 64540
rect 50250 64388 50306 64424
rect 50250 64368 50252 64388
rect 50252 64368 50304 64388
rect 50304 64368 50306 64388
rect 50300 63674 50356 63676
rect 50380 63674 50436 63676
rect 50460 63674 50516 63676
rect 50540 63674 50596 63676
rect 50300 63622 50326 63674
rect 50326 63622 50356 63674
rect 50380 63622 50390 63674
rect 50390 63622 50436 63674
rect 50460 63622 50506 63674
rect 50506 63622 50516 63674
rect 50540 63622 50570 63674
rect 50570 63622 50596 63674
rect 50300 63620 50356 63622
rect 50380 63620 50436 63622
rect 50460 63620 50516 63622
rect 50540 63620 50596 63622
rect 50300 62586 50356 62588
rect 50380 62586 50436 62588
rect 50460 62586 50516 62588
rect 50540 62586 50596 62588
rect 50300 62534 50326 62586
rect 50326 62534 50356 62586
rect 50380 62534 50390 62586
rect 50390 62534 50436 62586
rect 50460 62534 50506 62586
rect 50506 62534 50516 62586
rect 50540 62534 50570 62586
rect 50570 62534 50596 62586
rect 50300 62532 50356 62534
rect 50380 62532 50436 62534
rect 50460 62532 50516 62534
rect 50540 62532 50596 62534
rect 50300 61498 50356 61500
rect 50380 61498 50436 61500
rect 50460 61498 50516 61500
rect 50540 61498 50596 61500
rect 50300 61446 50326 61498
rect 50326 61446 50356 61498
rect 50380 61446 50390 61498
rect 50390 61446 50436 61498
rect 50460 61446 50506 61498
rect 50506 61446 50516 61498
rect 50540 61446 50570 61498
rect 50570 61446 50596 61498
rect 50300 61444 50356 61446
rect 50380 61444 50436 61446
rect 50460 61444 50516 61446
rect 50540 61444 50596 61446
rect 50300 60410 50356 60412
rect 50380 60410 50436 60412
rect 50460 60410 50516 60412
rect 50540 60410 50596 60412
rect 50300 60358 50326 60410
rect 50326 60358 50356 60410
rect 50380 60358 50390 60410
rect 50390 60358 50436 60410
rect 50460 60358 50506 60410
rect 50506 60358 50516 60410
rect 50540 60358 50570 60410
rect 50570 60358 50596 60410
rect 50300 60356 50356 60358
rect 50380 60356 50436 60358
rect 50460 60356 50516 60358
rect 50540 60356 50596 60358
rect 50300 59322 50356 59324
rect 50380 59322 50436 59324
rect 50460 59322 50516 59324
rect 50540 59322 50596 59324
rect 50300 59270 50326 59322
rect 50326 59270 50356 59322
rect 50380 59270 50390 59322
rect 50390 59270 50436 59322
rect 50460 59270 50506 59322
rect 50506 59270 50516 59322
rect 50540 59270 50570 59322
rect 50570 59270 50596 59322
rect 50300 59268 50356 59270
rect 50380 59268 50436 59270
rect 50460 59268 50516 59270
rect 50540 59268 50596 59270
rect 50300 58234 50356 58236
rect 50380 58234 50436 58236
rect 50460 58234 50516 58236
rect 50540 58234 50596 58236
rect 50300 58182 50326 58234
rect 50326 58182 50356 58234
rect 50380 58182 50390 58234
rect 50390 58182 50436 58234
rect 50460 58182 50506 58234
rect 50506 58182 50516 58234
rect 50540 58182 50570 58234
rect 50570 58182 50596 58234
rect 50300 58180 50356 58182
rect 50380 58180 50436 58182
rect 50460 58180 50516 58182
rect 50540 58180 50596 58182
rect 50300 57146 50356 57148
rect 50380 57146 50436 57148
rect 50460 57146 50516 57148
rect 50540 57146 50596 57148
rect 50300 57094 50326 57146
rect 50326 57094 50356 57146
rect 50380 57094 50390 57146
rect 50390 57094 50436 57146
rect 50460 57094 50506 57146
rect 50506 57094 50516 57146
rect 50540 57094 50570 57146
rect 50570 57094 50596 57146
rect 50300 57092 50356 57094
rect 50380 57092 50436 57094
rect 50460 57092 50516 57094
rect 50540 57092 50596 57094
rect 50300 56058 50356 56060
rect 50380 56058 50436 56060
rect 50460 56058 50516 56060
rect 50540 56058 50596 56060
rect 50300 56006 50326 56058
rect 50326 56006 50356 56058
rect 50380 56006 50390 56058
rect 50390 56006 50436 56058
rect 50460 56006 50506 56058
rect 50506 56006 50516 56058
rect 50540 56006 50570 56058
rect 50570 56006 50596 56058
rect 50300 56004 50356 56006
rect 50380 56004 50436 56006
rect 50460 56004 50516 56006
rect 50540 56004 50596 56006
rect 50300 54970 50356 54972
rect 50380 54970 50436 54972
rect 50460 54970 50516 54972
rect 50540 54970 50596 54972
rect 50300 54918 50326 54970
rect 50326 54918 50356 54970
rect 50380 54918 50390 54970
rect 50390 54918 50436 54970
rect 50460 54918 50506 54970
rect 50506 54918 50516 54970
rect 50540 54918 50570 54970
rect 50570 54918 50596 54970
rect 50300 54916 50356 54918
rect 50380 54916 50436 54918
rect 50460 54916 50516 54918
rect 50540 54916 50596 54918
rect 50300 53882 50356 53884
rect 50380 53882 50436 53884
rect 50460 53882 50516 53884
rect 50540 53882 50596 53884
rect 50300 53830 50326 53882
rect 50326 53830 50356 53882
rect 50380 53830 50390 53882
rect 50390 53830 50436 53882
rect 50460 53830 50506 53882
rect 50506 53830 50516 53882
rect 50540 53830 50570 53882
rect 50570 53830 50596 53882
rect 50300 53828 50356 53830
rect 50380 53828 50436 53830
rect 50460 53828 50516 53830
rect 50540 53828 50596 53830
rect 50300 52794 50356 52796
rect 50380 52794 50436 52796
rect 50460 52794 50516 52796
rect 50540 52794 50596 52796
rect 50300 52742 50326 52794
rect 50326 52742 50356 52794
rect 50380 52742 50390 52794
rect 50390 52742 50436 52794
rect 50460 52742 50506 52794
rect 50506 52742 50516 52794
rect 50540 52742 50570 52794
rect 50570 52742 50596 52794
rect 50300 52740 50356 52742
rect 50380 52740 50436 52742
rect 50460 52740 50516 52742
rect 50540 52740 50596 52742
rect 50300 51706 50356 51708
rect 50380 51706 50436 51708
rect 50460 51706 50516 51708
rect 50540 51706 50596 51708
rect 50300 51654 50326 51706
rect 50326 51654 50356 51706
rect 50380 51654 50390 51706
rect 50390 51654 50436 51706
rect 50460 51654 50506 51706
rect 50506 51654 50516 51706
rect 50540 51654 50570 51706
rect 50570 51654 50596 51706
rect 50300 51652 50356 51654
rect 50380 51652 50436 51654
rect 50460 51652 50516 51654
rect 50540 51652 50596 51654
rect 50300 50618 50356 50620
rect 50380 50618 50436 50620
rect 50460 50618 50516 50620
rect 50540 50618 50596 50620
rect 50300 50566 50326 50618
rect 50326 50566 50356 50618
rect 50380 50566 50390 50618
rect 50390 50566 50436 50618
rect 50460 50566 50506 50618
rect 50506 50566 50516 50618
rect 50540 50566 50570 50618
rect 50570 50566 50596 50618
rect 50300 50564 50356 50566
rect 50380 50564 50436 50566
rect 50460 50564 50516 50566
rect 50540 50564 50596 50566
rect 50300 49530 50356 49532
rect 50380 49530 50436 49532
rect 50460 49530 50516 49532
rect 50540 49530 50596 49532
rect 50300 49478 50326 49530
rect 50326 49478 50356 49530
rect 50380 49478 50390 49530
rect 50390 49478 50436 49530
rect 50460 49478 50506 49530
rect 50506 49478 50516 49530
rect 50540 49478 50570 49530
rect 50570 49478 50596 49530
rect 50300 49476 50356 49478
rect 50380 49476 50436 49478
rect 50460 49476 50516 49478
rect 50540 49476 50596 49478
rect 50300 48442 50356 48444
rect 50380 48442 50436 48444
rect 50460 48442 50516 48444
rect 50540 48442 50596 48444
rect 50300 48390 50326 48442
rect 50326 48390 50356 48442
rect 50380 48390 50390 48442
rect 50390 48390 50436 48442
rect 50460 48390 50506 48442
rect 50506 48390 50516 48442
rect 50540 48390 50570 48442
rect 50570 48390 50596 48442
rect 50300 48388 50356 48390
rect 50380 48388 50436 48390
rect 50460 48388 50516 48390
rect 50540 48388 50596 48390
rect 50300 47354 50356 47356
rect 50380 47354 50436 47356
rect 50460 47354 50516 47356
rect 50540 47354 50596 47356
rect 50300 47302 50326 47354
rect 50326 47302 50356 47354
rect 50380 47302 50390 47354
rect 50390 47302 50436 47354
rect 50460 47302 50506 47354
rect 50506 47302 50516 47354
rect 50540 47302 50570 47354
rect 50570 47302 50596 47354
rect 50300 47300 50356 47302
rect 50380 47300 50436 47302
rect 50460 47300 50516 47302
rect 50540 47300 50596 47302
rect 50300 46266 50356 46268
rect 50380 46266 50436 46268
rect 50460 46266 50516 46268
rect 50540 46266 50596 46268
rect 50300 46214 50326 46266
rect 50326 46214 50356 46266
rect 50380 46214 50390 46266
rect 50390 46214 50436 46266
rect 50460 46214 50506 46266
rect 50506 46214 50516 46266
rect 50540 46214 50570 46266
rect 50570 46214 50596 46266
rect 50300 46212 50356 46214
rect 50380 46212 50436 46214
rect 50460 46212 50516 46214
rect 50540 46212 50596 46214
rect 50300 45178 50356 45180
rect 50380 45178 50436 45180
rect 50460 45178 50516 45180
rect 50540 45178 50596 45180
rect 50300 45126 50326 45178
rect 50326 45126 50356 45178
rect 50380 45126 50390 45178
rect 50390 45126 50436 45178
rect 50460 45126 50506 45178
rect 50506 45126 50516 45178
rect 50540 45126 50570 45178
rect 50570 45126 50596 45178
rect 50300 45124 50356 45126
rect 50380 45124 50436 45126
rect 50460 45124 50516 45126
rect 50540 45124 50596 45126
rect 50300 44090 50356 44092
rect 50380 44090 50436 44092
rect 50460 44090 50516 44092
rect 50540 44090 50596 44092
rect 50300 44038 50326 44090
rect 50326 44038 50356 44090
rect 50380 44038 50390 44090
rect 50390 44038 50436 44090
rect 50460 44038 50506 44090
rect 50506 44038 50516 44090
rect 50540 44038 50570 44090
rect 50570 44038 50596 44090
rect 50300 44036 50356 44038
rect 50380 44036 50436 44038
rect 50460 44036 50516 44038
rect 50540 44036 50596 44038
rect 50300 43002 50356 43004
rect 50380 43002 50436 43004
rect 50460 43002 50516 43004
rect 50540 43002 50596 43004
rect 50300 42950 50326 43002
rect 50326 42950 50356 43002
rect 50380 42950 50390 43002
rect 50390 42950 50436 43002
rect 50460 42950 50506 43002
rect 50506 42950 50516 43002
rect 50540 42950 50570 43002
rect 50570 42950 50596 43002
rect 50300 42948 50356 42950
rect 50380 42948 50436 42950
rect 50460 42948 50516 42950
rect 50540 42948 50596 42950
rect 50300 41914 50356 41916
rect 50380 41914 50436 41916
rect 50460 41914 50516 41916
rect 50540 41914 50596 41916
rect 50300 41862 50326 41914
rect 50326 41862 50356 41914
rect 50380 41862 50390 41914
rect 50390 41862 50436 41914
rect 50460 41862 50506 41914
rect 50506 41862 50516 41914
rect 50540 41862 50570 41914
rect 50570 41862 50596 41914
rect 50300 41860 50356 41862
rect 50380 41860 50436 41862
rect 50460 41860 50516 41862
rect 50540 41860 50596 41862
rect 50300 40826 50356 40828
rect 50380 40826 50436 40828
rect 50460 40826 50516 40828
rect 50540 40826 50596 40828
rect 50300 40774 50326 40826
rect 50326 40774 50356 40826
rect 50380 40774 50390 40826
rect 50390 40774 50436 40826
rect 50460 40774 50506 40826
rect 50506 40774 50516 40826
rect 50540 40774 50570 40826
rect 50570 40774 50596 40826
rect 50300 40772 50356 40774
rect 50380 40772 50436 40774
rect 50460 40772 50516 40774
rect 50540 40772 50596 40774
rect 50300 39738 50356 39740
rect 50380 39738 50436 39740
rect 50460 39738 50516 39740
rect 50540 39738 50596 39740
rect 50300 39686 50326 39738
rect 50326 39686 50356 39738
rect 50380 39686 50390 39738
rect 50390 39686 50436 39738
rect 50460 39686 50506 39738
rect 50506 39686 50516 39738
rect 50540 39686 50570 39738
rect 50570 39686 50596 39738
rect 50300 39684 50356 39686
rect 50380 39684 50436 39686
rect 50460 39684 50516 39686
rect 50540 39684 50596 39686
rect 50300 38650 50356 38652
rect 50380 38650 50436 38652
rect 50460 38650 50516 38652
rect 50540 38650 50596 38652
rect 50300 38598 50326 38650
rect 50326 38598 50356 38650
rect 50380 38598 50390 38650
rect 50390 38598 50436 38650
rect 50460 38598 50506 38650
rect 50506 38598 50516 38650
rect 50540 38598 50570 38650
rect 50570 38598 50596 38650
rect 50300 38596 50356 38598
rect 50380 38596 50436 38598
rect 50460 38596 50516 38598
rect 50540 38596 50596 38598
rect 50300 37562 50356 37564
rect 50380 37562 50436 37564
rect 50460 37562 50516 37564
rect 50540 37562 50596 37564
rect 50300 37510 50326 37562
rect 50326 37510 50356 37562
rect 50380 37510 50390 37562
rect 50390 37510 50436 37562
rect 50460 37510 50506 37562
rect 50506 37510 50516 37562
rect 50540 37510 50570 37562
rect 50570 37510 50596 37562
rect 50300 37508 50356 37510
rect 50380 37508 50436 37510
rect 50460 37508 50516 37510
rect 50540 37508 50596 37510
rect 50300 36474 50356 36476
rect 50380 36474 50436 36476
rect 50460 36474 50516 36476
rect 50540 36474 50596 36476
rect 50300 36422 50326 36474
rect 50326 36422 50356 36474
rect 50380 36422 50390 36474
rect 50390 36422 50436 36474
rect 50460 36422 50506 36474
rect 50506 36422 50516 36474
rect 50540 36422 50570 36474
rect 50570 36422 50596 36474
rect 50300 36420 50356 36422
rect 50380 36420 50436 36422
rect 50460 36420 50516 36422
rect 50540 36420 50596 36422
rect 50300 35386 50356 35388
rect 50380 35386 50436 35388
rect 50460 35386 50516 35388
rect 50540 35386 50596 35388
rect 50300 35334 50326 35386
rect 50326 35334 50356 35386
rect 50380 35334 50390 35386
rect 50390 35334 50436 35386
rect 50460 35334 50506 35386
rect 50506 35334 50516 35386
rect 50540 35334 50570 35386
rect 50570 35334 50596 35386
rect 50300 35332 50356 35334
rect 50380 35332 50436 35334
rect 50460 35332 50516 35334
rect 50540 35332 50596 35334
rect 50300 34298 50356 34300
rect 50380 34298 50436 34300
rect 50460 34298 50516 34300
rect 50540 34298 50596 34300
rect 50300 34246 50326 34298
rect 50326 34246 50356 34298
rect 50380 34246 50390 34298
rect 50390 34246 50436 34298
rect 50460 34246 50506 34298
rect 50506 34246 50516 34298
rect 50540 34246 50570 34298
rect 50570 34246 50596 34298
rect 50300 34244 50356 34246
rect 50380 34244 50436 34246
rect 50460 34244 50516 34246
rect 50540 34244 50596 34246
rect 50300 33210 50356 33212
rect 50380 33210 50436 33212
rect 50460 33210 50516 33212
rect 50540 33210 50596 33212
rect 50300 33158 50326 33210
rect 50326 33158 50356 33210
rect 50380 33158 50390 33210
rect 50390 33158 50436 33210
rect 50460 33158 50506 33210
rect 50506 33158 50516 33210
rect 50540 33158 50570 33210
rect 50570 33158 50596 33210
rect 50300 33156 50356 33158
rect 50380 33156 50436 33158
rect 50460 33156 50516 33158
rect 50540 33156 50596 33158
rect 50300 32122 50356 32124
rect 50380 32122 50436 32124
rect 50460 32122 50516 32124
rect 50540 32122 50596 32124
rect 50300 32070 50326 32122
rect 50326 32070 50356 32122
rect 50380 32070 50390 32122
rect 50390 32070 50436 32122
rect 50460 32070 50506 32122
rect 50506 32070 50516 32122
rect 50540 32070 50570 32122
rect 50570 32070 50596 32122
rect 50300 32068 50356 32070
rect 50380 32068 50436 32070
rect 50460 32068 50516 32070
rect 50540 32068 50596 32070
rect 50300 31034 50356 31036
rect 50380 31034 50436 31036
rect 50460 31034 50516 31036
rect 50540 31034 50596 31036
rect 50300 30982 50326 31034
rect 50326 30982 50356 31034
rect 50380 30982 50390 31034
rect 50390 30982 50436 31034
rect 50460 30982 50506 31034
rect 50506 30982 50516 31034
rect 50540 30982 50570 31034
rect 50570 30982 50596 31034
rect 50300 30980 50356 30982
rect 50380 30980 50436 30982
rect 50460 30980 50516 30982
rect 50540 30980 50596 30982
rect 50300 29946 50356 29948
rect 50380 29946 50436 29948
rect 50460 29946 50516 29948
rect 50540 29946 50596 29948
rect 50300 29894 50326 29946
rect 50326 29894 50356 29946
rect 50380 29894 50390 29946
rect 50390 29894 50436 29946
rect 50460 29894 50506 29946
rect 50506 29894 50516 29946
rect 50540 29894 50570 29946
rect 50570 29894 50596 29946
rect 50300 29892 50356 29894
rect 50380 29892 50436 29894
rect 50460 29892 50516 29894
rect 50540 29892 50596 29894
rect 50300 28858 50356 28860
rect 50380 28858 50436 28860
rect 50460 28858 50516 28860
rect 50540 28858 50596 28860
rect 50300 28806 50326 28858
rect 50326 28806 50356 28858
rect 50380 28806 50390 28858
rect 50390 28806 50436 28858
rect 50460 28806 50506 28858
rect 50506 28806 50516 28858
rect 50540 28806 50570 28858
rect 50570 28806 50596 28858
rect 50300 28804 50356 28806
rect 50380 28804 50436 28806
rect 50460 28804 50516 28806
rect 50540 28804 50596 28806
rect 50300 27770 50356 27772
rect 50380 27770 50436 27772
rect 50460 27770 50516 27772
rect 50540 27770 50596 27772
rect 50300 27718 50326 27770
rect 50326 27718 50356 27770
rect 50380 27718 50390 27770
rect 50390 27718 50436 27770
rect 50460 27718 50506 27770
rect 50506 27718 50516 27770
rect 50540 27718 50570 27770
rect 50570 27718 50596 27770
rect 50300 27716 50356 27718
rect 50380 27716 50436 27718
rect 50460 27716 50516 27718
rect 50540 27716 50596 27718
rect 50300 26682 50356 26684
rect 50380 26682 50436 26684
rect 50460 26682 50516 26684
rect 50540 26682 50596 26684
rect 50300 26630 50326 26682
rect 50326 26630 50356 26682
rect 50380 26630 50390 26682
rect 50390 26630 50436 26682
rect 50460 26630 50506 26682
rect 50506 26630 50516 26682
rect 50540 26630 50570 26682
rect 50570 26630 50596 26682
rect 50300 26628 50356 26630
rect 50380 26628 50436 26630
rect 50460 26628 50516 26630
rect 50540 26628 50596 26630
rect 50300 25594 50356 25596
rect 50380 25594 50436 25596
rect 50460 25594 50516 25596
rect 50540 25594 50596 25596
rect 50300 25542 50326 25594
rect 50326 25542 50356 25594
rect 50380 25542 50390 25594
rect 50390 25542 50436 25594
rect 50460 25542 50506 25594
rect 50506 25542 50516 25594
rect 50540 25542 50570 25594
rect 50570 25542 50596 25594
rect 50300 25540 50356 25542
rect 50380 25540 50436 25542
rect 50460 25540 50516 25542
rect 50540 25540 50596 25542
rect 50300 24506 50356 24508
rect 50380 24506 50436 24508
rect 50460 24506 50516 24508
rect 50540 24506 50596 24508
rect 50300 24454 50326 24506
rect 50326 24454 50356 24506
rect 50380 24454 50390 24506
rect 50390 24454 50436 24506
rect 50460 24454 50506 24506
rect 50506 24454 50516 24506
rect 50540 24454 50570 24506
rect 50570 24454 50596 24506
rect 50300 24452 50356 24454
rect 50380 24452 50436 24454
rect 50460 24452 50516 24454
rect 50540 24452 50596 24454
rect 50300 23418 50356 23420
rect 50380 23418 50436 23420
rect 50460 23418 50516 23420
rect 50540 23418 50596 23420
rect 50300 23366 50326 23418
rect 50326 23366 50356 23418
rect 50380 23366 50390 23418
rect 50390 23366 50436 23418
rect 50460 23366 50506 23418
rect 50506 23366 50516 23418
rect 50540 23366 50570 23418
rect 50570 23366 50596 23418
rect 50300 23364 50356 23366
rect 50380 23364 50436 23366
rect 50460 23364 50516 23366
rect 50540 23364 50596 23366
rect 50300 22330 50356 22332
rect 50380 22330 50436 22332
rect 50460 22330 50516 22332
rect 50540 22330 50596 22332
rect 50300 22278 50326 22330
rect 50326 22278 50356 22330
rect 50380 22278 50390 22330
rect 50390 22278 50436 22330
rect 50460 22278 50506 22330
rect 50506 22278 50516 22330
rect 50540 22278 50570 22330
rect 50570 22278 50596 22330
rect 50300 22276 50356 22278
rect 50380 22276 50436 22278
rect 50460 22276 50516 22278
rect 50540 22276 50596 22278
rect 50300 21242 50356 21244
rect 50380 21242 50436 21244
rect 50460 21242 50516 21244
rect 50540 21242 50596 21244
rect 50300 21190 50326 21242
rect 50326 21190 50356 21242
rect 50380 21190 50390 21242
rect 50390 21190 50436 21242
rect 50460 21190 50506 21242
rect 50506 21190 50516 21242
rect 50540 21190 50570 21242
rect 50570 21190 50596 21242
rect 50300 21188 50356 21190
rect 50380 21188 50436 21190
rect 50460 21188 50516 21190
rect 50540 21188 50596 21190
rect 50300 20154 50356 20156
rect 50380 20154 50436 20156
rect 50460 20154 50516 20156
rect 50540 20154 50596 20156
rect 50300 20102 50326 20154
rect 50326 20102 50356 20154
rect 50380 20102 50390 20154
rect 50390 20102 50436 20154
rect 50460 20102 50506 20154
rect 50506 20102 50516 20154
rect 50540 20102 50570 20154
rect 50570 20102 50596 20154
rect 50300 20100 50356 20102
rect 50380 20100 50436 20102
rect 50460 20100 50516 20102
rect 50540 20100 50596 20102
rect 50300 19066 50356 19068
rect 50380 19066 50436 19068
rect 50460 19066 50516 19068
rect 50540 19066 50596 19068
rect 50300 19014 50326 19066
rect 50326 19014 50356 19066
rect 50380 19014 50390 19066
rect 50390 19014 50436 19066
rect 50460 19014 50506 19066
rect 50506 19014 50516 19066
rect 50540 19014 50570 19066
rect 50570 19014 50596 19066
rect 50300 19012 50356 19014
rect 50380 19012 50436 19014
rect 50460 19012 50516 19014
rect 50540 19012 50596 19014
rect 50300 17978 50356 17980
rect 50380 17978 50436 17980
rect 50460 17978 50516 17980
rect 50540 17978 50596 17980
rect 50300 17926 50326 17978
rect 50326 17926 50356 17978
rect 50380 17926 50390 17978
rect 50390 17926 50436 17978
rect 50460 17926 50506 17978
rect 50506 17926 50516 17978
rect 50540 17926 50570 17978
rect 50570 17926 50596 17978
rect 50300 17924 50356 17926
rect 50380 17924 50436 17926
rect 50460 17924 50516 17926
rect 50540 17924 50596 17926
rect 50300 16890 50356 16892
rect 50380 16890 50436 16892
rect 50460 16890 50516 16892
rect 50540 16890 50596 16892
rect 50300 16838 50326 16890
rect 50326 16838 50356 16890
rect 50380 16838 50390 16890
rect 50390 16838 50436 16890
rect 50460 16838 50506 16890
rect 50506 16838 50516 16890
rect 50540 16838 50570 16890
rect 50570 16838 50596 16890
rect 50300 16836 50356 16838
rect 50380 16836 50436 16838
rect 50460 16836 50516 16838
rect 50540 16836 50596 16838
rect 50300 15802 50356 15804
rect 50380 15802 50436 15804
rect 50460 15802 50516 15804
rect 50540 15802 50596 15804
rect 50300 15750 50326 15802
rect 50326 15750 50356 15802
rect 50380 15750 50390 15802
rect 50390 15750 50436 15802
rect 50460 15750 50506 15802
rect 50506 15750 50516 15802
rect 50540 15750 50570 15802
rect 50570 15750 50596 15802
rect 50300 15748 50356 15750
rect 50380 15748 50436 15750
rect 50460 15748 50516 15750
rect 50540 15748 50596 15750
rect 50300 14714 50356 14716
rect 50380 14714 50436 14716
rect 50460 14714 50516 14716
rect 50540 14714 50596 14716
rect 50300 14662 50326 14714
rect 50326 14662 50356 14714
rect 50380 14662 50390 14714
rect 50390 14662 50436 14714
rect 50460 14662 50506 14714
rect 50506 14662 50516 14714
rect 50540 14662 50570 14714
rect 50570 14662 50596 14714
rect 50300 14660 50356 14662
rect 50380 14660 50436 14662
rect 50460 14660 50516 14662
rect 50540 14660 50596 14662
rect 50300 13626 50356 13628
rect 50380 13626 50436 13628
rect 50460 13626 50516 13628
rect 50540 13626 50596 13628
rect 50300 13574 50326 13626
rect 50326 13574 50356 13626
rect 50380 13574 50390 13626
rect 50390 13574 50436 13626
rect 50460 13574 50506 13626
rect 50506 13574 50516 13626
rect 50540 13574 50570 13626
rect 50570 13574 50596 13626
rect 50300 13572 50356 13574
rect 50380 13572 50436 13574
rect 50460 13572 50516 13574
rect 50540 13572 50596 13574
rect 50300 12538 50356 12540
rect 50380 12538 50436 12540
rect 50460 12538 50516 12540
rect 50540 12538 50596 12540
rect 50300 12486 50326 12538
rect 50326 12486 50356 12538
rect 50380 12486 50390 12538
rect 50390 12486 50436 12538
rect 50460 12486 50506 12538
rect 50506 12486 50516 12538
rect 50540 12486 50570 12538
rect 50570 12486 50596 12538
rect 50300 12484 50356 12486
rect 50380 12484 50436 12486
rect 50460 12484 50516 12486
rect 50540 12484 50596 12486
rect 50300 11450 50356 11452
rect 50380 11450 50436 11452
rect 50460 11450 50516 11452
rect 50540 11450 50596 11452
rect 50300 11398 50326 11450
rect 50326 11398 50356 11450
rect 50380 11398 50390 11450
rect 50390 11398 50436 11450
rect 50460 11398 50506 11450
rect 50506 11398 50516 11450
rect 50540 11398 50570 11450
rect 50570 11398 50596 11450
rect 50300 11396 50356 11398
rect 50380 11396 50436 11398
rect 50460 11396 50516 11398
rect 50540 11396 50596 11398
rect 50300 10362 50356 10364
rect 50380 10362 50436 10364
rect 50460 10362 50516 10364
rect 50540 10362 50596 10364
rect 50300 10310 50326 10362
rect 50326 10310 50356 10362
rect 50380 10310 50390 10362
rect 50390 10310 50436 10362
rect 50460 10310 50506 10362
rect 50506 10310 50516 10362
rect 50540 10310 50570 10362
rect 50570 10310 50596 10362
rect 50300 10308 50356 10310
rect 50380 10308 50436 10310
rect 50460 10308 50516 10310
rect 50540 10308 50596 10310
rect 50300 9274 50356 9276
rect 50380 9274 50436 9276
rect 50460 9274 50516 9276
rect 50540 9274 50596 9276
rect 50300 9222 50326 9274
rect 50326 9222 50356 9274
rect 50380 9222 50390 9274
rect 50390 9222 50436 9274
rect 50460 9222 50506 9274
rect 50506 9222 50516 9274
rect 50540 9222 50570 9274
rect 50570 9222 50596 9274
rect 50300 9220 50356 9222
rect 50380 9220 50436 9222
rect 50460 9220 50516 9222
rect 50540 9220 50596 9222
rect 50300 8186 50356 8188
rect 50380 8186 50436 8188
rect 50460 8186 50516 8188
rect 50540 8186 50596 8188
rect 50300 8134 50326 8186
rect 50326 8134 50356 8186
rect 50380 8134 50390 8186
rect 50390 8134 50436 8186
rect 50460 8134 50506 8186
rect 50506 8134 50516 8186
rect 50540 8134 50570 8186
rect 50570 8134 50596 8186
rect 50300 8132 50356 8134
rect 50380 8132 50436 8134
rect 50460 8132 50516 8134
rect 50540 8132 50596 8134
rect 50300 7098 50356 7100
rect 50380 7098 50436 7100
rect 50460 7098 50516 7100
rect 50540 7098 50596 7100
rect 50300 7046 50326 7098
rect 50326 7046 50356 7098
rect 50380 7046 50390 7098
rect 50390 7046 50436 7098
rect 50460 7046 50506 7098
rect 50506 7046 50516 7098
rect 50540 7046 50570 7098
rect 50570 7046 50596 7098
rect 50300 7044 50356 7046
rect 50380 7044 50436 7046
rect 50460 7044 50516 7046
rect 50540 7044 50596 7046
rect 50300 6010 50356 6012
rect 50380 6010 50436 6012
rect 50460 6010 50516 6012
rect 50540 6010 50596 6012
rect 50300 5958 50326 6010
rect 50326 5958 50356 6010
rect 50380 5958 50390 6010
rect 50390 5958 50436 6010
rect 50460 5958 50506 6010
rect 50506 5958 50516 6010
rect 50540 5958 50570 6010
rect 50570 5958 50596 6010
rect 50300 5956 50356 5958
rect 50380 5956 50436 5958
rect 50460 5956 50516 5958
rect 50540 5956 50596 5958
rect 50300 4922 50356 4924
rect 50380 4922 50436 4924
rect 50460 4922 50516 4924
rect 50540 4922 50596 4924
rect 50300 4870 50326 4922
rect 50326 4870 50356 4922
rect 50380 4870 50390 4922
rect 50390 4870 50436 4922
rect 50460 4870 50506 4922
rect 50506 4870 50516 4922
rect 50540 4870 50570 4922
rect 50570 4870 50596 4922
rect 50300 4868 50356 4870
rect 50380 4868 50436 4870
rect 50460 4868 50516 4870
rect 50540 4868 50596 4870
rect 50300 3834 50356 3836
rect 50380 3834 50436 3836
rect 50460 3834 50516 3836
rect 50540 3834 50596 3836
rect 50300 3782 50326 3834
rect 50326 3782 50356 3834
rect 50380 3782 50390 3834
rect 50390 3782 50436 3834
rect 50460 3782 50506 3834
rect 50506 3782 50516 3834
rect 50540 3782 50570 3834
rect 50570 3782 50596 3834
rect 50300 3780 50356 3782
rect 50380 3780 50436 3782
rect 50460 3780 50516 3782
rect 50540 3780 50596 3782
rect 50300 2746 50356 2748
rect 50380 2746 50436 2748
rect 50460 2746 50516 2748
rect 50540 2746 50596 2748
rect 50300 2694 50326 2746
rect 50326 2694 50356 2746
rect 50380 2694 50390 2746
rect 50390 2694 50436 2746
rect 50460 2694 50506 2746
rect 50506 2694 50516 2746
rect 50540 2694 50570 2746
rect 50570 2694 50596 2746
rect 50300 2692 50356 2694
rect 50380 2692 50436 2694
rect 50460 2692 50516 2694
rect 50540 2692 50596 2694
rect 57426 70352 57482 70408
rect 57886 70352 57942 70408
rect 62670 63824 62726 63880
rect 62946 10004 62948 10024
rect 62948 10004 63000 10024
rect 63000 10004 63002 10024
rect 62946 9968 63002 10004
rect 62762 9832 62818 9888
rect 65660 96858 65716 96860
rect 65740 96858 65796 96860
rect 65820 96858 65876 96860
rect 65900 96858 65956 96860
rect 65660 96806 65686 96858
rect 65686 96806 65716 96858
rect 65740 96806 65750 96858
rect 65750 96806 65796 96858
rect 65820 96806 65866 96858
rect 65866 96806 65876 96858
rect 65900 96806 65930 96858
rect 65930 96806 65956 96858
rect 65660 96804 65716 96806
rect 65740 96804 65796 96806
rect 65820 96804 65876 96806
rect 65900 96804 65956 96806
rect 63590 9832 63646 9888
rect 63866 10004 63868 10024
rect 63868 10004 63920 10024
rect 63920 10004 63922 10024
rect 63866 9968 63922 10004
rect 65660 95770 65716 95772
rect 65740 95770 65796 95772
rect 65820 95770 65876 95772
rect 65900 95770 65956 95772
rect 65660 95718 65686 95770
rect 65686 95718 65716 95770
rect 65740 95718 65750 95770
rect 65750 95718 65796 95770
rect 65820 95718 65866 95770
rect 65866 95718 65876 95770
rect 65900 95718 65930 95770
rect 65930 95718 65956 95770
rect 65660 95716 65716 95718
rect 65740 95716 65796 95718
rect 65820 95716 65876 95718
rect 65900 95716 65956 95718
rect 65660 94682 65716 94684
rect 65740 94682 65796 94684
rect 65820 94682 65876 94684
rect 65900 94682 65956 94684
rect 65660 94630 65686 94682
rect 65686 94630 65716 94682
rect 65740 94630 65750 94682
rect 65750 94630 65796 94682
rect 65820 94630 65866 94682
rect 65866 94630 65876 94682
rect 65900 94630 65930 94682
rect 65930 94630 65956 94682
rect 65660 94628 65716 94630
rect 65740 94628 65796 94630
rect 65820 94628 65876 94630
rect 65900 94628 65956 94630
rect 65660 93594 65716 93596
rect 65740 93594 65796 93596
rect 65820 93594 65876 93596
rect 65900 93594 65956 93596
rect 65660 93542 65686 93594
rect 65686 93542 65716 93594
rect 65740 93542 65750 93594
rect 65750 93542 65796 93594
rect 65820 93542 65866 93594
rect 65866 93542 65876 93594
rect 65900 93542 65930 93594
rect 65930 93542 65956 93594
rect 65660 93540 65716 93542
rect 65740 93540 65796 93542
rect 65820 93540 65876 93542
rect 65900 93540 65956 93542
rect 65660 92506 65716 92508
rect 65740 92506 65796 92508
rect 65820 92506 65876 92508
rect 65900 92506 65956 92508
rect 65660 92454 65686 92506
rect 65686 92454 65716 92506
rect 65740 92454 65750 92506
rect 65750 92454 65796 92506
rect 65820 92454 65866 92506
rect 65866 92454 65876 92506
rect 65900 92454 65930 92506
rect 65930 92454 65956 92506
rect 65660 92452 65716 92454
rect 65740 92452 65796 92454
rect 65820 92452 65876 92454
rect 65900 92452 65956 92454
rect 65660 91418 65716 91420
rect 65740 91418 65796 91420
rect 65820 91418 65876 91420
rect 65900 91418 65956 91420
rect 65660 91366 65686 91418
rect 65686 91366 65716 91418
rect 65740 91366 65750 91418
rect 65750 91366 65796 91418
rect 65820 91366 65866 91418
rect 65866 91366 65876 91418
rect 65900 91366 65930 91418
rect 65930 91366 65956 91418
rect 65660 91364 65716 91366
rect 65740 91364 65796 91366
rect 65820 91364 65876 91366
rect 65900 91364 65956 91366
rect 65660 90330 65716 90332
rect 65740 90330 65796 90332
rect 65820 90330 65876 90332
rect 65900 90330 65956 90332
rect 65660 90278 65686 90330
rect 65686 90278 65716 90330
rect 65740 90278 65750 90330
rect 65750 90278 65796 90330
rect 65820 90278 65866 90330
rect 65866 90278 65876 90330
rect 65900 90278 65930 90330
rect 65930 90278 65956 90330
rect 65660 90276 65716 90278
rect 65740 90276 65796 90278
rect 65820 90276 65876 90278
rect 65900 90276 65956 90278
rect 65660 89242 65716 89244
rect 65740 89242 65796 89244
rect 65820 89242 65876 89244
rect 65900 89242 65956 89244
rect 65660 89190 65686 89242
rect 65686 89190 65716 89242
rect 65740 89190 65750 89242
rect 65750 89190 65796 89242
rect 65820 89190 65866 89242
rect 65866 89190 65876 89242
rect 65900 89190 65930 89242
rect 65930 89190 65956 89242
rect 65660 89188 65716 89190
rect 65740 89188 65796 89190
rect 65820 89188 65876 89190
rect 65900 89188 65956 89190
rect 65660 88154 65716 88156
rect 65740 88154 65796 88156
rect 65820 88154 65876 88156
rect 65900 88154 65956 88156
rect 65660 88102 65686 88154
rect 65686 88102 65716 88154
rect 65740 88102 65750 88154
rect 65750 88102 65796 88154
rect 65820 88102 65866 88154
rect 65866 88102 65876 88154
rect 65900 88102 65930 88154
rect 65930 88102 65956 88154
rect 65660 88100 65716 88102
rect 65740 88100 65796 88102
rect 65820 88100 65876 88102
rect 65900 88100 65956 88102
rect 65660 87066 65716 87068
rect 65740 87066 65796 87068
rect 65820 87066 65876 87068
rect 65900 87066 65956 87068
rect 65660 87014 65686 87066
rect 65686 87014 65716 87066
rect 65740 87014 65750 87066
rect 65750 87014 65796 87066
rect 65820 87014 65866 87066
rect 65866 87014 65876 87066
rect 65900 87014 65930 87066
rect 65930 87014 65956 87066
rect 65660 87012 65716 87014
rect 65740 87012 65796 87014
rect 65820 87012 65876 87014
rect 65900 87012 65956 87014
rect 65660 85978 65716 85980
rect 65740 85978 65796 85980
rect 65820 85978 65876 85980
rect 65900 85978 65956 85980
rect 65660 85926 65686 85978
rect 65686 85926 65716 85978
rect 65740 85926 65750 85978
rect 65750 85926 65796 85978
rect 65820 85926 65866 85978
rect 65866 85926 65876 85978
rect 65900 85926 65930 85978
rect 65930 85926 65956 85978
rect 65660 85924 65716 85926
rect 65740 85924 65796 85926
rect 65820 85924 65876 85926
rect 65900 85924 65956 85926
rect 65660 84890 65716 84892
rect 65740 84890 65796 84892
rect 65820 84890 65876 84892
rect 65900 84890 65956 84892
rect 65660 84838 65686 84890
rect 65686 84838 65716 84890
rect 65740 84838 65750 84890
rect 65750 84838 65796 84890
rect 65820 84838 65866 84890
rect 65866 84838 65876 84890
rect 65900 84838 65930 84890
rect 65930 84838 65956 84890
rect 65660 84836 65716 84838
rect 65740 84836 65796 84838
rect 65820 84836 65876 84838
rect 65900 84836 65956 84838
rect 65660 83802 65716 83804
rect 65740 83802 65796 83804
rect 65820 83802 65876 83804
rect 65900 83802 65956 83804
rect 65660 83750 65686 83802
rect 65686 83750 65716 83802
rect 65740 83750 65750 83802
rect 65750 83750 65796 83802
rect 65820 83750 65866 83802
rect 65866 83750 65876 83802
rect 65900 83750 65930 83802
rect 65930 83750 65956 83802
rect 65660 83748 65716 83750
rect 65740 83748 65796 83750
rect 65820 83748 65876 83750
rect 65900 83748 65956 83750
rect 65660 82714 65716 82716
rect 65740 82714 65796 82716
rect 65820 82714 65876 82716
rect 65900 82714 65956 82716
rect 65660 82662 65686 82714
rect 65686 82662 65716 82714
rect 65740 82662 65750 82714
rect 65750 82662 65796 82714
rect 65820 82662 65866 82714
rect 65866 82662 65876 82714
rect 65900 82662 65930 82714
rect 65930 82662 65956 82714
rect 65660 82660 65716 82662
rect 65740 82660 65796 82662
rect 65820 82660 65876 82662
rect 65900 82660 65956 82662
rect 65660 81626 65716 81628
rect 65740 81626 65796 81628
rect 65820 81626 65876 81628
rect 65900 81626 65956 81628
rect 65660 81574 65686 81626
rect 65686 81574 65716 81626
rect 65740 81574 65750 81626
rect 65750 81574 65796 81626
rect 65820 81574 65866 81626
rect 65866 81574 65876 81626
rect 65900 81574 65930 81626
rect 65930 81574 65956 81626
rect 65660 81572 65716 81574
rect 65740 81572 65796 81574
rect 65820 81572 65876 81574
rect 65900 81572 65956 81574
rect 65660 80538 65716 80540
rect 65740 80538 65796 80540
rect 65820 80538 65876 80540
rect 65900 80538 65956 80540
rect 65660 80486 65686 80538
rect 65686 80486 65716 80538
rect 65740 80486 65750 80538
rect 65750 80486 65796 80538
rect 65820 80486 65866 80538
rect 65866 80486 65876 80538
rect 65900 80486 65930 80538
rect 65930 80486 65956 80538
rect 65660 80484 65716 80486
rect 65740 80484 65796 80486
rect 65820 80484 65876 80486
rect 65900 80484 65956 80486
rect 65660 79450 65716 79452
rect 65740 79450 65796 79452
rect 65820 79450 65876 79452
rect 65900 79450 65956 79452
rect 65660 79398 65686 79450
rect 65686 79398 65716 79450
rect 65740 79398 65750 79450
rect 65750 79398 65796 79450
rect 65820 79398 65866 79450
rect 65866 79398 65876 79450
rect 65900 79398 65930 79450
rect 65930 79398 65956 79450
rect 65660 79396 65716 79398
rect 65740 79396 65796 79398
rect 65820 79396 65876 79398
rect 65900 79396 65956 79398
rect 65660 78362 65716 78364
rect 65740 78362 65796 78364
rect 65820 78362 65876 78364
rect 65900 78362 65956 78364
rect 65660 78310 65686 78362
rect 65686 78310 65716 78362
rect 65740 78310 65750 78362
rect 65750 78310 65796 78362
rect 65820 78310 65866 78362
rect 65866 78310 65876 78362
rect 65900 78310 65930 78362
rect 65930 78310 65956 78362
rect 65660 78308 65716 78310
rect 65740 78308 65796 78310
rect 65820 78308 65876 78310
rect 65900 78308 65956 78310
rect 65660 77274 65716 77276
rect 65740 77274 65796 77276
rect 65820 77274 65876 77276
rect 65900 77274 65956 77276
rect 65660 77222 65686 77274
rect 65686 77222 65716 77274
rect 65740 77222 65750 77274
rect 65750 77222 65796 77274
rect 65820 77222 65866 77274
rect 65866 77222 65876 77274
rect 65900 77222 65930 77274
rect 65930 77222 65956 77274
rect 65660 77220 65716 77222
rect 65740 77220 65796 77222
rect 65820 77220 65876 77222
rect 65900 77220 65956 77222
rect 65660 76186 65716 76188
rect 65740 76186 65796 76188
rect 65820 76186 65876 76188
rect 65900 76186 65956 76188
rect 65660 76134 65686 76186
rect 65686 76134 65716 76186
rect 65740 76134 65750 76186
rect 65750 76134 65796 76186
rect 65820 76134 65866 76186
rect 65866 76134 65876 76186
rect 65900 76134 65930 76186
rect 65930 76134 65956 76186
rect 65660 76132 65716 76134
rect 65740 76132 65796 76134
rect 65820 76132 65876 76134
rect 65900 76132 65956 76134
rect 65660 75098 65716 75100
rect 65740 75098 65796 75100
rect 65820 75098 65876 75100
rect 65900 75098 65956 75100
rect 65660 75046 65686 75098
rect 65686 75046 65716 75098
rect 65740 75046 65750 75098
rect 65750 75046 65796 75098
rect 65820 75046 65866 75098
rect 65866 75046 65876 75098
rect 65900 75046 65930 75098
rect 65930 75046 65956 75098
rect 65660 75044 65716 75046
rect 65740 75044 65796 75046
rect 65820 75044 65876 75046
rect 65900 75044 65956 75046
rect 65660 74010 65716 74012
rect 65740 74010 65796 74012
rect 65820 74010 65876 74012
rect 65900 74010 65956 74012
rect 65660 73958 65686 74010
rect 65686 73958 65716 74010
rect 65740 73958 65750 74010
rect 65750 73958 65796 74010
rect 65820 73958 65866 74010
rect 65866 73958 65876 74010
rect 65900 73958 65930 74010
rect 65930 73958 65956 74010
rect 65660 73956 65716 73958
rect 65740 73956 65796 73958
rect 65820 73956 65876 73958
rect 65900 73956 65956 73958
rect 65660 72922 65716 72924
rect 65740 72922 65796 72924
rect 65820 72922 65876 72924
rect 65900 72922 65956 72924
rect 65660 72870 65686 72922
rect 65686 72870 65716 72922
rect 65740 72870 65750 72922
rect 65750 72870 65796 72922
rect 65820 72870 65866 72922
rect 65866 72870 65876 72922
rect 65900 72870 65930 72922
rect 65930 72870 65956 72922
rect 65660 72868 65716 72870
rect 65740 72868 65796 72870
rect 65820 72868 65876 72870
rect 65900 72868 65956 72870
rect 65660 71834 65716 71836
rect 65740 71834 65796 71836
rect 65820 71834 65876 71836
rect 65900 71834 65956 71836
rect 65660 71782 65686 71834
rect 65686 71782 65716 71834
rect 65740 71782 65750 71834
rect 65750 71782 65796 71834
rect 65820 71782 65866 71834
rect 65866 71782 65876 71834
rect 65900 71782 65930 71834
rect 65930 71782 65956 71834
rect 65660 71780 65716 71782
rect 65740 71780 65796 71782
rect 65820 71780 65876 71782
rect 65900 71780 65956 71782
rect 65660 70746 65716 70748
rect 65740 70746 65796 70748
rect 65820 70746 65876 70748
rect 65900 70746 65956 70748
rect 65660 70694 65686 70746
rect 65686 70694 65716 70746
rect 65740 70694 65750 70746
rect 65750 70694 65796 70746
rect 65820 70694 65866 70746
rect 65866 70694 65876 70746
rect 65900 70694 65930 70746
rect 65930 70694 65956 70746
rect 65660 70692 65716 70694
rect 65740 70692 65796 70694
rect 65820 70692 65876 70694
rect 65900 70692 65956 70694
rect 65660 69658 65716 69660
rect 65740 69658 65796 69660
rect 65820 69658 65876 69660
rect 65900 69658 65956 69660
rect 65660 69606 65686 69658
rect 65686 69606 65716 69658
rect 65740 69606 65750 69658
rect 65750 69606 65796 69658
rect 65820 69606 65866 69658
rect 65866 69606 65876 69658
rect 65900 69606 65930 69658
rect 65930 69606 65956 69658
rect 65660 69604 65716 69606
rect 65740 69604 65796 69606
rect 65820 69604 65876 69606
rect 65900 69604 65956 69606
rect 65660 68570 65716 68572
rect 65740 68570 65796 68572
rect 65820 68570 65876 68572
rect 65900 68570 65956 68572
rect 65660 68518 65686 68570
rect 65686 68518 65716 68570
rect 65740 68518 65750 68570
rect 65750 68518 65796 68570
rect 65820 68518 65866 68570
rect 65866 68518 65876 68570
rect 65900 68518 65930 68570
rect 65930 68518 65956 68570
rect 65660 68516 65716 68518
rect 65740 68516 65796 68518
rect 65820 68516 65876 68518
rect 65900 68516 65956 68518
rect 65660 67482 65716 67484
rect 65740 67482 65796 67484
rect 65820 67482 65876 67484
rect 65900 67482 65956 67484
rect 65660 67430 65686 67482
rect 65686 67430 65716 67482
rect 65740 67430 65750 67482
rect 65750 67430 65796 67482
rect 65820 67430 65866 67482
rect 65866 67430 65876 67482
rect 65900 67430 65930 67482
rect 65930 67430 65956 67482
rect 65660 67428 65716 67430
rect 65740 67428 65796 67430
rect 65820 67428 65876 67430
rect 65900 67428 65956 67430
rect 65660 66394 65716 66396
rect 65740 66394 65796 66396
rect 65820 66394 65876 66396
rect 65900 66394 65956 66396
rect 65660 66342 65686 66394
rect 65686 66342 65716 66394
rect 65740 66342 65750 66394
rect 65750 66342 65796 66394
rect 65820 66342 65866 66394
rect 65866 66342 65876 66394
rect 65900 66342 65930 66394
rect 65930 66342 65956 66394
rect 65660 66340 65716 66342
rect 65740 66340 65796 66342
rect 65820 66340 65876 66342
rect 65900 66340 65956 66342
rect 65660 65306 65716 65308
rect 65740 65306 65796 65308
rect 65820 65306 65876 65308
rect 65900 65306 65956 65308
rect 65660 65254 65686 65306
rect 65686 65254 65716 65306
rect 65740 65254 65750 65306
rect 65750 65254 65796 65306
rect 65820 65254 65866 65306
rect 65866 65254 65876 65306
rect 65900 65254 65930 65306
rect 65930 65254 65956 65306
rect 65660 65252 65716 65254
rect 65740 65252 65796 65254
rect 65820 65252 65876 65254
rect 65900 65252 65956 65254
rect 65660 64218 65716 64220
rect 65740 64218 65796 64220
rect 65820 64218 65876 64220
rect 65900 64218 65956 64220
rect 65660 64166 65686 64218
rect 65686 64166 65716 64218
rect 65740 64166 65750 64218
rect 65750 64166 65796 64218
rect 65820 64166 65866 64218
rect 65866 64166 65876 64218
rect 65900 64166 65930 64218
rect 65930 64166 65956 64218
rect 65660 64164 65716 64166
rect 65740 64164 65796 64166
rect 65820 64164 65876 64166
rect 65900 64164 65956 64166
rect 65660 63130 65716 63132
rect 65740 63130 65796 63132
rect 65820 63130 65876 63132
rect 65900 63130 65956 63132
rect 65660 63078 65686 63130
rect 65686 63078 65716 63130
rect 65740 63078 65750 63130
rect 65750 63078 65796 63130
rect 65820 63078 65866 63130
rect 65866 63078 65876 63130
rect 65900 63078 65930 63130
rect 65930 63078 65956 63130
rect 65660 63076 65716 63078
rect 65740 63076 65796 63078
rect 65820 63076 65876 63078
rect 65900 63076 65956 63078
rect 65660 62042 65716 62044
rect 65740 62042 65796 62044
rect 65820 62042 65876 62044
rect 65900 62042 65956 62044
rect 65660 61990 65686 62042
rect 65686 61990 65716 62042
rect 65740 61990 65750 62042
rect 65750 61990 65796 62042
rect 65820 61990 65866 62042
rect 65866 61990 65876 62042
rect 65900 61990 65930 62042
rect 65930 61990 65956 62042
rect 65660 61988 65716 61990
rect 65740 61988 65796 61990
rect 65820 61988 65876 61990
rect 65900 61988 65956 61990
rect 65660 60954 65716 60956
rect 65740 60954 65796 60956
rect 65820 60954 65876 60956
rect 65900 60954 65956 60956
rect 65660 60902 65686 60954
rect 65686 60902 65716 60954
rect 65740 60902 65750 60954
rect 65750 60902 65796 60954
rect 65820 60902 65866 60954
rect 65866 60902 65876 60954
rect 65900 60902 65930 60954
rect 65930 60902 65956 60954
rect 65660 60900 65716 60902
rect 65740 60900 65796 60902
rect 65820 60900 65876 60902
rect 65900 60900 65956 60902
rect 65660 59866 65716 59868
rect 65740 59866 65796 59868
rect 65820 59866 65876 59868
rect 65900 59866 65956 59868
rect 65660 59814 65686 59866
rect 65686 59814 65716 59866
rect 65740 59814 65750 59866
rect 65750 59814 65796 59866
rect 65820 59814 65866 59866
rect 65866 59814 65876 59866
rect 65900 59814 65930 59866
rect 65930 59814 65956 59866
rect 65660 59812 65716 59814
rect 65740 59812 65796 59814
rect 65820 59812 65876 59814
rect 65900 59812 65956 59814
rect 65660 58778 65716 58780
rect 65740 58778 65796 58780
rect 65820 58778 65876 58780
rect 65900 58778 65956 58780
rect 65660 58726 65686 58778
rect 65686 58726 65716 58778
rect 65740 58726 65750 58778
rect 65750 58726 65796 58778
rect 65820 58726 65866 58778
rect 65866 58726 65876 58778
rect 65900 58726 65930 58778
rect 65930 58726 65956 58778
rect 65660 58724 65716 58726
rect 65740 58724 65796 58726
rect 65820 58724 65876 58726
rect 65900 58724 65956 58726
rect 65660 57690 65716 57692
rect 65740 57690 65796 57692
rect 65820 57690 65876 57692
rect 65900 57690 65956 57692
rect 65660 57638 65686 57690
rect 65686 57638 65716 57690
rect 65740 57638 65750 57690
rect 65750 57638 65796 57690
rect 65820 57638 65866 57690
rect 65866 57638 65876 57690
rect 65900 57638 65930 57690
rect 65930 57638 65956 57690
rect 65660 57636 65716 57638
rect 65740 57636 65796 57638
rect 65820 57636 65876 57638
rect 65900 57636 65956 57638
rect 65660 56602 65716 56604
rect 65740 56602 65796 56604
rect 65820 56602 65876 56604
rect 65900 56602 65956 56604
rect 65660 56550 65686 56602
rect 65686 56550 65716 56602
rect 65740 56550 65750 56602
rect 65750 56550 65796 56602
rect 65820 56550 65866 56602
rect 65866 56550 65876 56602
rect 65900 56550 65930 56602
rect 65930 56550 65956 56602
rect 65660 56548 65716 56550
rect 65740 56548 65796 56550
rect 65820 56548 65876 56550
rect 65900 56548 65956 56550
rect 65660 55514 65716 55516
rect 65740 55514 65796 55516
rect 65820 55514 65876 55516
rect 65900 55514 65956 55516
rect 65660 55462 65686 55514
rect 65686 55462 65716 55514
rect 65740 55462 65750 55514
rect 65750 55462 65796 55514
rect 65820 55462 65866 55514
rect 65866 55462 65876 55514
rect 65900 55462 65930 55514
rect 65930 55462 65956 55514
rect 65660 55460 65716 55462
rect 65740 55460 65796 55462
rect 65820 55460 65876 55462
rect 65900 55460 65956 55462
rect 65660 54426 65716 54428
rect 65740 54426 65796 54428
rect 65820 54426 65876 54428
rect 65900 54426 65956 54428
rect 65660 54374 65686 54426
rect 65686 54374 65716 54426
rect 65740 54374 65750 54426
rect 65750 54374 65796 54426
rect 65820 54374 65866 54426
rect 65866 54374 65876 54426
rect 65900 54374 65930 54426
rect 65930 54374 65956 54426
rect 65660 54372 65716 54374
rect 65740 54372 65796 54374
rect 65820 54372 65876 54374
rect 65900 54372 65956 54374
rect 65660 53338 65716 53340
rect 65740 53338 65796 53340
rect 65820 53338 65876 53340
rect 65900 53338 65956 53340
rect 65660 53286 65686 53338
rect 65686 53286 65716 53338
rect 65740 53286 65750 53338
rect 65750 53286 65796 53338
rect 65820 53286 65866 53338
rect 65866 53286 65876 53338
rect 65900 53286 65930 53338
rect 65930 53286 65956 53338
rect 65660 53284 65716 53286
rect 65740 53284 65796 53286
rect 65820 53284 65876 53286
rect 65900 53284 65956 53286
rect 65660 52250 65716 52252
rect 65740 52250 65796 52252
rect 65820 52250 65876 52252
rect 65900 52250 65956 52252
rect 65660 52198 65686 52250
rect 65686 52198 65716 52250
rect 65740 52198 65750 52250
rect 65750 52198 65796 52250
rect 65820 52198 65866 52250
rect 65866 52198 65876 52250
rect 65900 52198 65930 52250
rect 65930 52198 65956 52250
rect 65660 52196 65716 52198
rect 65740 52196 65796 52198
rect 65820 52196 65876 52198
rect 65900 52196 65956 52198
rect 65660 51162 65716 51164
rect 65740 51162 65796 51164
rect 65820 51162 65876 51164
rect 65900 51162 65956 51164
rect 65660 51110 65686 51162
rect 65686 51110 65716 51162
rect 65740 51110 65750 51162
rect 65750 51110 65796 51162
rect 65820 51110 65866 51162
rect 65866 51110 65876 51162
rect 65900 51110 65930 51162
rect 65930 51110 65956 51162
rect 65660 51108 65716 51110
rect 65740 51108 65796 51110
rect 65820 51108 65876 51110
rect 65900 51108 65956 51110
rect 65660 50074 65716 50076
rect 65740 50074 65796 50076
rect 65820 50074 65876 50076
rect 65900 50074 65956 50076
rect 65660 50022 65686 50074
rect 65686 50022 65716 50074
rect 65740 50022 65750 50074
rect 65750 50022 65796 50074
rect 65820 50022 65866 50074
rect 65866 50022 65876 50074
rect 65900 50022 65930 50074
rect 65930 50022 65956 50074
rect 65660 50020 65716 50022
rect 65740 50020 65796 50022
rect 65820 50020 65876 50022
rect 65900 50020 65956 50022
rect 65660 48986 65716 48988
rect 65740 48986 65796 48988
rect 65820 48986 65876 48988
rect 65900 48986 65956 48988
rect 65660 48934 65686 48986
rect 65686 48934 65716 48986
rect 65740 48934 65750 48986
rect 65750 48934 65796 48986
rect 65820 48934 65866 48986
rect 65866 48934 65876 48986
rect 65900 48934 65930 48986
rect 65930 48934 65956 48986
rect 65660 48932 65716 48934
rect 65740 48932 65796 48934
rect 65820 48932 65876 48934
rect 65900 48932 65956 48934
rect 65660 47898 65716 47900
rect 65740 47898 65796 47900
rect 65820 47898 65876 47900
rect 65900 47898 65956 47900
rect 65660 47846 65686 47898
rect 65686 47846 65716 47898
rect 65740 47846 65750 47898
rect 65750 47846 65796 47898
rect 65820 47846 65866 47898
rect 65866 47846 65876 47898
rect 65900 47846 65930 47898
rect 65930 47846 65956 47898
rect 65660 47844 65716 47846
rect 65740 47844 65796 47846
rect 65820 47844 65876 47846
rect 65900 47844 65956 47846
rect 65660 46810 65716 46812
rect 65740 46810 65796 46812
rect 65820 46810 65876 46812
rect 65900 46810 65956 46812
rect 65660 46758 65686 46810
rect 65686 46758 65716 46810
rect 65740 46758 65750 46810
rect 65750 46758 65796 46810
rect 65820 46758 65866 46810
rect 65866 46758 65876 46810
rect 65900 46758 65930 46810
rect 65930 46758 65956 46810
rect 65660 46756 65716 46758
rect 65740 46756 65796 46758
rect 65820 46756 65876 46758
rect 65900 46756 65956 46758
rect 65660 45722 65716 45724
rect 65740 45722 65796 45724
rect 65820 45722 65876 45724
rect 65900 45722 65956 45724
rect 65660 45670 65686 45722
rect 65686 45670 65716 45722
rect 65740 45670 65750 45722
rect 65750 45670 65796 45722
rect 65820 45670 65866 45722
rect 65866 45670 65876 45722
rect 65900 45670 65930 45722
rect 65930 45670 65956 45722
rect 65660 45668 65716 45670
rect 65740 45668 65796 45670
rect 65820 45668 65876 45670
rect 65900 45668 65956 45670
rect 65660 44634 65716 44636
rect 65740 44634 65796 44636
rect 65820 44634 65876 44636
rect 65900 44634 65956 44636
rect 65660 44582 65686 44634
rect 65686 44582 65716 44634
rect 65740 44582 65750 44634
rect 65750 44582 65796 44634
rect 65820 44582 65866 44634
rect 65866 44582 65876 44634
rect 65900 44582 65930 44634
rect 65930 44582 65956 44634
rect 65660 44580 65716 44582
rect 65740 44580 65796 44582
rect 65820 44580 65876 44582
rect 65900 44580 65956 44582
rect 65660 43546 65716 43548
rect 65740 43546 65796 43548
rect 65820 43546 65876 43548
rect 65900 43546 65956 43548
rect 65660 43494 65686 43546
rect 65686 43494 65716 43546
rect 65740 43494 65750 43546
rect 65750 43494 65796 43546
rect 65820 43494 65866 43546
rect 65866 43494 65876 43546
rect 65900 43494 65930 43546
rect 65930 43494 65956 43546
rect 65660 43492 65716 43494
rect 65740 43492 65796 43494
rect 65820 43492 65876 43494
rect 65900 43492 65956 43494
rect 65660 42458 65716 42460
rect 65740 42458 65796 42460
rect 65820 42458 65876 42460
rect 65900 42458 65956 42460
rect 65660 42406 65686 42458
rect 65686 42406 65716 42458
rect 65740 42406 65750 42458
rect 65750 42406 65796 42458
rect 65820 42406 65866 42458
rect 65866 42406 65876 42458
rect 65900 42406 65930 42458
rect 65930 42406 65956 42458
rect 65660 42404 65716 42406
rect 65740 42404 65796 42406
rect 65820 42404 65876 42406
rect 65900 42404 65956 42406
rect 65660 41370 65716 41372
rect 65740 41370 65796 41372
rect 65820 41370 65876 41372
rect 65900 41370 65956 41372
rect 65660 41318 65686 41370
rect 65686 41318 65716 41370
rect 65740 41318 65750 41370
rect 65750 41318 65796 41370
rect 65820 41318 65866 41370
rect 65866 41318 65876 41370
rect 65900 41318 65930 41370
rect 65930 41318 65956 41370
rect 65660 41316 65716 41318
rect 65740 41316 65796 41318
rect 65820 41316 65876 41318
rect 65900 41316 65956 41318
rect 65660 40282 65716 40284
rect 65740 40282 65796 40284
rect 65820 40282 65876 40284
rect 65900 40282 65956 40284
rect 65660 40230 65686 40282
rect 65686 40230 65716 40282
rect 65740 40230 65750 40282
rect 65750 40230 65796 40282
rect 65820 40230 65866 40282
rect 65866 40230 65876 40282
rect 65900 40230 65930 40282
rect 65930 40230 65956 40282
rect 65660 40228 65716 40230
rect 65740 40228 65796 40230
rect 65820 40228 65876 40230
rect 65900 40228 65956 40230
rect 65660 39194 65716 39196
rect 65740 39194 65796 39196
rect 65820 39194 65876 39196
rect 65900 39194 65956 39196
rect 65660 39142 65686 39194
rect 65686 39142 65716 39194
rect 65740 39142 65750 39194
rect 65750 39142 65796 39194
rect 65820 39142 65866 39194
rect 65866 39142 65876 39194
rect 65900 39142 65930 39194
rect 65930 39142 65956 39194
rect 65660 39140 65716 39142
rect 65740 39140 65796 39142
rect 65820 39140 65876 39142
rect 65900 39140 65956 39142
rect 65660 38106 65716 38108
rect 65740 38106 65796 38108
rect 65820 38106 65876 38108
rect 65900 38106 65956 38108
rect 65660 38054 65686 38106
rect 65686 38054 65716 38106
rect 65740 38054 65750 38106
rect 65750 38054 65796 38106
rect 65820 38054 65866 38106
rect 65866 38054 65876 38106
rect 65900 38054 65930 38106
rect 65930 38054 65956 38106
rect 65660 38052 65716 38054
rect 65740 38052 65796 38054
rect 65820 38052 65876 38054
rect 65900 38052 65956 38054
rect 65660 37018 65716 37020
rect 65740 37018 65796 37020
rect 65820 37018 65876 37020
rect 65900 37018 65956 37020
rect 65660 36966 65686 37018
rect 65686 36966 65716 37018
rect 65740 36966 65750 37018
rect 65750 36966 65796 37018
rect 65820 36966 65866 37018
rect 65866 36966 65876 37018
rect 65900 36966 65930 37018
rect 65930 36966 65956 37018
rect 65660 36964 65716 36966
rect 65740 36964 65796 36966
rect 65820 36964 65876 36966
rect 65900 36964 65956 36966
rect 65660 35930 65716 35932
rect 65740 35930 65796 35932
rect 65820 35930 65876 35932
rect 65900 35930 65956 35932
rect 65660 35878 65686 35930
rect 65686 35878 65716 35930
rect 65740 35878 65750 35930
rect 65750 35878 65796 35930
rect 65820 35878 65866 35930
rect 65866 35878 65876 35930
rect 65900 35878 65930 35930
rect 65930 35878 65956 35930
rect 65660 35876 65716 35878
rect 65740 35876 65796 35878
rect 65820 35876 65876 35878
rect 65900 35876 65956 35878
rect 65660 34842 65716 34844
rect 65740 34842 65796 34844
rect 65820 34842 65876 34844
rect 65900 34842 65956 34844
rect 65660 34790 65686 34842
rect 65686 34790 65716 34842
rect 65740 34790 65750 34842
rect 65750 34790 65796 34842
rect 65820 34790 65866 34842
rect 65866 34790 65876 34842
rect 65900 34790 65930 34842
rect 65930 34790 65956 34842
rect 65660 34788 65716 34790
rect 65740 34788 65796 34790
rect 65820 34788 65876 34790
rect 65900 34788 65956 34790
rect 65660 33754 65716 33756
rect 65740 33754 65796 33756
rect 65820 33754 65876 33756
rect 65900 33754 65956 33756
rect 65660 33702 65686 33754
rect 65686 33702 65716 33754
rect 65740 33702 65750 33754
rect 65750 33702 65796 33754
rect 65820 33702 65866 33754
rect 65866 33702 65876 33754
rect 65900 33702 65930 33754
rect 65930 33702 65956 33754
rect 65660 33700 65716 33702
rect 65740 33700 65796 33702
rect 65820 33700 65876 33702
rect 65900 33700 65956 33702
rect 65660 32666 65716 32668
rect 65740 32666 65796 32668
rect 65820 32666 65876 32668
rect 65900 32666 65956 32668
rect 65660 32614 65686 32666
rect 65686 32614 65716 32666
rect 65740 32614 65750 32666
rect 65750 32614 65796 32666
rect 65820 32614 65866 32666
rect 65866 32614 65876 32666
rect 65900 32614 65930 32666
rect 65930 32614 65956 32666
rect 65660 32612 65716 32614
rect 65740 32612 65796 32614
rect 65820 32612 65876 32614
rect 65900 32612 65956 32614
rect 65660 31578 65716 31580
rect 65740 31578 65796 31580
rect 65820 31578 65876 31580
rect 65900 31578 65956 31580
rect 65660 31526 65686 31578
rect 65686 31526 65716 31578
rect 65740 31526 65750 31578
rect 65750 31526 65796 31578
rect 65820 31526 65866 31578
rect 65866 31526 65876 31578
rect 65900 31526 65930 31578
rect 65930 31526 65956 31578
rect 65660 31524 65716 31526
rect 65740 31524 65796 31526
rect 65820 31524 65876 31526
rect 65900 31524 65956 31526
rect 65660 30490 65716 30492
rect 65740 30490 65796 30492
rect 65820 30490 65876 30492
rect 65900 30490 65956 30492
rect 65660 30438 65686 30490
rect 65686 30438 65716 30490
rect 65740 30438 65750 30490
rect 65750 30438 65796 30490
rect 65820 30438 65866 30490
rect 65866 30438 65876 30490
rect 65900 30438 65930 30490
rect 65930 30438 65956 30490
rect 65660 30436 65716 30438
rect 65740 30436 65796 30438
rect 65820 30436 65876 30438
rect 65900 30436 65956 30438
rect 65660 29402 65716 29404
rect 65740 29402 65796 29404
rect 65820 29402 65876 29404
rect 65900 29402 65956 29404
rect 65660 29350 65686 29402
rect 65686 29350 65716 29402
rect 65740 29350 65750 29402
rect 65750 29350 65796 29402
rect 65820 29350 65866 29402
rect 65866 29350 65876 29402
rect 65900 29350 65930 29402
rect 65930 29350 65956 29402
rect 65660 29348 65716 29350
rect 65740 29348 65796 29350
rect 65820 29348 65876 29350
rect 65900 29348 65956 29350
rect 65660 28314 65716 28316
rect 65740 28314 65796 28316
rect 65820 28314 65876 28316
rect 65900 28314 65956 28316
rect 65660 28262 65686 28314
rect 65686 28262 65716 28314
rect 65740 28262 65750 28314
rect 65750 28262 65796 28314
rect 65820 28262 65866 28314
rect 65866 28262 65876 28314
rect 65900 28262 65930 28314
rect 65930 28262 65956 28314
rect 65660 28260 65716 28262
rect 65740 28260 65796 28262
rect 65820 28260 65876 28262
rect 65900 28260 65956 28262
rect 65660 27226 65716 27228
rect 65740 27226 65796 27228
rect 65820 27226 65876 27228
rect 65900 27226 65956 27228
rect 65660 27174 65686 27226
rect 65686 27174 65716 27226
rect 65740 27174 65750 27226
rect 65750 27174 65796 27226
rect 65820 27174 65866 27226
rect 65866 27174 65876 27226
rect 65900 27174 65930 27226
rect 65930 27174 65956 27226
rect 65660 27172 65716 27174
rect 65740 27172 65796 27174
rect 65820 27172 65876 27174
rect 65900 27172 65956 27174
rect 65660 26138 65716 26140
rect 65740 26138 65796 26140
rect 65820 26138 65876 26140
rect 65900 26138 65956 26140
rect 65660 26086 65686 26138
rect 65686 26086 65716 26138
rect 65740 26086 65750 26138
rect 65750 26086 65796 26138
rect 65820 26086 65866 26138
rect 65866 26086 65876 26138
rect 65900 26086 65930 26138
rect 65930 26086 65956 26138
rect 65660 26084 65716 26086
rect 65740 26084 65796 26086
rect 65820 26084 65876 26086
rect 65900 26084 65956 26086
rect 65660 25050 65716 25052
rect 65740 25050 65796 25052
rect 65820 25050 65876 25052
rect 65900 25050 65956 25052
rect 65660 24998 65686 25050
rect 65686 24998 65716 25050
rect 65740 24998 65750 25050
rect 65750 24998 65796 25050
rect 65820 24998 65866 25050
rect 65866 24998 65876 25050
rect 65900 24998 65930 25050
rect 65930 24998 65956 25050
rect 65660 24996 65716 24998
rect 65740 24996 65796 24998
rect 65820 24996 65876 24998
rect 65900 24996 65956 24998
rect 65660 23962 65716 23964
rect 65740 23962 65796 23964
rect 65820 23962 65876 23964
rect 65900 23962 65956 23964
rect 65660 23910 65686 23962
rect 65686 23910 65716 23962
rect 65740 23910 65750 23962
rect 65750 23910 65796 23962
rect 65820 23910 65866 23962
rect 65866 23910 65876 23962
rect 65900 23910 65930 23962
rect 65930 23910 65956 23962
rect 65660 23908 65716 23910
rect 65740 23908 65796 23910
rect 65820 23908 65876 23910
rect 65900 23908 65956 23910
rect 65660 22874 65716 22876
rect 65740 22874 65796 22876
rect 65820 22874 65876 22876
rect 65900 22874 65956 22876
rect 65660 22822 65686 22874
rect 65686 22822 65716 22874
rect 65740 22822 65750 22874
rect 65750 22822 65796 22874
rect 65820 22822 65866 22874
rect 65866 22822 65876 22874
rect 65900 22822 65930 22874
rect 65930 22822 65956 22874
rect 65660 22820 65716 22822
rect 65740 22820 65796 22822
rect 65820 22820 65876 22822
rect 65900 22820 65956 22822
rect 65660 21786 65716 21788
rect 65740 21786 65796 21788
rect 65820 21786 65876 21788
rect 65900 21786 65956 21788
rect 65660 21734 65686 21786
rect 65686 21734 65716 21786
rect 65740 21734 65750 21786
rect 65750 21734 65796 21786
rect 65820 21734 65866 21786
rect 65866 21734 65876 21786
rect 65900 21734 65930 21786
rect 65930 21734 65956 21786
rect 65660 21732 65716 21734
rect 65740 21732 65796 21734
rect 65820 21732 65876 21734
rect 65900 21732 65956 21734
rect 65660 20698 65716 20700
rect 65740 20698 65796 20700
rect 65820 20698 65876 20700
rect 65900 20698 65956 20700
rect 65660 20646 65686 20698
rect 65686 20646 65716 20698
rect 65740 20646 65750 20698
rect 65750 20646 65796 20698
rect 65820 20646 65866 20698
rect 65866 20646 65876 20698
rect 65900 20646 65930 20698
rect 65930 20646 65956 20698
rect 65660 20644 65716 20646
rect 65740 20644 65796 20646
rect 65820 20644 65876 20646
rect 65900 20644 65956 20646
rect 65660 19610 65716 19612
rect 65740 19610 65796 19612
rect 65820 19610 65876 19612
rect 65900 19610 65956 19612
rect 65660 19558 65686 19610
rect 65686 19558 65716 19610
rect 65740 19558 65750 19610
rect 65750 19558 65796 19610
rect 65820 19558 65866 19610
rect 65866 19558 65876 19610
rect 65900 19558 65930 19610
rect 65930 19558 65956 19610
rect 65660 19556 65716 19558
rect 65740 19556 65796 19558
rect 65820 19556 65876 19558
rect 65900 19556 65956 19558
rect 65660 18522 65716 18524
rect 65740 18522 65796 18524
rect 65820 18522 65876 18524
rect 65900 18522 65956 18524
rect 65660 18470 65686 18522
rect 65686 18470 65716 18522
rect 65740 18470 65750 18522
rect 65750 18470 65796 18522
rect 65820 18470 65866 18522
rect 65866 18470 65876 18522
rect 65900 18470 65930 18522
rect 65930 18470 65956 18522
rect 65660 18468 65716 18470
rect 65740 18468 65796 18470
rect 65820 18468 65876 18470
rect 65900 18468 65956 18470
rect 65660 17434 65716 17436
rect 65740 17434 65796 17436
rect 65820 17434 65876 17436
rect 65900 17434 65956 17436
rect 65660 17382 65686 17434
rect 65686 17382 65716 17434
rect 65740 17382 65750 17434
rect 65750 17382 65796 17434
rect 65820 17382 65866 17434
rect 65866 17382 65876 17434
rect 65900 17382 65930 17434
rect 65930 17382 65956 17434
rect 65660 17380 65716 17382
rect 65740 17380 65796 17382
rect 65820 17380 65876 17382
rect 65900 17380 65956 17382
rect 66350 63960 66406 64016
rect 66994 63996 66996 64016
rect 66996 63996 67048 64016
rect 67048 63996 67050 64016
rect 66994 63960 67050 63996
rect 65660 16346 65716 16348
rect 65740 16346 65796 16348
rect 65820 16346 65876 16348
rect 65900 16346 65956 16348
rect 65660 16294 65686 16346
rect 65686 16294 65716 16346
rect 65740 16294 65750 16346
rect 65750 16294 65796 16346
rect 65820 16294 65866 16346
rect 65866 16294 65876 16346
rect 65900 16294 65930 16346
rect 65930 16294 65956 16346
rect 65660 16292 65716 16294
rect 65740 16292 65796 16294
rect 65820 16292 65876 16294
rect 65900 16292 65956 16294
rect 65660 15258 65716 15260
rect 65740 15258 65796 15260
rect 65820 15258 65876 15260
rect 65900 15258 65956 15260
rect 65660 15206 65686 15258
rect 65686 15206 65716 15258
rect 65740 15206 65750 15258
rect 65750 15206 65796 15258
rect 65820 15206 65866 15258
rect 65866 15206 65876 15258
rect 65900 15206 65930 15258
rect 65930 15206 65956 15258
rect 65660 15204 65716 15206
rect 65740 15204 65796 15206
rect 65820 15204 65876 15206
rect 65900 15204 65956 15206
rect 65660 14170 65716 14172
rect 65740 14170 65796 14172
rect 65820 14170 65876 14172
rect 65900 14170 65956 14172
rect 65660 14118 65686 14170
rect 65686 14118 65716 14170
rect 65740 14118 65750 14170
rect 65750 14118 65796 14170
rect 65820 14118 65866 14170
rect 65866 14118 65876 14170
rect 65900 14118 65930 14170
rect 65930 14118 65956 14170
rect 65660 14116 65716 14118
rect 65740 14116 65796 14118
rect 65820 14116 65876 14118
rect 65900 14116 65956 14118
rect 65660 13082 65716 13084
rect 65740 13082 65796 13084
rect 65820 13082 65876 13084
rect 65900 13082 65956 13084
rect 65660 13030 65686 13082
rect 65686 13030 65716 13082
rect 65740 13030 65750 13082
rect 65750 13030 65796 13082
rect 65820 13030 65866 13082
rect 65866 13030 65876 13082
rect 65900 13030 65930 13082
rect 65930 13030 65956 13082
rect 65660 13028 65716 13030
rect 65740 13028 65796 13030
rect 65820 13028 65876 13030
rect 65900 13028 65956 13030
rect 65660 11994 65716 11996
rect 65740 11994 65796 11996
rect 65820 11994 65876 11996
rect 65900 11994 65956 11996
rect 65660 11942 65686 11994
rect 65686 11942 65716 11994
rect 65740 11942 65750 11994
rect 65750 11942 65796 11994
rect 65820 11942 65866 11994
rect 65866 11942 65876 11994
rect 65900 11942 65930 11994
rect 65930 11942 65956 11994
rect 65660 11940 65716 11942
rect 65740 11940 65796 11942
rect 65820 11940 65876 11942
rect 65900 11940 65956 11942
rect 65660 10906 65716 10908
rect 65740 10906 65796 10908
rect 65820 10906 65876 10908
rect 65900 10906 65956 10908
rect 65660 10854 65686 10906
rect 65686 10854 65716 10906
rect 65740 10854 65750 10906
rect 65750 10854 65796 10906
rect 65820 10854 65866 10906
rect 65866 10854 65876 10906
rect 65900 10854 65930 10906
rect 65930 10854 65956 10906
rect 65660 10852 65716 10854
rect 65740 10852 65796 10854
rect 65820 10852 65876 10854
rect 65900 10852 65956 10854
rect 65660 9818 65716 9820
rect 65740 9818 65796 9820
rect 65820 9818 65876 9820
rect 65900 9818 65956 9820
rect 65660 9766 65686 9818
rect 65686 9766 65716 9818
rect 65740 9766 65750 9818
rect 65750 9766 65796 9818
rect 65820 9766 65866 9818
rect 65866 9766 65876 9818
rect 65900 9766 65930 9818
rect 65930 9766 65956 9818
rect 65660 9764 65716 9766
rect 65740 9764 65796 9766
rect 65820 9764 65876 9766
rect 65900 9764 65956 9766
rect 65660 8730 65716 8732
rect 65740 8730 65796 8732
rect 65820 8730 65876 8732
rect 65900 8730 65956 8732
rect 65660 8678 65686 8730
rect 65686 8678 65716 8730
rect 65740 8678 65750 8730
rect 65750 8678 65796 8730
rect 65820 8678 65866 8730
rect 65866 8678 65876 8730
rect 65900 8678 65930 8730
rect 65930 8678 65956 8730
rect 65660 8676 65716 8678
rect 65740 8676 65796 8678
rect 65820 8676 65876 8678
rect 65900 8676 65956 8678
rect 65660 7642 65716 7644
rect 65740 7642 65796 7644
rect 65820 7642 65876 7644
rect 65900 7642 65956 7644
rect 65660 7590 65686 7642
rect 65686 7590 65716 7642
rect 65740 7590 65750 7642
rect 65750 7590 65796 7642
rect 65820 7590 65866 7642
rect 65866 7590 65876 7642
rect 65900 7590 65930 7642
rect 65930 7590 65956 7642
rect 65660 7588 65716 7590
rect 65740 7588 65796 7590
rect 65820 7588 65876 7590
rect 65900 7588 65956 7590
rect 65660 6554 65716 6556
rect 65740 6554 65796 6556
rect 65820 6554 65876 6556
rect 65900 6554 65956 6556
rect 65660 6502 65686 6554
rect 65686 6502 65716 6554
rect 65740 6502 65750 6554
rect 65750 6502 65796 6554
rect 65820 6502 65866 6554
rect 65866 6502 65876 6554
rect 65900 6502 65930 6554
rect 65930 6502 65956 6554
rect 65660 6500 65716 6502
rect 65740 6500 65796 6502
rect 65820 6500 65876 6502
rect 65900 6500 65956 6502
rect 65660 5466 65716 5468
rect 65740 5466 65796 5468
rect 65820 5466 65876 5468
rect 65900 5466 65956 5468
rect 65660 5414 65686 5466
rect 65686 5414 65716 5466
rect 65740 5414 65750 5466
rect 65750 5414 65796 5466
rect 65820 5414 65866 5466
rect 65866 5414 65876 5466
rect 65900 5414 65930 5466
rect 65930 5414 65956 5466
rect 65660 5412 65716 5414
rect 65740 5412 65796 5414
rect 65820 5412 65876 5414
rect 65900 5412 65956 5414
rect 65660 4378 65716 4380
rect 65740 4378 65796 4380
rect 65820 4378 65876 4380
rect 65900 4378 65956 4380
rect 65660 4326 65686 4378
rect 65686 4326 65716 4378
rect 65740 4326 65750 4378
rect 65750 4326 65796 4378
rect 65820 4326 65866 4378
rect 65866 4326 65876 4378
rect 65900 4326 65930 4378
rect 65930 4326 65956 4378
rect 65660 4324 65716 4326
rect 65740 4324 65796 4326
rect 65820 4324 65876 4326
rect 65900 4324 65956 4326
rect 65660 3290 65716 3292
rect 65740 3290 65796 3292
rect 65820 3290 65876 3292
rect 65900 3290 65956 3292
rect 65660 3238 65686 3290
rect 65686 3238 65716 3290
rect 65740 3238 65750 3290
rect 65750 3238 65796 3290
rect 65820 3238 65866 3290
rect 65866 3238 65876 3290
rect 65900 3238 65930 3290
rect 65930 3238 65956 3290
rect 65660 3236 65716 3238
rect 65740 3236 65796 3238
rect 65820 3236 65876 3238
rect 65900 3236 65956 3238
rect 65660 2202 65716 2204
rect 65740 2202 65796 2204
rect 65820 2202 65876 2204
rect 65900 2202 65956 2204
rect 65660 2150 65686 2202
rect 65686 2150 65716 2202
rect 65740 2150 65750 2202
rect 65750 2150 65796 2202
rect 65820 2150 65866 2202
rect 65866 2150 65876 2202
rect 65900 2150 65930 2202
rect 65930 2150 65956 2202
rect 65660 2148 65716 2150
rect 65740 2148 65796 2150
rect 65820 2148 65876 2150
rect 65900 2148 65956 2150
rect 67454 63960 67510 64016
rect 67270 63824 67326 63880
rect 67730 18284 67786 18320
rect 67730 18264 67732 18284
rect 67732 18264 67784 18284
rect 67784 18264 67786 18284
rect 70490 18148 70546 18184
rect 70490 18128 70492 18148
rect 70492 18128 70544 18148
rect 70544 18128 70546 18148
rect 71134 18300 71136 18320
rect 71136 18300 71188 18320
rect 71188 18300 71190 18320
rect 71134 18264 71190 18300
rect 71318 18148 71374 18184
rect 71318 18128 71320 18148
rect 71320 18128 71372 18148
rect 71372 18128 71374 18148
rect 81020 97402 81076 97404
rect 81100 97402 81156 97404
rect 81180 97402 81236 97404
rect 81260 97402 81316 97404
rect 81020 97350 81046 97402
rect 81046 97350 81076 97402
rect 81100 97350 81110 97402
rect 81110 97350 81156 97402
rect 81180 97350 81226 97402
rect 81226 97350 81236 97402
rect 81260 97350 81290 97402
rect 81290 97350 81316 97402
rect 81020 97348 81076 97350
rect 81100 97348 81156 97350
rect 81180 97348 81236 97350
rect 81260 97348 81316 97350
rect 81020 96314 81076 96316
rect 81100 96314 81156 96316
rect 81180 96314 81236 96316
rect 81260 96314 81316 96316
rect 81020 96262 81046 96314
rect 81046 96262 81076 96314
rect 81100 96262 81110 96314
rect 81110 96262 81156 96314
rect 81180 96262 81226 96314
rect 81226 96262 81236 96314
rect 81260 96262 81290 96314
rect 81290 96262 81316 96314
rect 81020 96260 81076 96262
rect 81100 96260 81156 96262
rect 81180 96260 81236 96262
rect 81260 96260 81316 96262
rect 81020 95226 81076 95228
rect 81100 95226 81156 95228
rect 81180 95226 81236 95228
rect 81260 95226 81316 95228
rect 81020 95174 81046 95226
rect 81046 95174 81076 95226
rect 81100 95174 81110 95226
rect 81110 95174 81156 95226
rect 81180 95174 81226 95226
rect 81226 95174 81236 95226
rect 81260 95174 81290 95226
rect 81290 95174 81316 95226
rect 81020 95172 81076 95174
rect 81100 95172 81156 95174
rect 81180 95172 81236 95174
rect 81260 95172 81316 95174
rect 81020 94138 81076 94140
rect 81100 94138 81156 94140
rect 81180 94138 81236 94140
rect 81260 94138 81316 94140
rect 81020 94086 81046 94138
rect 81046 94086 81076 94138
rect 81100 94086 81110 94138
rect 81110 94086 81156 94138
rect 81180 94086 81226 94138
rect 81226 94086 81236 94138
rect 81260 94086 81290 94138
rect 81290 94086 81316 94138
rect 81020 94084 81076 94086
rect 81100 94084 81156 94086
rect 81180 94084 81236 94086
rect 81260 94084 81316 94086
rect 81020 93050 81076 93052
rect 81100 93050 81156 93052
rect 81180 93050 81236 93052
rect 81260 93050 81316 93052
rect 81020 92998 81046 93050
rect 81046 92998 81076 93050
rect 81100 92998 81110 93050
rect 81110 92998 81156 93050
rect 81180 92998 81226 93050
rect 81226 92998 81236 93050
rect 81260 92998 81290 93050
rect 81290 92998 81316 93050
rect 81020 92996 81076 92998
rect 81100 92996 81156 92998
rect 81180 92996 81236 92998
rect 81260 92996 81316 92998
rect 81020 91962 81076 91964
rect 81100 91962 81156 91964
rect 81180 91962 81236 91964
rect 81260 91962 81316 91964
rect 81020 91910 81046 91962
rect 81046 91910 81076 91962
rect 81100 91910 81110 91962
rect 81110 91910 81156 91962
rect 81180 91910 81226 91962
rect 81226 91910 81236 91962
rect 81260 91910 81290 91962
rect 81290 91910 81316 91962
rect 81020 91908 81076 91910
rect 81100 91908 81156 91910
rect 81180 91908 81236 91910
rect 81260 91908 81316 91910
rect 81020 90874 81076 90876
rect 81100 90874 81156 90876
rect 81180 90874 81236 90876
rect 81260 90874 81316 90876
rect 81020 90822 81046 90874
rect 81046 90822 81076 90874
rect 81100 90822 81110 90874
rect 81110 90822 81156 90874
rect 81180 90822 81226 90874
rect 81226 90822 81236 90874
rect 81260 90822 81290 90874
rect 81290 90822 81316 90874
rect 81020 90820 81076 90822
rect 81100 90820 81156 90822
rect 81180 90820 81236 90822
rect 81260 90820 81316 90822
rect 81020 89786 81076 89788
rect 81100 89786 81156 89788
rect 81180 89786 81236 89788
rect 81260 89786 81316 89788
rect 81020 89734 81046 89786
rect 81046 89734 81076 89786
rect 81100 89734 81110 89786
rect 81110 89734 81156 89786
rect 81180 89734 81226 89786
rect 81226 89734 81236 89786
rect 81260 89734 81290 89786
rect 81290 89734 81316 89786
rect 81020 89732 81076 89734
rect 81100 89732 81156 89734
rect 81180 89732 81236 89734
rect 81260 89732 81316 89734
rect 81020 88698 81076 88700
rect 81100 88698 81156 88700
rect 81180 88698 81236 88700
rect 81260 88698 81316 88700
rect 81020 88646 81046 88698
rect 81046 88646 81076 88698
rect 81100 88646 81110 88698
rect 81110 88646 81156 88698
rect 81180 88646 81226 88698
rect 81226 88646 81236 88698
rect 81260 88646 81290 88698
rect 81290 88646 81316 88698
rect 81020 88644 81076 88646
rect 81100 88644 81156 88646
rect 81180 88644 81236 88646
rect 81260 88644 81316 88646
rect 81020 87610 81076 87612
rect 81100 87610 81156 87612
rect 81180 87610 81236 87612
rect 81260 87610 81316 87612
rect 81020 87558 81046 87610
rect 81046 87558 81076 87610
rect 81100 87558 81110 87610
rect 81110 87558 81156 87610
rect 81180 87558 81226 87610
rect 81226 87558 81236 87610
rect 81260 87558 81290 87610
rect 81290 87558 81316 87610
rect 81020 87556 81076 87558
rect 81100 87556 81156 87558
rect 81180 87556 81236 87558
rect 81260 87556 81316 87558
rect 81020 86522 81076 86524
rect 81100 86522 81156 86524
rect 81180 86522 81236 86524
rect 81260 86522 81316 86524
rect 81020 86470 81046 86522
rect 81046 86470 81076 86522
rect 81100 86470 81110 86522
rect 81110 86470 81156 86522
rect 81180 86470 81226 86522
rect 81226 86470 81236 86522
rect 81260 86470 81290 86522
rect 81290 86470 81316 86522
rect 81020 86468 81076 86470
rect 81100 86468 81156 86470
rect 81180 86468 81236 86470
rect 81260 86468 81316 86470
rect 81020 85434 81076 85436
rect 81100 85434 81156 85436
rect 81180 85434 81236 85436
rect 81260 85434 81316 85436
rect 81020 85382 81046 85434
rect 81046 85382 81076 85434
rect 81100 85382 81110 85434
rect 81110 85382 81156 85434
rect 81180 85382 81226 85434
rect 81226 85382 81236 85434
rect 81260 85382 81290 85434
rect 81290 85382 81316 85434
rect 81020 85380 81076 85382
rect 81100 85380 81156 85382
rect 81180 85380 81236 85382
rect 81260 85380 81316 85382
rect 81020 84346 81076 84348
rect 81100 84346 81156 84348
rect 81180 84346 81236 84348
rect 81260 84346 81316 84348
rect 81020 84294 81046 84346
rect 81046 84294 81076 84346
rect 81100 84294 81110 84346
rect 81110 84294 81156 84346
rect 81180 84294 81226 84346
rect 81226 84294 81236 84346
rect 81260 84294 81290 84346
rect 81290 84294 81316 84346
rect 81020 84292 81076 84294
rect 81100 84292 81156 84294
rect 81180 84292 81236 84294
rect 81260 84292 81316 84294
rect 81020 83258 81076 83260
rect 81100 83258 81156 83260
rect 81180 83258 81236 83260
rect 81260 83258 81316 83260
rect 81020 83206 81046 83258
rect 81046 83206 81076 83258
rect 81100 83206 81110 83258
rect 81110 83206 81156 83258
rect 81180 83206 81226 83258
rect 81226 83206 81236 83258
rect 81260 83206 81290 83258
rect 81290 83206 81316 83258
rect 81020 83204 81076 83206
rect 81100 83204 81156 83206
rect 81180 83204 81236 83206
rect 81260 83204 81316 83206
rect 81020 82170 81076 82172
rect 81100 82170 81156 82172
rect 81180 82170 81236 82172
rect 81260 82170 81316 82172
rect 81020 82118 81046 82170
rect 81046 82118 81076 82170
rect 81100 82118 81110 82170
rect 81110 82118 81156 82170
rect 81180 82118 81226 82170
rect 81226 82118 81236 82170
rect 81260 82118 81290 82170
rect 81290 82118 81316 82170
rect 81020 82116 81076 82118
rect 81100 82116 81156 82118
rect 81180 82116 81236 82118
rect 81260 82116 81316 82118
rect 81020 81082 81076 81084
rect 81100 81082 81156 81084
rect 81180 81082 81236 81084
rect 81260 81082 81316 81084
rect 81020 81030 81046 81082
rect 81046 81030 81076 81082
rect 81100 81030 81110 81082
rect 81110 81030 81156 81082
rect 81180 81030 81226 81082
rect 81226 81030 81236 81082
rect 81260 81030 81290 81082
rect 81290 81030 81316 81082
rect 81020 81028 81076 81030
rect 81100 81028 81156 81030
rect 81180 81028 81236 81030
rect 81260 81028 81316 81030
rect 81020 79994 81076 79996
rect 81100 79994 81156 79996
rect 81180 79994 81236 79996
rect 81260 79994 81316 79996
rect 81020 79942 81046 79994
rect 81046 79942 81076 79994
rect 81100 79942 81110 79994
rect 81110 79942 81156 79994
rect 81180 79942 81226 79994
rect 81226 79942 81236 79994
rect 81260 79942 81290 79994
rect 81290 79942 81316 79994
rect 81020 79940 81076 79942
rect 81100 79940 81156 79942
rect 81180 79940 81236 79942
rect 81260 79940 81316 79942
rect 81020 78906 81076 78908
rect 81100 78906 81156 78908
rect 81180 78906 81236 78908
rect 81260 78906 81316 78908
rect 81020 78854 81046 78906
rect 81046 78854 81076 78906
rect 81100 78854 81110 78906
rect 81110 78854 81156 78906
rect 81180 78854 81226 78906
rect 81226 78854 81236 78906
rect 81260 78854 81290 78906
rect 81290 78854 81316 78906
rect 81020 78852 81076 78854
rect 81100 78852 81156 78854
rect 81180 78852 81236 78854
rect 81260 78852 81316 78854
rect 81020 77818 81076 77820
rect 81100 77818 81156 77820
rect 81180 77818 81236 77820
rect 81260 77818 81316 77820
rect 81020 77766 81046 77818
rect 81046 77766 81076 77818
rect 81100 77766 81110 77818
rect 81110 77766 81156 77818
rect 81180 77766 81226 77818
rect 81226 77766 81236 77818
rect 81260 77766 81290 77818
rect 81290 77766 81316 77818
rect 81020 77764 81076 77766
rect 81100 77764 81156 77766
rect 81180 77764 81236 77766
rect 81260 77764 81316 77766
rect 81020 76730 81076 76732
rect 81100 76730 81156 76732
rect 81180 76730 81236 76732
rect 81260 76730 81316 76732
rect 81020 76678 81046 76730
rect 81046 76678 81076 76730
rect 81100 76678 81110 76730
rect 81110 76678 81156 76730
rect 81180 76678 81226 76730
rect 81226 76678 81236 76730
rect 81260 76678 81290 76730
rect 81290 76678 81316 76730
rect 81020 76676 81076 76678
rect 81100 76676 81156 76678
rect 81180 76676 81236 76678
rect 81260 76676 81316 76678
rect 81020 75642 81076 75644
rect 81100 75642 81156 75644
rect 81180 75642 81236 75644
rect 81260 75642 81316 75644
rect 81020 75590 81046 75642
rect 81046 75590 81076 75642
rect 81100 75590 81110 75642
rect 81110 75590 81156 75642
rect 81180 75590 81226 75642
rect 81226 75590 81236 75642
rect 81260 75590 81290 75642
rect 81290 75590 81316 75642
rect 81020 75588 81076 75590
rect 81100 75588 81156 75590
rect 81180 75588 81236 75590
rect 81260 75588 81316 75590
rect 81020 74554 81076 74556
rect 81100 74554 81156 74556
rect 81180 74554 81236 74556
rect 81260 74554 81316 74556
rect 81020 74502 81046 74554
rect 81046 74502 81076 74554
rect 81100 74502 81110 74554
rect 81110 74502 81156 74554
rect 81180 74502 81226 74554
rect 81226 74502 81236 74554
rect 81260 74502 81290 74554
rect 81290 74502 81316 74554
rect 81020 74500 81076 74502
rect 81100 74500 81156 74502
rect 81180 74500 81236 74502
rect 81260 74500 81316 74502
rect 81020 73466 81076 73468
rect 81100 73466 81156 73468
rect 81180 73466 81236 73468
rect 81260 73466 81316 73468
rect 81020 73414 81046 73466
rect 81046 73414 81076 73466
rect 81100 73414 81110 73466
rect 81110 73414 81156 73466
rect 81180 73414 81226 73466
rect 81226 73414 81236 73466
rect 81260 73414 81290 73466
rect 81290 73414 81316 73466
rect 81020 73412 81076 73414
rect 81100 73412 81156 73414
rect 81180 73412 81236 73414
rect 81260 73412 81316 73414
rect 81020 72378 81076 72380
rect 81100 72378 81156 72380
rect 81180 72378 81236 72380
rect 81260 72378 81316 72380
rect 81020 72326 81046 72378
rect 81046 72326 81076 72378
rect 81100 72326 81110 72378
rect 81110 72326 81156 72378
rect 81180 72326 81226 72378
rect 81226 72326 81236 72378
rect 81260 72326 81290 72378
rect 81290 72326 81316 72378
rect 81020 72324 81076 72326
rect 81100 72324 81156 72326
rect 81180 72324 81236 72326
rect 81260 72324 81316 72326
rect 81020 71290 81076 71292
rect 81100 71290 81156 71292
rect 81180 71290 81236 71292
rect 81260 71290 81316 71292
rect 81020 71238 81046 71290
rect 81046 71238 81076 71290
rect 81100 71238 81110 71290
rect 81110 71238 81156 71290
rect 81180 71238 81226 71290
rect 81226 71238 81236 71290
rect 81260 71238 81290 71290
rect 81290 71238 81316 71290
rect 81020 71236 81076 71238
rect 81100 71236 81156 71238
rect 81180 71236 81236 71238
rect 81260 71236 81316 71238
rect 81020 70202 81076 70204
rect 81100 70202 81156 70204
rect 81180 70202 81236 70204
rect 81260 70202 81316 70204
rect 81020 70150 81046 70202
rect 81046 70150 81076 70202
rect 81100 70150 81110 70202
rect 81110 70150 81156 70202
rect 81180 70150 81226 70202
rect 81226 70150 81236 70202
rect 81260 70150 81290 70202
rect 81290 70150 81316 70202
rect 81020 70148 81076 70150
rect 81100 70148 81156 70150
rect 81180 70148 81236 70150
rect 81260 70148 81316 70150
rect 81020 69114 81076 69116
rect 81100 69114 81156 69116
rect 81180 69114 81236 69116
rect 81260 69114 81316 69116
rect 81020 69062 81046 69114
rect 81046 69062 81076 69114
rect 81100 69062 81110 69114
rect 81110 69062 81156 69114
rect 81180 69062 81226 69114
rect 81226 69062 81236 69114
rect 81260 69062 81290 69114
rect 81290 69062 81316 69114
rect 81020 69060 81076 69062
rect 81100 69060 81156 69062
rect 81180 69060 81236 69062
rect 81260 69060 81316 69062
rect 81020 68026 81076 68028
rect 81100 68026 81156 68028
rect 81180 68026 81236 68028
rect 81260 68026 81316 68028
rect 81020 67974 81046 68026
rect 81046 67974 81076 68026
rect 81100 67974 81110 68026
rect 81110 67974 81156 68026
rect 81180 67974 81226 68026
rect 81226 67974 81236 68026
rect 81260 67974 81290 68026
rect 81290 67974 81316 68026
rect 81020 67972 81076 67974
rect 81100 67972 81156 67974
rect 81180 67972 81236 67974
rect 81260 67972 81316 67974
rect 81020 66938 81076 66940
rect 81100 66938 81156 66940
rect 81180 66938 81236 66940
rect 81260 66938 81316 66940
rect 81020 66886 81046 66938
rect 81046 66886 81076 66938
rect 81100 66886 81110 66938
rect 81110 66886 81156 66938
rect 81180 66886 81226 66938
rect 81226 66886 81236 66938
rect 81260 66886 81290 66938
rect 81290 66886 81316 66938
rect 81020 66884 81076 66886
rect 81100 66884 81156 66886
rect 81180 66884 81236 66886
rect 81260 66884 81316 66886
rect 81020 65850 81076 65852
rect 81100 65850 81156 65852
rect 81180 65850 81236 65852
rect 81260 65850 81316 65852
rect 81020 65798 81046 65850
rect 81046 65798 81076 65850
rect 81100 65798 81110 65850
rect 81110 65798 81156 65850
rect 81180 65798 81226 65850
rect 81226 65798 81236 65850
rect 81260 65798 81290 65850
rect 81290 65798 81316 65850
rect 81020 65796 81076 65798
rect 81100 65796 81156 65798
rect 81180 65796 81236 65798
rect 81260 65796 81316 65798
rect 81020 64762 81076 64764
rect 81100 64762 81156 64764
rect 81180 64762 81236 64764
rect 81260 64762 81316 64764
rect 81020 64710 81046 64762
rect 81046 64710 81076 64762
rect 81100 64710 81110 64762
rect 81110 64710 81156 64762
rect 81180 64710 81226 64762
rect 81226 64710 81236 64762
rect 81260 64710 81290 64762
rect 81290 64710 81316 64762
rect 81020 64708 81076 64710
rect 81100 64708 81156 64710
rect 81180 64708 81236 64710
rect 81260 64708 81316 64710
rect 81020 63674 81076 63676
rect 81100 63674 81156 63676
rect 81180 63674 81236 63676
rect 81260 63674 81316 63676
rect 81020 63622 81046 63674
rect 81046 63622 81076 63674
rect 81100 63622 81110 63674
rect 81110 63622 81156 63674
rect 81180 63622 81226 63674
rect 81226 63622 81236 63674
rect 81260 63622 81290 63674
rect 81290 63622 81316 63674
rect 81020 63620 81076 63622
rect 81100 63620 81156 63622
rect 81180 63620 81236 63622
rect 81260 63620 81316 63622
rect 81020 62586 81076 62588
rect 81100 62586 81156 62588
rect 81180 62586 81236 62588
rect 81260 62586 81316 62588
rect 81020 62534 81046 62586
rect 81046 62534 81076 62586
rect 81100 62534 81110 62586
rect 81110 62534 81156 62586
rect 81180 62534 81226 62586
rect 81226 62534 81236 62586
rect 81260 62534 81290 62586
rect 81290 62534 81316 62586
rect 81020 62532 81076 62534
rect 81100 62532 81156 62534
rect 81180 62532 81236 62534
rect 81260 62532 81316 62534
rect 81020 61498 81076 61500
rect 81100 61498 81156 61500
rect 81180 61498 81236 61500
rect 81260 61498 81316 61500
rect 81020 61446 81046 61498
rect 81046 61446 81076 61498
rect 81100 61446 81110 61498
rect 81110 61446 81156 61498
rect 81180 61446 81226 61498
rect 81226 61446 81236 61498
rect 81260 61446 81290 61498
rect 81290 61446 81316 61498
rect 81020 61444 81076 61446
rect 81100 61444 81156 61446
rect 81180 61444 81236 61446
rect 81260 61444 81316 61446
rect 81020 60410 81076 60412
rect 81100 60410 81156 60412
rect 81180 60410 81236 60412
rect 81260 60410 81316 60412
rect 81020 60358 81046 60410
rect 81046 60358 81076 60410
rect 81100 60358 81110 60410
rect 81110 60358 81156 60410
rect 81180 60358 81226 60410
rect 81226 60358 81236 60410
rect 81260 60358 81290 60410
rect 81290 60358 81316 60410
rect 81020 60356 81076 60358
rect 81100 60356 81156 60358
rect 81180 60356 81236 60358
rect 81260 60356 81316 60358
rect 81020 59322 81076 59324
rect 81100 59322 81156 59324
rect 81180 59322 81236 59324
rect 81260 59322 81316 59324
rect 81020 59270 81046 59322
rect 81046 59270 81076 59322
rect 81100 59270 81110 59322
rect 81110 59270 81156 59322
rect 81180 59270 81226 59322
rect 81226 59270 81236 59322
rect 81260 59270 81290 59322
rect 81290 59270 81316 59322
rect 81020 59268 81076 59270
rect 81100 59268 81156 59270
rect 81180 59268 81236 59270
rect 81260 59268 81316 59270
rect 81020 58234 81076 58236
rect 81100 58234 81156 58236
rect 81180 58234 81236 58236
rect 81260 58234 81316 58236
rect 81020 58182 81046 58234
rect 81046 58182 81076 58234
rect 81100 58182 81110 58234
rect 81110 58182 81156 58234
rect 81180 58182 81226 58234
rect 81226 58182 81236 58234
rect 81260 58182 81290 58234
rect 81290 58182 81316 58234
rect 81020 58180 81076 58182
rect 81100 58180 81156 58182
rect 81180 58180 81236 58182
rect 81260 58180 81316 58182
rect 81020 57146 81076 57148
rect 81100 57146 81156 57148
rect 81180 57146 81236 57148
rect 81260 57146 81316 57148
rect 81020 57094 81046 57146
rect 81046 57094 81076 57146
rect 81100 57094 81110 57146
rect 81110 57094 81156 57146
rect 81180 57094 81226 57146
rect 81226 57094 81236 57146
rect 81260 57094 81290 57146
rect 81290 57094 81316 57146
rect 81020 57092 81076 57094
rect 81100 57092 81156 57094
rect 81180 57092 81236 57094
rect 81260 57092 81316 57094
rect 81020 56058 81076 56060
rect 81100 56058 81156 56060
rect 81180 56058 81236 56060
rect 81260 56058 81316 56060
rect 81020 56006 81046 56058
rect 81046 56006 81076 56058
rect 81100 56006 81110 56058
rect 81110 56006 81156 56058
rect 81180 56006 81226 56058
rect 81226 56006 81236 56058
rect 81260 56006 81290 56058
rect 81290 56006 81316 56058
rect 81020 56004 81076 56006
rect 81100 56004 81156 56006
rect 81180 56004 81236 56006
rect 81260 56004 81316 56006
rect 81020 54970 81076 54972
rect 81100 54970 81156 54972
rect 81180 54970 81236 54972
rect 81260 54970 81316 54972
rect 81020 54918 81046 54970
rect 81046 54918 81076 54970
rect 81100 54918 81110 54970
rect 81110 54918 81156 54970
rect 81180 54918 81226 54970
rect 81226 54918 81236 54970
rect 81260 54918 81290 54970
rect 81290 54918 81316 54970
rect 81020 54916 81076 54918
rect 81100 54916 81156 54918
rect 81180 54916 81236 54918
rect 81260 54916 81316 54918
rect 81020 53882 81076 53884
rect 81100 53882 81156 53884
rect 81180 53882 81236 53884
rect 81260 53882 81316 53884
rect 81020 53830 81046 53882
rect 81046 53830 81076 53882
rect 81100 53830 81110 53882
rect 81110 53830 81156 53882
rect 81180 53830 81226 53882
rect 81226 53830 81236 53882
rect 81260 53830 81290 53882
rect 81290 53830 81316 53882
rect 81020 53828 81076 53830
rect 81100 53828 81156 53830
rect 81180 53828 81236 53830
rect 81260 53828 81316 53830
rect 81020 52794 81076 52796
rect 81100 52794 81156 52796
rect 81180 52794 81236 52796
rect 81260 52794 81316 52796
rect 81020 52742 81046 52794
rect 81046 52742 81076 52794
rect 81100 52742 81110 52794
rect 81110 52742 81156 52794
rect 81180 52742 81226 52794
rect 81226 52742 81236 52794
rect 81260 52742 81290 52794
rect 81290 52742 81316 52794
rect 81020 52740 81076 52742
rect 81100 52740 81156 52742
rect 81180 52740 81236 52742
rect 81260 52740 81316 52742
rect 81020 51706 81076 51708
rect 81100 51706 81156 51708
rect 81180 51706 81236 51708
rect 81260 51706 81316 51708
rect 81020 51654 81046 51706
rect 81046 51654 81076 51706
rect 81100 51654 81110 51706
rect 81110 51654 81156 51706
rect 81180 51654 81226 51706
rect 81226 51654 81236 51706
rect 81260 51654 81290 51706
rect 81290 51654 81316 51706
rect 81020 51652 81076 51654
rect 81100 51652 81156 51654
rect 81180 51652 81236 51654
rect 81260 51652 81316 51654
rect 81020 50618 81076 50620
rect 81100 50618 81156 50620
rect 81180 50618 81236 50620
rect 81260 50618 81316 50620
rect 81020 50566 81046 50618
rect 81046 50566 81076 50618
rect 81100 50566 81110 50618
rect 81110 50566 81156 50618
rect 81180 50566 81226 50618
rect 81226 50566 81236 50618
rect 81260 50566 81290 50618
rect 81290 50566 81316 50618
rect 81020 50564 81076 50566
rect 81100 50564 81156 50566
rect 81180 50564 81236 50566
rect 81260 50564 81316 50566
rect 81020 49530 81076 49532
rect 81100 49530 81156 49532
rect 81180 49530 81236 49532
rect 81260 49530 81316 49532
rect 81020 49478 81046 49530
rect 81046 49478 81076 49530
rect 81100 49478 81110 49530
rect 81110 49478 81156 49530
rect 81180 49478 81226 49530
rect 81226 49478 81236 49530
rect 81260 49478 81290 49530
rect 81290 49478 81316 49530
rect 81020 49476 81076 49478
rect 81100 49476 81156 49478
rect 81180 49476 81236 49478
rect 81260 49476 81316 49478
rect 81020 48442 81076 48444
rect 81100 48442 81156 48444
rect 81180 48442 81236 48444
rect 81260 48442 81316 48444
rect 81020 48390 81046 48442
rect 81046 48390 81076 48442
rect 81100 48390 81110 48442
rect 81110 48390 81156 48442
rect 81180 48390 81226 48442
rect 81226 48390 81236 48442
rect 81260 48390 81290 48442
rect 81290 48390 81316 48442
rect 81020 48388 81076 48390
rect 81100 48388 81156 48390
rect 81180 48388 81236 48390
rect 81260 48388 81316 48390
rect 81020 47354 81076 47356
rect 81100 47354 81156 47356
rect 81180 47354 81236 47356
rect 81260 47354 81316 47356
rect 81020 47302 81046 47354
rect 81046 47302 81076 47354
rect 81100 47302 81110 47354
rect 81110 47302 81156 47354
rect 81180 47302 81226 47354
rect 81226 47302 81236 47354
rect 81260 47302 81290 47354
rect 81290 47302 81316 47354
rect 81020 47300 81076 47302
rect 81100 47300 81156 47302
rect 81180 47300 81236 47302
rect 81260 47300 81316 47302
rect 81020 46266 81076 46268
rect 81100 46266 81156 46268
rect 81180 46266 81236 46268
rect 81260 46266 81316 46268
rect 81020 46214 81046 46266
rect 81046 46214 81076 46266
rect 81100 46214 81110 46266
rect 81110 46214 81156 46266
rect 81180 46214 81226 46266
rect 81226 46214 81236 46266
rect 81260 46214 81290 46266
rect 81290 46214 81316 46266
rect 81020 46212 81076 46214
rect 81100 46212 81156 46214
rect 81180 46212 81236 46214
rect 81260 46212 81316 46214
rect 81020 45178 81076 45180
rect 81100 45178 81156 45180
rect 81180 45178 81236 45180
rect 81260 45178 81316 45180
rect 81020 45126 81046 45178
rect 81046 45126 81076 45178
rect 81100 45126 81110 45178
rect 81110 45126 81156 45178
rect 81180 45126 81226 45178
rect 81226 45126 81236 45178
rect 81260 45126 81290 45178
rect 81290 45126 81316 45178
rect 81020 45124 81076 45126
rect 81100 45124 81156 45126
rect 81180 45124 81236 45126
rect 81260 45124 81316 45126
rect 81020 44090 81076 44092
rect 81100 44090 81156 44092
rect 81180 44090 81236 44092
rect 81260 44090 81316 44092
rect 81020 44038 81046 44090
rect 81046 44038 81076 44090
rect 81100 44038 81110 44090
rect 81110 44038 81156 44090
rect 81180 44038 81226 44090
rect 81226 44038 81236 44090
rect 81260 44038 81290 44090
rect 81290 44038 81316 44090
rect 81020 44036 81076 44038
rect 81100 44036 81156 44038
rect 81180 44036 81236 44038
rect 81260 44036 81316 44038
rect 81020 43002 81076 43004
rect 81100 43002 81156 43004
rect 81180 43002 81236 43004
rect 81260 43002 81316 43004
rect 81020 42950 81046 43002
rect 81046 42950 81076 43002
rect 81100 42950 81110 43002
rect 81110 42950 81156 43002
rect 81180 42950 81226 43002
rect 81226 42950 81236 43002
rect 81260 42950 81290 43002
rect 81290 42950 81316 43002
rect 81020 42948 81076 42950
rect 81100 42948 81156 42950
rect 81180 42948 81236 42950
rect 81260 42948 81316 42950
rect 81020 41914 81076 41916
rect 81100 41914 81156 41916
rect 81180 41914 81236 41916
rect 81260 41914 81316 41916
rect 81020 41862 81046 41914
rect 81046 41862 81076 41914
rect 81100 41862 81110 41914
rect 81110 41862 81156 41914
rect 81180 41862 81226 41914
rect 81226 41862 81236 41914
rect 81260 41862 81290 41914
rect 81290 41862 81316 41914
rect 81020 41860 81076 41862
rect 81100 41860 81156 41862
rect 81180 41860 81236 41862
rect 81260 41860 81316 41862
rect 81020 40826 81076 40828
rect 81100 40826 81156 40828
rect 81180 40826 81236 40828
rect 81260 40826 81316 40828
rect 81020 40774 81046 40826
rect 81046 40774 81076 40826
rect 81100 40774 81110 40826
rect 81110 40774 81156 40826
rect 81180 40774 81226 40826
rect 81226 40774 81236 40826
rect 81260 40774 81290 40826
rect 81290 40774 81316 40826
rect 81020 40772 81076 40774
rect 81100 40772 81156 40774
rect 81180 40772 81236 40774
rect 81260 40772 81316 40774
rect 81020 39738 81076 39740
rect 81100 39738 81156 39740
rect 81180 39738 81236 39740
rect 81260 39738 81316 39740
rect 81020 39686 81046 39738
rect 81046 39686 81076 39738
rect 81100 39686 81110 39738
rect 81110 39686 81156 39738
rect 81180 39686 81226 39738
rect 81226 39686 81236 39738
rect 81260 39686 81290 39738
rect 81290 39686 81316 39738
rect 81020 39684 81076 39686
rect 81100 39684 81156 39686
rect 81180 39684 81236 39686
rect 81260 39684 81316 39686
rect 81020 38650 81076 38652
rect 81100 38650 81156 38652
rect 81180 38650 81236 38652
rect 81260 38650 81316 38652
rect 81020 38598 81046 38650
rect 81046 38598 81076 38650
rect 81100 38598 81110 38650
rect 81110 38598 81156 38650
rect 81180 38598 81226 38650
rect 81226 38598 81236 38650
rect 81260 38598 81290 38650
rect 81290 38598 81316 38650
rect 81020 38596 81076 38598
rect 81100 38596 81156 38598
rect 81180 38596 81236 38598
rect 81260 38596 81316 38598
rect 81020 37562 81076 37564
rect 81100 37562 81156 37564
rect 81180 37562 81236 37564
rect 81260 37562 81316 37564
rect 81020 37510 81046 37562
rect 81046 37510 81076 37562
rect 81100 37510 81110 37562
rect 81110 37510 81156 37562
rect 81180 37510 81226 37562
rect 81226 37510 81236 37562
rect 81260 37510 81290 37562
rect 81290 37510 81316 37562
rect 81020 37508 81076 37510
rect 81100 37508 81156 37510
rect 81180 37508 81236 37510
rect 81260 37508 81316 37510
rect 81020 36474 81076 36476
rect 81100 36474 81156 36476
rect 81180 36474 81236 36476
rect 81260 36474 81316 36476
rect 81020 36422 81046 36474
rect 81046 36422 81076 36474
rect 81100 36422 81110 36474
rect 81110 36422 81156 36474
rect 81180 36422 81226 36474
rect 81226 36422 81236 36474
rect 81260 36422 81290 36474
rect 81290 36422 81316 36474
rect 81020 36420 81076 36422
rect 81100 36420 81156 36422
rect 81180 36420 81236 36422
rect 81260 36420 81316 36422
rect 81020 35386 81076 35388
rect 81100 35386 81156 35388
rect 81180 35386 81236 35388
rect 81260 35386 81316 35388
rect 81020 35334 81046 35386
rect 81046 35334 81076 35386
rect 81100 35334 81110 35386
rect 81110 35334 81156 35386
rect 81180 35334 81226 35386
rect 81226 35334 81236 35386
rect 81260 35334 81290 35386
rect 81290 35334 81316 35386
rect 81020 35332 81076 35334
rect 81100 35332 81156 35334
rect 81180 35332 81236 35334
rect 81260 35332 81316 35334
rect 81020 34298 81076 34300
rect 81100 34298 81156 34300
rect 81180 34298 81236 34300
rect 81260 34298 81316 34300
rect 81020 34246 81046 34298
rect 81046 34246 81076 34298
rect 81100 34246 81110 34298
rect 81110 34246 81156 34298
rect 81180 34246 81226 34298
rect 81226 34246 81236 34298
rect 81260 34246 81290 34298
rect 81290 34246 81316 34298
rect 81020 34244 81076 34246
rect 81100 34244 81156 34246
rect 81180 34244 81236 34246
rect 81260 34244 81316 34246
rect 81020 33210 81076 33212
rect 81100 33210 81156 33212
rect 81180 33210 81236 33212
rect 81260 33210 81316 33212
rect 81020 33158 81046 33210
rect 81046 33158 81076 33210
rect 81100 33158 81110 33210
rect 81110 33158 81156 33210
rect 81180 33158 81226 33210
rect 81226 33158 81236 33210
rect 81260 33158 81290 33210
rect 81290 33158 81316 33210
rect 81020 33156 81076 33158
rect 81100 33156 81156 33158
rect 81180 33156 81236 33158
rect 81260 33156 81316 33158
rect 81020 32122 81076 32124
rect 81100 32122 81156 32124
rect 81180 32122 81236 32124
rect 81260 32122 81316 32124
rect 81020 32070 81046 32122
rect 81046 32070 81076 32122
rect 81100 32070 81110 32122
rect 81110 32070 81156 32122
rect 81180 32070 81226 32122
rect 81226 32070 81236 32122
rect 81260 32070 81290 32122
rect 81290 32070 81316 32122
rect 81020 32068 81076 32070
rect 81100 32068 81156 32070
rect 81180 32068 81236 32070
rect 81260 32068 81316 32070
rect 81020 31034 81076 31036
rect 81100 31034 81156 31036
rect 81180 31034 81236 31036
rect 81260 31034 81316 31036
rect 81020 30982 81046 31034
rect 81046 30982 81076 31034
rect 81100 30982 81110 31034
rect 81110 30982 81156 31034
rect 81180 30982 81226 31034
rect 81226 30982 81236 31034
rect 81260 30982 81290 31034
rect 81290 30982 81316 31034
rect 81020 30980 81076 30982
rect 81100 30980 81156 30982
rect 81180 30980 81236 30982
rect 81260 30980 81316 30982
rect 81020 29946 81076 29948
rect 81100 29946 81156 29948
rect 81180 29946 81236 29948
rect 81260 29946 81316 29948
rect 81020 29894 81046 29946
rect 81046 29894 81076 29946
rect 81100 29894 81110 29946
rect 81110 29894 81156 29946
rect 81180 29894 81226 29946
rect 81226 29894 81236 29946
rect 81260 29894 81290 29946
rect 81290 29894 81316 29946
rect 81020 29892 81076 29894
rect 81100 29892 81156 29894
rect 81180 29892 81236 29894
rect 81260 29892 81316 29894
rect 81020 28858 81076 28860
rect 81100 28858 81156 28860
rect 81180 28858 81236 28860
rect 81260 28858 81316 28860
rect 81020 28806 81046 28858
rect 81046 28806 81076 28858
rect 81100 28806 81110 28858
rect 81110 28806 81156 28858
rect 81180 28806 81226 28858
rect 81226 28806 81236 28858
rect 81260 28806 81290 28858
rect 81290 28806 81316 28858
rect 81020 28804 81076 28806
rect 81100 28804 81156 28806
rect 81180 28804 81236 28806
rect 81260 28804 81316 28806
rect 81020 27770 81076 27772
rect 81100 27770 81156 27772
rect 81180 27770 81236 27772
rect 81260 27770 81316 27772
rect 81020 27718 81046 27770
rect 81046 27718 81076 27770
rect 81100 27718 81110 27770
rect 81110 27718 81156 27770
rect 81180 27718 81226 27770
rect 81226 27718 81236 27770
rect 81260 27718 81290 27770
rect 81290 27718 81316 27770
rect 81020 27716 81076 27718
rect 81100 27716 81156 27718
rect 81180 27716 81236 27718
rect 81260 27716 81316 27718
rect 81020 26682 81076 26684
rect 81100 26682 81156 26684
rect 81180 26682 81236 26684
rect 81260 26682 81316 26684
rect 81020 26630 81046 26682
rect 81046 26630 81076 26682
rect 81100 26630 81110 26682
rect 81110 26630 81156 26682
rect 81180 26630 81226 26682
rect 81226 26630 81236 26682
rect 81260 26630 81290 26682
rect 81290 26630 81316 26682
rect 81020 26628 81076 26630
rect 81100 26628 81156 26630
rect 81180 26628 81236 26630
rect 81260 26628 81316 26630
rect 81020 25594 81076 25596
rect 81100 25594 81156 25596
rect 81180 25594 81236 25596
rect 81260 25594 81316 25596
rect 81020 25542 81046 25594
rect 81046 25542 81076 25594
rect 81100 25542 81110 25594
rect 81110 25542 81156 25594
rect 81180 25542 81226 25594
rect 81226 25542 81236 25594
rect 81260 25542 81290 25594
rect 81290 25542 81316 25594
rect 81020 25540 81076 25542
rect 81100 25540 81156 25542
rect 81180 25540 81236 25542
rect 81260 25540 81316 25542
rect 81020 24506 81076 24508
rect 81100 24506 81156 24508
rect 81180 24506 81236 24508
rect 81260 24506 81316 24508
rect 81020 24454 81046 24506
rect 81046 24454 81076 24506
rect 81100 24454 81110 24506
rect 81110 24454 81156 24506
rect 81180 24454 81226 24506
rect 81226 24454 81236 24506
rect 81260 24454 81290 24506
rect 81290 24454 81316 24506
rect 81020 24452 81076 24454
rect 81100 24452 81156 24454
rect 81180 24452 81236 24454
rect 81260 24452 81316 24454
rect 81020 23418 81076 23420
rect 81100 23418 81156 23420
rect 81180 23418 81236 23420
rect 81260 23418 81316 23420
rect 81020 23366 81046 23418
rect 81046 23366 81076 23418
rect 81100 23366 81110 23418
rect 81110 23366 81156 23418
rect 81180 23366 81226 23418
rect 81226 23366 81236 23418
rect 81260 23366 81290 23418
rect 81290 23366 81316 23418
rect 81020 23364 81076 23366
rect 81100 23364 81156 23366
rect 81180 23364 81236 23366
rect 81260 23364 81316 23366
rect 81020 22330 81076 22332
rect 81100 22330 81156 22332
rect 81180 22330 81236 22332
rect 81260 22330 81316 22332
rect 81020 22278 81046 22330
rect 81046 22278 81076 22330
rect 81100 22278 81110 22330
rect 81110 22278 81156 22330
rect 81180 22278 81226 22330
rect 81226 22278 81236 22330
rect 81260 22278 81290 22330
rect 81290 22278 81316 22330
rect 81020 22276 81076 22278
rect 81100 22276 81156 22278
rect 81180 22276 81236 22278
rect 81260 22276 81316 22278
rect 81020 21242 81076 21244
rect 81100 21242 81156 21244
rect 81180 21242 81236 21244
rect 81260 21242 81316 21244
rect 81020 21190 81046 21242
rect 81046 21190 81076 21242
rect 81100 21190 81110 21242
rect 81110 21190 81156 21242
rect 81180 21190 81226 21242
rect 81226 21190 81236 21242
rect 81260 21190 81290 21242
rect 81290 21190 81316 21242
rect 81020 21188 81076 21190
rect 81100 21188 81156 21190
rect 81180 21188 81236 21190
rect 81260 21188 81316 21190
rect 81020 20154 81076 20156
rect 81100 20154 81156 20156
rect 81180 20154 81236 20156
rect 81260 20154 81316 20156
rect 81020 20102 81046 20154
rect 81046 20102 81076 20154
rect 81100 20102 81110 20154
rect 81110 20102 81156 20154
rect 81180 20102 81226 20154
rect 81226 20102 81236 20154
rect 81260 20102 81290 20154
rect 81290 20102 81316 20154
rect 81020 20100 81076 20102
rect 81100 20100 81156 20102
rect 81180 20100 81236 20102
rect 81260 20100 81316 20102
rect 81020 19066 81076 19068
rect 81100 19066 81156 19068
rect 81180 19066 81236 19068
rect 81260 19066 81316 19068
rect 81020 19014 81046 19066
rect 81046 19014 81076 19066
rect 81100 19014 81110 19066
rect 81110 19014 81156 19066
rect 81180 19014 81226 19066
rect 81226 19014 81236 19066
rect 81260 19014 81290 19066
rect 81290 19014 81316 19066
rect 81020 19012 81076 19014
rect 81100 19012 81156 19014
rect 81180 19012 81236 19014
rect 81260 19012 81316 19014
rect 81020 17978 81076 17980
rect 81100 17978 81156 17980
rect 81180 17978 81236 17980
rect 81260 17978 81316 17980
rect 81020 17926 81046 17978
rect 81046 17926 81076 17978
rect 81100 17926 81110 17978
rect 81110 17926 81156 17978
rect 81180 17926 81226 17978
rect 81226 17926 81236 17978
rect 81260 17926 81290 17978
rect 81290 17926 81316 17978
rect 81020 17924 81076 17926
rect 81100 17924 81156 17926
rect 81180 17924 81236 17926
rect 81260 17924 81316 17926
rect 81020 16890 81076 16892
rect 81100 16890 81156 16892
rect 81180 16890 81236 16892
rect 81260 16890 81316 16892
rect 81020 16838 81046 16890
rect 81046 16838 81076 16890
rect 81100 16838 81110 16890
rect 81110 16838 81156 16890
rect 81180 16838 81226 16890
rect 81226 16838 81236 16890
rect 81260 16838 81290 16890
rect 81290 16838 81316 16890
rect 81020 16836 81076 16838
rect 81100 16836 81156 16838
rect 81180 16836 81236 16838
rect 81260 16836 81316 16838
rect 81020 15802 81076 15804
rect 81100 15802 81156 15804
rect 81180 15802 81236 15804
rect 81260 15802 81316 15804
rect 81020 15750 81046 15802
rect 81046 15750 81076 15802
rect 81100 15750 81110 15802
rect 81110 15750 81156 15802
rect 81180 15750 81226 15802
rect 81226 15750 81236 15802
rect 81260 15750 81290 15802
rect 81290 15750 81316 15802
rect 81020 15748 81076 15750
rect 81100 15748 81156 15750
rect 81180 15748 81236 15750
rect 81260 15748 81316 15750
rect 81020 14714 81076 14716
rect 81100 14714 81156 14716
rect 81180 14714 81236 14716
rect 81260 14714 81316 14716
rect 81020 14662 81046 14714
rect 81046 14662 81076 14714
rect 81100 14662 81110 14714
rect 81110 14662 81156 14714
rect 81180 14662 81226 14714
rect 81226 14662 81236 14714
rect 81260 14662 81290 14714
rect 81290 14662 81316 14714
rect 81020 14660 81076 14662
rect 81100 14660 81156 14662
rect 81180 14660 81236 14662
rect 81260 14660 81316 14662
rect 81020 13626 81076 13628
rect 81100 13626 81156 13628
rect 81180 13626 81236 13628
rect 81260 13626 81316 13628
rect 81020 13574 81046 13626
rect 81046 13574 81076 13626
rect 81100 13574 81110 13626
rect 81110 13574 81156 13626
rect 81180 13574 81226 13626
rect 81226 13574 81236 13626
rect 81260 13574 81290 13626
rect 81290 13574 81316 13626
rect 81020 13572 81076 13574
rect 81100 13572 81156 13574
rect 81180 13572 81236 13574
rect 81260 13572 81316 13574
rect 81020 12538 81076 12540
rect 81100 12538 81156 12540
rect 81180 12538 81236 12540
rect 81260 12538 81316 12540
rect 81020 12486 81046 12538
rect 81046 12486 81076 12538
rect 81100 12486 81110 12538
rect 81110 12486 81156 12538
rect 81180 12486 81226 12538
rect 81226 12486 81236 12538
rect 81260 12486 81290 12538
rect 81290 12486 81316 12538
rect 81020 12484 81076 12486
rect 81100 12484 81156 12486
rect 81180 12484 81236 12486
rect 81260 12484 81316 12486
rect 81020 11450 81076 11452
rect 81100 11450 81156 11452
rect 81180 11450 81236 11452
rect 81260 11450 81316 11452
rect 81020 11398 81046 11450
rect 81046 11398 81076 11450
rect 81100 11398 81110 11450
rect 81110 11398 81156 11450
rect 81180 11398 81226 11450
rect 81226 11398 81236 11450
rect 81260 11398 81290 11450
rect 81290 11398 81316 11450
rect 81020 11396 81076 11398
rect 81100 11396 81156 11398
rect 81180 11396 81236 11398
rect 81260 11396 81316 11398
rect 81020 10362 81076 10364
rect 81100 10362 81156 10364
rect 81180 10362 81236 10364
rect 81260 10362 81316 10364
rect 81020 10310 81046 10362
rect 81046 10310 81076 10362
rect 81100 10310 81110 10362
rect 81110 10310 81156 10362
rect 81180 10310 81226 10362
rect 81226 10310 81236 10362
rect 81260 10310 81290 10362
rect 81290 10310 81316 10362
rect 81020 10308 81076 10310
rect 81100 10308 81156 10310
rect 81180 10308 81236 10310
rect 81260 10308 81316 10310
rect 81020 9274 81076 9276
rect 81100 9274 81156 9276
rect 81180 9274 81236 9276
rect 81260 9274 81316 9276
rect 81020 9222 81046 9274
rect 81046 9222 81076 9274
rect 81100 9222 81110 9274
rect 81110 9222 81156 9274
rect 81180 9222 81226 9274
rect 81226 9222 81236 9274
rect 81260 9222 81290 9274
rect 81290 9222 81316 9274
rect 81020 9220 81076 9222
rect 81100 9220 81156 9222
rect 81180 9220 81236 9222
rect 81260 9220 81316 9222
rect 81020 8186 81076 8188
rect 81100 8186 81156 8188
rect 81180 8186 81236 8188
rect 81260 8186 81316 8188
rect 81020 8134 81046 8186
rect 81046 8134 81076 8186
rect 81100 8134 81110 8186
rect 81110 8134 81156 8186
rect 81180 8134 81226 8186
rect 81226 8134 81236 8186
rect 81260 8134 81290 8186
rect 81290 8134 81316 8186
rect 81020 8132 81076 8134
rect 81100 8132 81156 8134
rect 81180 8132 81236 8134
rect 81260 8132 81316 8134
rect 81020 7098 81076 7100
rect 81100 7098 81156 7100
rect 81180 7098 81236 7100
rect 81260 7098 81316 7100
rect 81020 7046 81046 7098
rect 81046 7046 81076 7098
rect 81100 7046 81110 7098
rect 81110 7046 81156 7098
rect 81180 7046 81226 7098
rect 81226 7046 81236 7098
rect 81260 7046 81290 7098
rect 81290 7046 81316 7098
rect 81020 7044 81076 7046
rect 81100 7044 81156 7046
rect 81180 7044 81236 7046
rect 81260 7044 81316 7046
rect 81020 6010 81076 6012
rect 81100 6010 81156 6012
rect 81180 6010 81236 6012
rect 81260 6010 81316 6012
rect 81020 5958 81046 6010
rect 81046 5958 81076 6010
rect 81100 5958 81110 6010
rect 81110 5958 81156 6010
rect 81180 5958 81226 6010
rect 81226 5958 81236 6010
rect 81260 5958 81290 6010
rect 81290 5958 81316 6010
rect 81020 5956 81076 5958
rect 81100 5956 81156 5958
rect 81180 5956 81236 5958
rect 81260 5956 81316 5958
rect 81020 4922 81076 4924
rect 81100 4922 81156 4924
rect 81180 4922 81236 4924
rect 81260 4922 81316 4924
rect 81020 4870 81046 4922
rect 81046 4870 81076 4922
rect 81100 4870 81110 4922
rect 81110 4870 81156 4922
rect 81180 4870 81226 4922
rect 81226 4870 81236 4922
rect 81260 4870 81290 4922
rect 81290 4870 81316 4922
rect 81020 4868 81076 4870
rect 81100 4868 81156 4870
rect 81180 4868 81236 4870
rect 81260 4868 81316 4870
rect 81020 3834 81076 3836
rect 81100 3834 81156 3836
rect 81180 3834 81236 3836
rect 81260 3834 81316 3836
rect 81020 3782 81046 3834
rect 81046 3782 81076 3834
rect 81100 3782 81110 3834
rect 81110 3782 81156 3834
rect 81180 3782 81226 3834
rect 81226 3782 81236 3834
rect 81260 3782 81290 3834
rect 81290 3782 81316 3834
rect 81020 3780 81076 3782
rect 81100 3780 81156 3782
rect 81180 3780 81236 3782
rect 81260 3780 81316 3782
rect 81020 2746 81076 2748
rect 81100 2746 81156 2748
rect 81180 2746 81236 2748
rect 81260 2746 81316 2748
rect 81020 2694 81046 2746
rect 81046 2694 81076 2746
rect 81100 2694 81110 2746
rect 81110 2694 81156 2746
rect 81180 2694 81226 2746
rect 81226 2694 81236 2746
rect 81260 2694 81290 2746
rect 81290 2694 81316 2746
rect 81020 2692 81076 2694
rect 81100 2692 81156 2694
rect 81180 2692 81236 2694
rect 81260 2692 81316 2694
rect 96380 96858 96436 96860
rect 96460 96858 96516 96860
rect 96540 96858 96596 96860
rect 96620 96858 96676 96860
rect 96380 96806 96406 96858
rect 96406 96806 96436 96858
rect 96460 96806 96470 96858
rect 96470 96806 96516 96858
rect 96540 96806 96586 96858
rect 96586 96806 96596 96858
rect 96620 96806 96650 96858
rect 96650 96806 96676 96858
rect 96380 96804 96436 96806
rect 96460 96804 96516 96806
rect 96540 96804 96596 96806
rect 96620 96804 96676 96806
rect 96380 95770 96436 95772
rect 96460 95770 96516 95772
rect 96540 95770 96596 95772
rect 96620 95770 96676 95772
rect 96380 95718 96406 95770
rect 96406 95718 96436 95770
rect 96460 95718 96470 95770
rect 96470 95718 96516 95770
rect 96540 95718 96586 95770
rect 96586 95718 96596 95770
rect 96620 95718 96650 95770
rect 96650 95718 96676 95770
rect 96380 95716 96436 95718
rect 96460 95716 96516 95718
rect 96540 95716 96596 95718
rect 96620 95716 96676 95718
rect 96380 94682 96436 94684
rect 96460 94682 96516 94684
rect 96540 94682 96596 94684
rect 96620 94682 96676 94684
rect 96380 94630 96406 94682
rect 96406 94630 96436 94682
rect 96460 94630 96470 94682
rect 96470 94630 96516 94682
rect 96540 94630 96586 94682
rect 96586 94630 96596 94682
rect 96620 94630 96650 94682
rect 96650 94630 96676 94682
rect 96380 94628 96436 94630
rect 96460 94628 96516 94630
rect 96540 94628 96596 94630
rect 96620 94628 96676 94630
rect 96380 93594 96436 93596
rect 96460 93594 96516 93596
rect 96540 93594 96596 93596
rect 96620 93594 96676 93596
rect 96380 93542 96406 93594
rect 96406 93542 96436 93594
rect 96460 93542 96470 93594
rect 96470 93542 96516 93594
rect 96540 93542 96586 93594
rect 96586 93542 96596 93594
rect 96620 93542 96650 93594
rect 96650 93542 96676 93594
rect 96380 93540 96436 93542
rect 96460 93540 96516 93542
rect 96540 93540 96596 93542
rect 96620 93540 96676 93542
rect 96380 92506 96436 92508
rect 96460 92506 96516 92508
rect 96540 92506 96596 92508
rect 96620 92506 96676 92508
rect 96380 92454 96406 92506
rect 96406 92454 96436 92506
rect 96460 92454 96470 92506
rect 96470 92454 96516 92506
rect 96540 92454 96586 92506
rect 96586 92454 96596 92506
rect 96620 92454 96650 92506
rect 96650 92454 96676 92506
rect 96380 92452 96436 92454
rect 96460 92452 96516 92454
rect 96540 92452 96596 92454
rect 96620 92452 96676 92454
rect 96380 91418 96436 91420
rect 96460 91418 96516 91420
rect 96540 91418 96596 91420
rect 96620 91418 96676 91420
rect 96380 91366 96406 91418
rect 96406 91366 96436 91418
rect 96460 91366 96470 91418
rect 96470 91366 96516 91418
rect 96540 91366 96586 91418
rect 96586 91366 96596 91418
rect 96620 91366 96650 91418
rect 96650 91366 96676 91418
rect 96380 91364 96436 91366
rect 96460 91364 96516 91366
rect 96540 91364 96596 91366
rect 96620 91364 96676 91366
rect 96380 90330 96436 90332
rect 96460 90330 96516 90332
rect 96540 90330 96596 90332
rect 96620 90330 96676 90332
rect 96380 90278 96406 90330
rect 96406 90278 96436 90330
rect 96460 90278 96470 90330
rect 96470 90278 96516 90330
rect 96540 90278 96586 90330
rect 96586 90278 96596 90330
rect 96620 90278 96650 90330
rect 96650 90278 96676 90330
rect 96380 90276 96436 90278
rect 96460 90276 96516 90278
rect 96540 90276 96596 90278
rect 96620 90276 96676 90278
rect 96380 89242 96436 89244
rect 96460 89242 96516 89244
rect 96540 89242 96596 89244
rect 96620 89242 96676 89244
rect 96380 89190 96406 89242
rect 96406 89190 96436 89242
rect 96460 89190 96470 89242
rect 96470 89190 96516 89242
rect 96540 89190 96586 89242
rect 96586 89190 96596 89242
rect 96620 89190 96650 89242
rect 96650 89190 96676 89242
rect 96380 89188 96436 89190
rect 96460 89188 96516 89190
rect 96540 89188 96596 89190
rect 96620 89188 96676 89190
rect 96380 88154 96436 88156
rect 96460 88154 96516 88156
rect 96540 88154 96596 88156
rect 96620 88154 96676 88156
rect 96380 88102 96406 88154
rect 96406 88102 96436 88154
rect 96460 88102 96470 88154
rect 96470 88102 96516 88154
rect 96540 88102 96586 88154
rect 96586 88102 96596 88154
rect 96620 88102 96650 88154
rect 96650 88102 96676 88154
rect 96380 88100 96436 88102
rect 96460 88100 96516 88102
rect 96540 88100 96596 88102
rect 96620 88100 96676 88102
rect 96380 87066 96436 87068
rect 96460 87066 96516 87068
rect 96540 87066 96596 87068
rect 96620 87066 96676 87068
rect 96380 87014 96406 87066
rect 96406 87014 96436 87066
rect 96460 87014 96470 87066
rect 96470 87014 96516 87066
rect 96540 87014 96586 87066
rect 96586 87014 96596 87066
rect 96620 87014 96650 87066
rect 96650 87014 96676 87066
rect 96380 87012 96436 87014
rect 96460 87012 96516 87014
rect 96540 87012 96596 87014
rect 96620 87012 96676 87014
rect 96380 85978 96436 85980
rect 96460 85978 96516 85980
rect 96540 85978 96596 85980
rect 96620 85978 96676 85980
rect 96380 85926 96406 85978
rect 96406 85926 96436 85978
rect 96460 85926 96470 85978
rect 96470 85926 96516 85978
rect 96540 85926 96586 85978
rect 96586 85926 96596 85978
rect 96620 85926 96650 85978
rect 96650 85926 96676 85978
rect 96380 85924 96436 85926
rect 96460 85924 96516 85926
rect 96540 85924 96596 85926
rect 96620 85924 96676 85926
rect 96380 84890 96436 84892
rect 96460 84890 96516 84892
rect 96540 84890 96596 84892
rect 96620 84890 96676 84892
rect 96380 84838 96406 84890
rect 96406 84838 96436 84890
rect 96460 84838 96470 84890
rect 96470 84838 96516 84890
rect 96540 84838 96586 84890
rect 96586 84838 96596 84890
rect 96620 84838 96650 84890
rect 96650 84838 96676 84890
rect 96380 84836 96436 84838
rect 96460 84836 96516 84838
rect 96540 84836 96596 84838
rect 96620 84836 96676 84838
rect 96380 83802 96436 83804
rect 96460 83802 96516 83804
rect 96540 83802 96596 83804
rect 96620 83802 96676 83804
rect 96380 83750 96406 83802
rect 96406 83750 96436 83802
rect 96460 83750 96470 83802
rect 96470 83750 96516 83802
rect 96540 83750 96586 83802
rect 96586 83750 96596 83802
rect 96620 83750 96650 83802
rect 96650 83750 96676 83802
rect 96380 83748 96436 83750
rect 96460 83748 96516 83750
rect 96540 83748 96596 83750
rect 96620 83748 96676 83750
rect 96380 82714 96436 82716
rect 96460 82714 96516 82716
rect 96540 82714 96596 82716
rect 96620 82714 96676 82716
rect 96380 82662 96406 82714
rect 96406 82662 96436 82714
rect 96460 82662 96470 82714
rect 96470 82662 96516 82714
rect 96540 82662 96586 82714
rect 96586 82662 96596 82714
rect 96620 82662 96650 82714
rect 96650 82662 96676 82714
rect 96380 82660 96436 82662
rect 96460 82660 96516 82662
rect 96540 82660 96596 82662
rect 96620 82660 96676 82662
rect 96380 81626 96436 81628
rect 96460 81626 96516 81628
rect 96540 81626 96596 81628
rect 96620 81626 96676 81628
rect 96380 81574 96406 81626
rect 96406 81574 96436 81626
rect 96460 81574 96470 81626
rect 96470 81574 96516 81626
rect 96540 81574 96586 81626
rect 96586 81574 96596 81626
rect 96620 81574 96650 81626
rect 96650 81574 96676 81626
rect 96380 81572 96436 81574
rect 96460 81572 96516 81574
rect 96540 81572 96596 81574
rect 96620 81572 96676 81574
rect 96380 80538 96436 80540
rect 96460 80538 96516 80540
rect 96540 80538 96596 80540
rect 96620 80538 96676 80540
rect 96380 80486 96406 80538
rect 96406 80486 96436 80538
rect 96460 80486 96470 80538
rect 96470 80486 96516 80538
rect 96540 80486 96586 80538
rect 96586 80486 96596 80538
rect 96620 80486 96650 80538
rect 96650 80486 96676 80538
rect 96380 80484 96436 80486
rect 96460 80484 96516 80486
rect 96540 80484 96596 80486
rect 96620 80484 96676 80486
rect 96380 79450 96436 79452
rect 96460 79450 96516 79452
rect 96540 79450 96596 79452
rect 96620 79450 96676 79452
rect 96380 79398 96406 79450
rect 96406 79398 96436 79450
rect 96460 79398 96470 79450
rect 96470 79398 96516 79450
rect 96540 79398 96586 79450
rect 96586 79398 96596 79450
rect 96620 79398 96650 79450
rect 96650 79398 96676 79450
rect 96380 79396 96436 79398
rect 96460 79396 96516 79398
rect 96540 79396 96596 79398
rect 96620 79396 96676 79398
rect 96380 78362 96436 78364
rect 96460 78362 96516 78364
rect 96540 78362 96596 78364
rect 96620 78362 96676 78364
rect 96380 78310 96406 78362
rect 96406 78310 96436 78362
rect 96460 78310 96470 78362
rect 96470 78310 96516 78362
rect 96540 78310 96586 78362
rect 96586 78310 96596 78362
rect 96620 78310 96650 78362
rect 96650 78310 96676 78362
rect 96380 78308 96436 78310
rect 96460 78308 96516 78310
rect 96540 78308 96596 78310
rect 96620 78308 96676 78310
rect 96380 77274 96436 77276
rect 96460 77274 96516 77276
rect 96540 77274 96596 77276
rect 96620 77274 96676 77276
rect 96380 77222 96406 77274
rect 96406 77222 96436 77274
rect 96460 77222 96470 77274
rect 96470 77222 96516 77274
rect 96540 77222 96586 77274
rect 96586 77222 96596 77274
rect 96620 77222 96650 77274
rect 96650 77222 96676 77274
rect 96380 77220 96436 77222
rect 96460 77220 96516 77222
rect 96540 77220 96596 77222
rect 96620 77220 96676 77222
rect 96380 76186 96436 76188
rect 96460 76186 96516 76188
rect 96540 76186 96596 76188
rect 96620 76186 96676 76188
rect 96380 76134 96406 76186
rect 96406 76134 96436 76186
rect 96460 76134 96470 76186
rect 96470 76134 96516 76186
rect 96540 76134 96586 76186
rect 96586 76134 96596 76186
rect 96620 76134 96650 76186
rect 96650 76134 96676 76186
rect 96380 76132 96436 76134
rect 96460 76132 96516 76134
rect 96540 76132 96596 76134
rect 96620 76132 96676 76134
rect 96380 75098 96436 75100
rect 96460 75098 96516 75100
rect 96540 75098 96596 75100
rect 96620 75098 96676 75100
rect 96380 75046 96406 75098
rect 96406 75046 96436 75098
rect 96460 75046 96470 75098
rect 96470 75046 96516 75098
rect 96540 75046 96586 75098
rect 96586 75046 96596 75098
rect 96620 75046 96650 75098
rect 96650 75046 96676 75098
rect 96380 75044 96436 75046
rect 96460 75044 96516 75046
rect 96540 75044 96596 75046
rect 96620 75044 96676 75046
rect 96380 74010 96436 74012
rect 96460 74010 96516 74012
rect 96540 74010 96596 74012
rect 96620 74010 96676 74012
rect 96380 73958 96406 74010
rect 96406 73958 96436 74010
rect 96460 73958 96470 74010
rect 96470 73958 96516 74010
rect 96540 73958 96586 74010
rect 96586 73958 96596 74010
rect 96620 73958 96650 74010
rect 96650 73958 96676 74010
rect 96380 73956 96436 73958
rect 96460 73956 96516 73958
rect 96540 73956 96596 73958
rect 96620 73956 96676 73958
rect 96380 72922 96436 72924
rect 96460 72922 96516 72924
rect 96540 72922 96596 72924
rect 96620 72922 96676 72924
rect 96380 72870 96406 72922
rect 96406 72870 96436 72922
rect 96460 72870 96470 72922
rect 96470 72870 96516 72922
rect 96540 72870 96586 72922
rect 96586 72870 96596 72922
rect 96620 72870 96650 72922
rect 96650 72870 96676 72922
rect 96380 72868 96436 72870
rect 96460 72868 96516 72870
rect 96540 72868 96596 72870
rect 96620 72868 96676 72870
rect 96380 71834 96436 71836
rect 96460 71834 96516 71836
rect 96540 71834 96596 71836
rect 96620 71834 96676 71836
rect 96380 71782 96406 71834
rect 96406 71782 96436 71834
rect 96460 71782 96470 71834
rect 96470 71782 96516 71834
rect 96540 71782 96586 71834
rect 96586 71782 96596 71834
rect 96620 71782 96650 71834
rect 96650 71782 96676 71834
rect 96380 71780 96436 71782
rect 96460 71780 96516 71782
rect 96540 71780 96596 71782
rect 96620 71780 96676 71782
rect 96380 70746 96436 70748
rect 96460 70746 96516 70748
rect 96540 70746 96596 70748
rect 96620 70746 96676 70748
rect 96380 70694 96406 70746
rect 96406 70694 96436 70746
rect 96460 70694 96470 70746
rect 96470 70694 96516 70746
rect 96540 70694 96586 70746
rect 96586 70694 96596 70746
rect 96620 70694 96650 70746
rect 96650 70694 96676 70746
rect 96380 70692 96436 70694
rect 96460 70692 96516 70694
rect 96540 70692 96596 70694
rect 96620 70692 96676 70694
rect 96380 69658 96436 69660
rect 96460 69658 96516 69660
rect 96540 69658 96596 69660
rect 96620 69658 96676 69660
rect 96380 69606 96406 69658
rect 96406 69606 96436 69658
rect 96460 69606 96470 69658
rect 96470 69606 96516 69658
rect 96540 69606 96586 69658
rect 96586 69606 96596 69658
rect 96620 69606 96650 69658
rect 96650 69606 96676 69658
rect 96380 69604 96436 69606
rect 96460 69604 96516 69606
rect 96540 69604 96596 69606
rect 96620 69604 96676 69606
rect 96380 68570 96436 68572
rect 96460 68570 96516 68572
rect 96540 68570 96596 68572
rect 96620 68570 96676 68572
rect 96380 68518 96406 68570
rect 96406 68518 96436 68570
rect 96460 68518 96470 68570
rect 96470 68518 96516 68570
rect 96540 68518 96586 68570
rect 96586 68518 96596 68570
rect 96620 68518 96650 68570
rect 96650 68518 96676 68570
rect 96380 68516 96436 68518
rect 96460 68516 96516 68518
rect 96540 68516 96596 68518
rect 96620 68516 96676 68518
rect 96380 67482 96436 67484
rect 96460 67482 96516 67484
rect 96540 67482 96596 67484
rect 96620 67482 96676 67484
rect 96380 67430 96406 67482
rect 96406 67430 96436 67482
rect 96460 67430 96470 67482
rect 96470 67430 96516 67482
rect 96540 67430 96586 67482
rect 96586 67430 96596 67482
rect 96620 67430 96650 67482
rect 96650 67430 96676 67482
rect 96380 67428 96436 67430
rect 96460 67428 96516 67430
rect 96540 67428 96596 67430
rect 96620 67428 96676 67430
rect 96380 66394 96436 66396
rect 96460 66394 96516 66396
rect 96540 66394 96596 66396
rect 96620 66394 96676 66396
rect 96380 66342 96406 66394
rect 96406 66342 96436 66394
rect 96460 66342 96470 66394
rect 96470 66342 96516 66394
rect 96540 66342 96586 66394
rect 96586 66342 96596 66394
rect 96620 66342 96650 66394
rect 96650 66342 96676 66394
rect 96380 66340 96436 66342
rect 96460 66340 96516 66342
rect 96540 66340 96596 66342
rect 96620 66340 96676 66342
rect 96380 65306 96436 65308
rect 96460 65306 96516 65308
rect 96540 65306 96596 65308
rect 96620 65306 96676 65308
rect 96380 65254 96406 65306
rect 96406 65254 96436 65306
rect 96460 65254 96470 65306
rect 96470 65254 96516 65306
rect 96540 65254 96586 65306
rect 96586 65254 96596 65306
rect 96620 65254 96650 65306
rect 96650 65254 96676 65306
rect 96380 65252 96436 65254
rect 96460 65252 96516 65254
rect 96540 65252 96596 65254
rect 96620 65252 96676 65254
rect 96380 64218 96436 64220
rect 96460 64218 96516 64220
rect 96540 64218 96596 64220
rect 96620 64218 96676 64220
rect 96380 64166 96406 64218
rect 96406 64166 96436 64218
rect 96460 64166 96470 64218
rect 96470 64166 96516 64218
rect 96540 64166 96586 64218
rect 96586 64166 96596 64218
rect 96620 64166 96650 64218
rect 96650 64166 96676 64218
rect 96380 64164 96436 64166
rect 96460 64164 96516 64166
rect 96540 64164 96596 64166
rect 96620 64164 96676 64166
rect 96380 63130 96436 63132
rect 96460 63130 96516 63132
rect 96540 63130 96596 63132
rect 96620 63130 96676 63132
rect 96380 63078 96406 63130
rect 96406 63078 96436 63130
rect 96460 63078 96470 63130
rect 96470 63078 96516 63130
rect 96540 63078 96586 63130
rect 96586 63078 96596 63130
rect 96620 63078 96650 63130
rect 96650 63078 96676 63130
rect 96380 63076 96436 63078
rect 96460 63076 96516 63078
rect 96540 63076 96596 63078
rect 96620 63076 96676 63078
rect 96380 62042 96436 62044
rect 96460 62042 96516 62044
rect 96540 62042 96596 62044
rect 96620 62042 96676 62044
rect 96380 61990 96406 62042
rect 96406 61990 96436 62042
rect 96460 61990 96470 62042
rect 96470 61990 96516 62042
rect 96540 61990 96586 62042
rect 96586 61990 96596 62042
rect 96620 61990 96650 62042
rect 96650 61990 96676 62042
rect 96380 61988 96436 61990
rect 96460 61988 96516 61990
rect 96540 61988 96596 61990
rect 96620 61988 96676 61990
rect 96380 60954 96436 60956
rect 96460 60954 96516 60956
rect 96540 60954 96596 60956
rect 96620 60954 96676 60956
rect 96380 60902 96406 60954
rect 96406 60902 96436 60954
rect 96460 60902 96470 60954
rect 96470 60902 96516 60954
rect 96540 60902 96586 60954
rect 96586 60902 96596 60954
rect 96620 60902 96650 60954
rect 96650 60902 96676 60954
rect 96380 60900 96436 60902
rect 96460 60900 96516 60902
rect 96540 60900 96596 60902
rect 96620 60900 96676 60902
rect 96380 59866 96436 59868
rect 96460 59866 96516 59868
rect 96540 59866 96596 59868
rect 96620 59866 96676 59868
rect 96380 59814 96406 59866
rect 96406 59814 96436 59866
rect 96460 59814 96470 59866
rect 96470 59814 96516 59866
rect 96540 59814 96586 59866
rect 96586 59814 96596 59866
rect 96620 59814 96650 59866
rect 96650 59814 96676 59866
rect 96380 59812 96436 59814
rect 96460 59812 96516 59814
rect 96540 59812 96596 59814
rect 96620 59812 96676 59814
rect 96380 58778 96436 58780
rect 96460 58778 96516 58780
rect 96540 58778 96596 58780
rect 96620 58778 96676 58780
rect 96380 58726 96406 58778
rect 96406 58726 96436 58778
rect 96460 58726 96470 58778
rect 96470 58726 96516 58778
rect 96540 58726 96586 58778
rect 96586 58726 96596 58778
rect 96620 58726 96650 58778
rect 96650 58726 96676 58778
rect 96380 58724 96436 58726
rect 96460 58724 96516 58726
rect 96540 58724 96596 58726
rect 96620 58724 96676 58726
rect 96380 57690 96436 57692
rect 96460 57690 96516 57692
rect 96540 57690 96596 57692
rect 96620 57690 96676 57692
rect 96380 57638 96406 57690
rect 96406 57638 96436 57690
rect 96460 57638 96470 57690
rect 96470 57638 96516 57690
rect 96540 57638 96586 57690
rect 96586 57638 96596 57690
rect 96620 57638 96650 57690
rect 96650 57638 96676 57690
rect 96380 57636 96436 57638
rect 96460 57636 96516 57638
rect 96540 57636 96596 57638
rect 96620 57636 96676 57638
rect 96380 56602 96436 56604
rect 96460 56602 96516 56604
rect 96540 56602 96596 56604
rect 96620 56602 96676 56604
rect 96380 56550 96406 56602
rect 96406 56550 96436 56602
rect 96460 56550 96470 56602
rect 96470 56550 96516 56602
rect 96540 56550 96586 56602
rect 96586 56550 96596 56602
rect 96620 56550 96650 56602
rect 96650 56550 96676 56602
rect 96380 56548 96436 56550
rect 96460 56548 96516 56550
rect 96540 56548 96596 56550
rect 96620 56548 96676 56550
rect 96380 55514 96436 55516
rect 96460 55514 96516 55516
rect 96540 55514 96596 55516
rect 96620 55514 96676 55516
rect 96380 55462 96406 55514
rect 96406 55462 96436 55514
rect 96460 55462 96470 55514
rect 96470 55462 96516 55514
rect 96540 55462 96586 55514
rect 96586 55462 96596 55514
rect 96620 55462 96650 55514
rect 96650 55462 96676 55514
rect 96380 55460 96436 55462
rect 96460 55460 96516 55462
rect 96540 55460 96596 55462
rect 96620 55460 96676 55462
rect 96380 54426 96436 54428
rect 96460 54426 96516 54428
rect 96540 54426 96596 54428
rect 96620 54426 96676 54428
rect 96380 54374 96406 54426
rect 96406 54374 96436 54426
rect 96460 54374 96470 54426
rect 96470 54374 96516 54426
rect 96540 54374 96586 54426
rect 96586 54374 96596 54426
rect 96620 54374 96650 54426
rect 96650 54374 96676 54426
rect 96380 54372 96436 54374
rect 96460 54372 96516 54374
rect 96540 54372 96596 54374
rect 96620 54372 96676 54374
rect 96380 53338 96436 53340
rect 96460 53338 96516 53340
rect 96540 53338 96596 53340
rect 96620 53338 96676 53340
rect 96380 53286 96406 53338
rect 96406 53286 96436 53338
rect 96460 53286 96470 53338
rect 96470 53286 96516 53338
rect 96540 53286 96586 53338
rect 96586 53286 96596 53338
rect 96620 53286 96650 53338
rect 96650 53286 96676 53338
rect 96380 53284 96436 53286
rect 96460 53284 96516 53286
rect 96540 53284 96596 53286
rect 96620 53284 96676 53286
rect 96380 52250 96436 52252
rect 96460 52250 96516 52252
rect 96540 52250 96596 52252
rect 96620 52250 96676 52252
rect 96380 52198 96406 52250
rect 96406 52198 96436 52250
rect 96460 52198 96470 52250
rect 96470 52198 96516 52250
rect 96540 52198 96586 52250
rect 96586 52198 96596 52250
rect 96620 52198 96650 52250
rect 96650 52198 96676 52250
rect 96380 52196 96436 52198
rect 96460 52196 96516 52198
rect 96540 52196 96596 52198
rect 96620 52196 96676 52198
rect 96380 51162 96436 51164
rect 96460 51162 96516 51164
rect 96540 51162 96596 51164
rect 96620 51162 96676 51164
rect 96380 51110 96406 51162
rect 96406 51110 96436 51162
rect 96460 51110 96470 51162
rect 96470 51110 96516 51162
rect 96540 51110 96586 51162
rect 96586 51110 96596 51162
rect 96620 51110 96650 51162
rect 96650 51110 96676 51162
rect 96380 51108 96436 51110
rect 96460 51108 96516 51110
rect 96540 51108 96596 51110
rect 96620 51108 96676 51110
rect 96380 50074 96436 50076
rect 96460 50074 96516 50076
rect 96540 50074 96596 50076
rect 96620 50074 96676 50076
rect 96380 50022 96406 50074
rect 96406 50022 96436 50074
rect 96460 50022 96470 50074
rect 96470 50022 96516 50074
rect 96540 50022 96586 50074
rect 96586 50022 96596 50074
rect 96620 50022 96650 50074
rect 96650 50022 96676 50074
rect 96380 50020 96436 50022
rect 96460 50020 96516 50022
rect 96540 50020 96596 50022
rect 96620 50020 96676 50022
rect 96380 48986 96436 48988
rect 96460 48986 96516 48988
rect 96540 48986 96596 48988
rect 96620 48986 96676 48988
rect 96380 48934 96406 48986
rect 96406 48934 96436 48986
rect 96460 48934 96470 48986
rect 96470 48934 96516 48986
rect 96540 48934 96586 48986
rect 96586 48934 96596 48986
rect 96620 48934 96650 48986
rect 96650 48934 96676 48986
rect 96380 48932 96436 48934
rect 96460 48932 96516 48934
rect 96540 48932 96596 48934
rect 96620 48932 96676 48934
rect 96380 47898 96436 47900
rect 96460 47898 96516 47900
rect 96540 47898 96596 47900
rect 96620 47898 96676 47900
rect 96380 47846 96406 47898
rect 96406 47846 96436 47898
rect 96460 47846 96470 47898
rect 96470 47846 96516 47898
rect 96540 47846 96586 47898
rect 96586 47846 96596 47898
rect 96620 47846 96650 47898
rect 96650 47846 96676 47898
rect 96380 47844 96436 47846
rect 96460 47844 96516 47846
rect 96540 47844 96596 47846
rect 96620 47844 96676 47846
rect 96380 46810 96436 46812
rect 96460 46810 96516 46812
rect 96540 46810 96596 46812
rect 96620 46810 96676 46812
rect 96380 46758 96406 46810
rect 96406 46758 96436 46810
rect 96460 46758 96470 46810
rect 96470 46758 96516 46810
rect 96540 46758 96586 46810
rect 96586 46758 96596 46810
rect 96620 46758 96650 46810
rect 96650 46758 96676 46810
rect 96380 46756 96436 46758
rect 96460 46756 96516 46758
rect 96540 46756 96596 46758
rect 96620 46756 96676 46758
rect 96380 45722 96436 45724
rect 96460 45722 96516 45724
rect 96540 45722 96596 45724
rect 96620 45722 96676 45724
rect 96380 45670 96406 45722
rect 96406 45670 96436 45722
rect 96460 45670 96470 45722
rect 96470 45670 96516 45722
rect 96540 45670 96586 45722
rect 96586 45670 96596 45722
rect 96620 45670 96650 45722
rect 96650 45670 96676 45722
rect 96380 45668 96436 45670
rect 96460 45668 96516 45670
rect 96540 45668 96596 45670
rect 96620 45668 96676 45670
rect 96380 44634 96436 44636
rect 96460 44634 96516 44636
rect 96540 44634 96596 44636
rect 96620 44634 96676 44636
rect 96380 44582 96406 44634
rect 96406 44582 96436 44634
rect 96460 44582 96470 44634
rect 96470 44582 96516 44634
rect 96540 44582 96586 44634
rect 96586 44582 96596 44634
rect 96620 44582 96650 44634
rect 96650 44582 96676 44634
rect 96380 44580 96436 44582
rect 96460 44580 96516 44582
rect 96540 44580 96596 44582
rect 96620 44580 96676 44582
rect 96380 43546 96436 43548
rect 96460 43546 96516 43548
rect 96540 43546 96596 43548
rect 96620 43546 96676 43548
rect 96380 43494 96406 43546
rect 96406 43494 96436 43546
rect 96460 43494 96470 43546
rect 96470 43494 96516 43546
rect 96540 43494 96586 43546
rect 96586 43494 96596 43546
rect 96620 43494 96650 43546
rect 96650 43494 96676 43546
rect 96380 43492 96436 43494
rect 96460 43492 96516 43494
rect 96540 43492 96596 43494
rect 96620 43492 96676 43494
rect 96380 42458 96436 42460
rect 96460 42458 96516 42460
rect 96540 42458 96596 42460
rect 96620 42458 96676 42460
rect 96380 42406 96406 42458
rect 96406 42406 96436 42458
rect 96460 42406 96470 42458
rect 96470 42406 96516 42458
rect 96540 42406 96586 42458
rect 96586 42406 96596 42458
rect 96620 42406 96650 42458
rect 96650 42406 96676 42458
rect 96380 42404 96436 42406
rect 96460 42404 96516 42406
rect 96540 42404 96596 42406
rect 96620 42404 96676 42406
rect 96380 41370 96436 41372
rect 96460 41370 96516 41372
rect 96540 41370 96596 41372
rect 96620 41370 96676 41372
rect 96380 41318 96406 41370
rect 96406 41318 96436 41370
rect 96460 41318 96470 41370
rect 96470 41318 96516 41370
rect 96540 41318 96586 41370
rect 96586 41318 96596 41370
rect 96620 41318 96650 41370
rect 96650 41318 96676 41370
rect 96380 41316 96436 41318
rect 96460 41316 96516 41318
rect 96540 41316 96596 41318
rect 96620 41316 96676 41318
rect 96380 40282 96436 40284
rect 96460 40282 96516 40284
rect 96540 40282 96596 40284
rect 96620 40282 96676 40284
rect 96380 40230 96406 40282
rect 96406 40230 96436 40282
rect 96460 40230 96470 40282
rect 96470 40230 96516 40282
rect 96540 40230 96586 40282
rect 96586 40230 96596 40282
rect 96620 40230 96650 40282
rect 96650 40230 96676 40282
rect 96380 40228 96436 40230
rect 96460 40228 96516 40230
rect 96540 40228 96596 40230
rect 96620 40228 96676 40230
rect 96380 39194 96436 39196
rect 96460 39194 96516 39196
rect 96540 39194 96596 39196
rect 96620 39194 96676 39196
rect 96380 39142 96406 39194
rect 96406 39142 96436 39194
rect 96460 39142 96470 39194
rect 96470 39142 96516 39194
rect 96540 39142 96586 39194
rect 96586 39142 96596 39194
rect 96620 39142 96650 39194
rect 96650 39142 96676 39194
rect 96380 39140 96436 39142
rect 96460 39140 96516 39142
rect 96540 39140 96596 39142
rect 96620 39140 96676 39142
rect 96380 38106 96436 38108
rect 96460 38106 96516 38108
rect 96540 38106 96596 38108
rect 96620 38106 96676 38108
rect 96380 38054 96406 38106
rect 96406 38054 96436 38106
rect 96460 38054 96470 38106
rect 96470 38054 96516 38106
rect 96540 38054 96586 38106
rect 96586 38054 96596 38106
rect 96620 38054 96650 38106
rect 96650 38054 96676 38106
rect 96380 38052 96436 38054
rect 96460 38052 96516 38054
rect 96540 38052 96596 38054
rect 96620 38052 96676 38054
rect 96380 37018 96436 37020
rect 96460 37018 96516 37020
rect 96540 37018 96596 37020
rect 96620 37018 96676 37020
rect 96380 36966 96406 37018
rect 96406 36966 96436 37018
rect 96460 36966 96470 37018
rect 96470 36966 96516 37018
rect 96540 36966 96586 37018
rect 96586 36966 96596 37018
rect 96620 36966 96650 37018
rect 96650 36966 96676 37018
rect 96380 36964 96436 36966
rect 96460 36964 96516 36966
rect 96540 36964 96596 36966
rect 96620 36964 96676 36966
rect 96380 35930 96436 35932
rect 96460 35930 96516 35932
rect 96540 35930 96596 35932
rect 96620 35930 96676 35932
rect 96380 35878 96406 35930
rect 96406 35878 96436 35930
rect 96460 35878 96470 35930
rect 96470 35878 96516 35930
rect 96540 35878 96586 35930
rect 96586 35878 96596 35930
rect 96620 35878 96650 35930
rect 96650 35878 96676 35930
rect 96380 35876 96436 35878
rect 96460 35876 96516 35878
rect 96540 35876 96596 35878
rect 96620 35876 96676 35878
rect 96380 34842 96436 34844
rect 96460 34842 96516 34844
rect 96540 34842 96596 34844
rect 96620 34842 96676 34844
rect 96380 34790 96406 34842
rect 96406 34790 96436 34842
rect 96460 34790 96470 34842
rect 96470 34790 96516 34842
rect 96540 34790 96586 34842
rect 96586 34790 96596 34842
rect 96620 34790 96650 34842
rect 96650 34790 96676 34842
rect 96380 34788 96436 34790
rect 96460 34788 96516 34790
rect 96540 34788 96596 34790
rect 96620 34788 96676 34790
rect 96380 33754 96436 33756
rect 96460 33754 96516 33756
rect 96540 33754 96596 33756
rect 96620 33754 96676 33756
rect 96380 33702 96406 33754
rect 96406 33702 96436 33754
rect 96460 33702 96470 33754
rect 96470 33702 96516 33754
rect 96540 33702 96586 33754
rect 96586 33702 96596 33754
rect 96620 33702 96650 33754
rect 96650 33702 96676 33754
rect 96380 33700 96436 33702
rect 96460 33700 96516 33702
rect 96540 33700 96596 33702
rect 96620 33700 96676 33702
rect 96380 32666 96436 32668
rect 96460 32666 96516 32668
rect 96540 32666 96596 32668
rect 96620 32666 96676 32668
rect 96380 32614 96406 32666
rect 96406 32614 96436 32666
rect 96460 32614 96470 32666
rect 96470 32614 96516 32666
rect 96540 32614 96586 32666
rect 96586 32614 96596 32666
rect 96620 32614 96650 32666
rect 96650 32614 96676 32666
rect 96380 32612 96436 32614
rect 96460 32612 96516 32614
rect 96540 32612 96596 32614
rect 96620 32612 96676 32614
rect 96380 31578 96436 31580
rect 96460 31578 96516 31580
rect 96540 31578 96596 31580
rect 96620 31578 96676 31580
rect 96380 31526 96406 31578
rect 96406 31526 96436 31578
rect 96460 31526 96470 31578
rect 96470 31526 96516 31578
rect 96540 31526 96586 31578
rect 96586 31526 96596 31578
rect 96620 31526 96650 31578
rect 96650 31526 96676 31578
rect 96380 31524 96436 31526
rect 96460 31524 96516 31526
rect 96540 31524 96596 31526
rect 96620 31524 96676 31526
rect 96380 30490 96436 30492
rect 96460 30490 96516 30492
rect 96540 30490 96596 30492
rect 96620 30490 96676 30492
rect 96380 30438 96406 30490
rect 96406 30438 96436 30490
rect 96460 30438 96470 30490
rect 96470 30438 96516 30490
rect 96540 30438 96586 30490
rect 96586 30438 96596 30490
rect 96620 30438 96650 30490
rect 96650 30438 96676 30490
rect 96380 30436 96436 30438
rect 96460 30436 96516 30438
rect 96540 30436 96596 30438
rect 96620 30436 96676 30438
rect 96380 29402 96436 29404
rect 96460 29402 96516 29404
rect 96540 29402 96596 29404
rect 96620 29402 96676 29404
rect 96380 29350 96406 29402
rect 96406 29350 96436 29402
rect 96460 29350 96470 29402
rect 96470 29350 96516 29402
rect 96540 29350 96586 29402
rect 96586 29350 96596 29402
rect 96620 29350 96650 29402
rect 96650 29350 96676 29402
rect 96380 29348 96436 29350
rect 96460 29348 96516 29350
rect 96540 29348 96596 29350
rect 96620 29348 96676 29350
rect 96380 28314 96436 28316
rect 96460 28314 96516 28316
rect 96540 28314 96596 28316
rect 96620 28314 96676 28316
rect 96380 28262 96406 28314
rect 96406 28262 96436 28314
rect 96460 28262 96470 28314
rect 96470 28262 96516 28314
rect 96540 28262 96586 28314
rect 96586 28262 96596 28314
rect 96620 28262 96650 28314
rect 96650 28262 96676 28314
rect 96380 28260 96436 28262
rect 96460 28260 96516 28262
rect 96540 28260 96596 28262
rect 96620 28260 96676 28262
rect 96380 27226 96436 27228
rect 96460 27226 96516 27228
rect 96540 27226 96596 27228
rect 96620 27226 96676 27228
rect 96380 27174 96406 27226
rect 96406 27174 96436 27226
rect 96460 27174 96470 27226
rect 96470 27174 96516 27226
rect 96540 27174 96586 27226
rect 96586 27174 96596 27226
rect 96620 27174 96650 27226
rect 96650 27174 96676 27226
rect 96380 27172 96436 27174
rect 96460 27172 96516 27174
rect 96540 27172 96596 27174
rect 96620 27172 96676 27174
rect 96380 26138 96436 26140
rect 96460 26138 96516 26140
rect 96540 26138 96596 26140
rect 96620 26138 96676 26140
rect 96380 26086 96406 26138
rect 96406 26086 96436 26138
rect 96460 26086 96470 26138
rect 96470 26086 96516 26138
rect 96540 26086 96586 26138
rect 96586 26086 96596 26138
rect 96620 26086 96650 26138
rect 96650 26086 96676 26138
rect 96380 26084 96436 26086
rect 96460 26084 96516 26086
rect 96540 26084 96596 26086
rect 96620 26084 96676 26086
rect 96380 25050 96436 25052
rect 96460 25050 96516 25052
rect 96540 25050 96596 25052
rect 96620 25050 96676 25052
rect 96380 24998 96406 25050
rect 96406 24998 96436 25050
rect 96460 24998 96470 25050
rect 96470 24998 96516 25050
rect 96540 24998 96586 25050
rect 96586 24998 96596 25050
rect 96620 24998 96650 25050
rect 96650 24998 96676 25050
rect 96380 24996 96436 24998
rect 96460 24996 96516 24998
rect 96540 24996 96596 24998
rect 96620 24996 96676 24998
rect 96380 23962 96436 23964
rect 96460 23962 96516 23964
rect 96540 23962 96596 23964
rect 96620 23962 96676 23964
rect 96380 23910 96406 23962
rect 96406 23910 96436 23962
rect 96460 23910 96470 23962
rect 96470 23910 96516 23962
rect 96540 23910 96586 23962
rect 96586 23910 96596 23962
rect 96620 23910 96650 23962
rect 96650 23910 96676 23962
rect 96380 23908 96436 23910
rect 96460 23908 96516 23910
rect 96540 23908 96596 23910
rect 96620 23908 96676 23910
rect 96380 22874 96436 22876
rect 96460 22874 96516 22876
rect 96540 22874 96596 22876
rect 96620 22874 96676 22876
rect 96380 22822 96406 22874
rect 96406 22822 96436 22874
rect 96460 22822 96470 22874
rect 96470 22822 96516 22874
rect 96540 22822 96586 22874
rect 96586 22822 96596 22874
rect 96620 22822 96650 22874
rect 96650 22822 96676 22874
rect 96380 22820 96436 22822
rect 96460 22820 96516 22822
rect 96540 22820 96596 22822
rect 96620 22820 96676 22822
rect 96380 21786 96436 21788
rect 96460 21786 96516 21788
rect 96540 21786 96596 21788
rect 96620 21786 96676 21788
rect 96380 21734 96406 21786
rect 96406 21734 96436 21786
rect 96460 21734 96470 21786
rect 96470 21734 96516 21786
rect 96540 21734 96586 21786
rect 96586 21734 96596 21786
rect 96620 21734 96650 21786
rect 96650 21734 96676 21786
rect 96380 21732 96436 21734
rect 96460 21732 96516 21734
rect 96540 21732 96596 21734
rect 96620 21732 96676 21734
rect 96380 20698 96436 20700
rect 96460 20698 96516 20700
rect 96540 20698 96596 20700
rect 96620 20698 96676 20700
rect 96380 20646 96406 20698
rect 96406 20646 96436 20698
rect 96460 20646 96470 20698
rect 96470 20646 96516 20698
rect 96540 20646 96586 20698
rect 96586 20646 96596 20698
rect 96620 20646 96650 20698
rect 96650 20646 96676 20698
rect 96380 20644 96436 20646
rect 96460 20644 96516 20646
rect 96540 20644 96596 20646
rect 96620 20644 96676 20646
rect 96380 19610 96436 19612
rect 96460 19610 96516 19612
rect 96540 19610 96596 19612
rect 96620 19610 96676 19612
rect 96380 19558 96406 19610
rect 96406 19558 96436 19610
rect 96460 19558 96470 19610
rect 96470 19558 96516 19610
rect 96540 19558 96586 19610
rect 96586 19558 96596 19610
rect 96620 19558 96650 19610
rect 96650 19558 96676 19610
rect 96380 19556 96436 19558
rect 96460 19556 96516 19558
rect 96540 19556 96596 19558
rect 96620 19556 96676 19558
rect 96380 18522 96436 18524
rect 96460 18522 96516 18524
rect 96540 18522 96596 18524
rect 96620 18522 96676 18524
rect 96380 18470 96406 18522
rect 96406 18470 96436 18522
rect 96460 18470 96470 18522
rect 96470 18470 96516 18522
rect 96540 18470 96586 18522
rect 96586 18470 96596 18522
rect 96620 18470 96650 18522
rect 96650 18470 96676 18522
rect 96380 18468 96436 18470
rect 96460 18468 96516 18470
rect 96540 18468 96596 18470
rect 96620 18468 96676 18470
rect 96380 17434 96436 17436
rect 96460 17434 96516 17436
rect 96540 17434 96596 17436
rect 96620 17434 96676 17436
rect 96380 17382 96406 17434
rect 96406 17382 96436 17434
rect 96460 17382 96470 17434
rect 96470 17382 96516 17434
rect 96540 17382 96586 17434
rect 96586 17382 96596 17434
rect 96620 17382 96650 17434
rect 96650 17382 96676 17434
rect 96380 17380 96436 17382
rect 96460 17380 96516 17382
rect 96540 17380 96596 17382
rect 96620 17380 96676 17382
rect 96380 16346 96436 16348
rect 96460 16346 96516 16348
rect 96540 16346 96596 16348
rect 96620 16346 96676 16348
rect 96380 16294 96406 16346
rect 96406 16294 96436 16346
rect 96460 16294 96470 16346
rect 96470 16294 96516 16346
rect 96540 16294 96586 16346
rect 96586 16294 96596 16346
rect 96620 16294 96650 16346
rect 96650 16294 96676 16346
rect 96380 16292 96436 16294
rect 96460 16292 96516 16294
rect 96540 16292 96596 16294
rect 96620 16292 96676 16294
rect 96380 15258 96436 15260
rect 96460 15258 96516 15260
rect 96540 15258 96596 15260
rect 96620 15258 96676 15260
rect 96380 15206 96406 15258
rect 96406 15206 96436 15258
rect 96460 15206 96470 15258
rect 96470 15206 96516 15258
rect 96540 15206 96586 15258
rect 96586 15206 96596 15258
rect 96620 15206 96650 15258
rect 96650 15206 96676 15258
rect 96380 15204 96436 15206
rect 96460 15204 96516 15206
rect 96540 15204 96596 15206
rect 96620 15204 96676 15206
rect 96380 14170 96436 14172
rect 96460 14170 96516 14172
rect 96540 14170 96596 14172
rect 96620 14170 96676 14172
rect 96380 14118 96406 14170
rect 96406 14118 96436 14170
rect 96460 14118 96470 14170
rect 96470 14118 96516 14170
rect 96540 14118 96586 14170
rect 96586 14118 96596 14170
rect 96620 14118 96650 14170
rect 96650 14118 96676 14170
rect 96380 14116 96436 14118
rect 96460 14116 96516 14118
rect 96540 14116 96596 14118
rect 96620 14116 96676 14118
rect 96380 13082 96436 13084
rect 96460 13082 96516 13084
rect 96540 13082 96596 13084
rect 96620 13082 96676 13084
rect 96380 13030 96406 13082
rect 96406 13030 96436 13082
rect 96460 13030 96470 13082
rect 96470 13030 96516 13082
rect 96540 13030 96586 13082
rect 96586 13030 96596 13082
rect 96620 13030 96650 13082
rect 96650 13030 96676 13082
rect 96380 13028 96436 13030
rect 96460 13028 96516 13030
rect 96540 13028 96596 13030
rect 96620 13028 96676 13030
rect 96380 11994 96436 11996
rect 96460 11994 96516 11996
rect 96540 11994 96596 11996
rect 96620 11994 96676 11996
rect 96380 11942 96406 11994
rect 96406 11942 96436 11994
rect 96460 11942 96470 11994
rect 96470 11942 96516 11994
rect 96540 11942 96586 11994
rect 96586 11942 96596 11994
rect 96620 11942 96650 11994
rect 96650 11942 96676 11994
rect 96380 11940 96436 11942
rect 96460 11940 96516 11942
rect 96540 11940 96596 11942
rect 96620 11940 96676 11942
rect 96380 10906 96436 10908
rect 96460 10906 96516 10908
rect 96540 10906 96596 10908
rect 96620 10906 96676 10908
rect 96380 10854 96406 10906
rect 96406 10854 96436 10906
rect 96460 10854 96470 10906
rect 96470 10854 96516 10906
rect 96540 10854 96586 10906
rect 96586 10854 96596 10906
rect 96620 10854 96650 10906
rect 96650 10854 96676 10906
rect 96380 10852 96436 10854
rect 96460 10852 96516 10854
rect 96540 10852 96596 10854
rect 96620 10852 96676 10854
rect 96380 9818 96436 9820
rect 96460 9818 96516 9820
rect 96540 9818 96596 9820
rect 96620 9818 96676 9820
rect 96380 9766 96406 9818
rect 96406 9766 96436 9818
rect 96460 9766 96470 9818
rect 96470 9766 96516 9818
rect 96540 9766 96586 9818
rect 96586 9766 96596 9818
rect 96620 9766 96650 9818
rect 96650 9766 96676 9818
rect 96380 9764 96436 9766
rect 96460 9764 96516 9766
rect 96540 9764 96596 9766
rect 96620 9764 96676 9766
rect 96380 8730 96436 8732
rect 96460 8730 96516 8732
rect 96540 8730 96596 8732
rect 96620 8730 96676 8732
rect 96380 8678 96406 8730
rect 96406 8678 96436 8730
rect 96460 8678 96470 8730
rect 96470 8678 96516 8730
rect 96540 8678 96586 8730
rect 96586 8678 96596 8730
rect 96620 8678 96650 8730
rect 96650 8678 96676 8730
rect 96380 8676 96436 8678
rect 96460 8676 96516 8678
rect 96540 8676 96596 8678
rect 96620 8676 96676 8678
rect 96380 7642 96436 7644
rect 96460 7642 96516 7644
rect 96540 7642 96596 7644
rect 96620 7642 96676 7644
rect 96380 7590 96406 7642
rect 96406 7590 96436 7642
rect 96460 7590 96470 7642
rect 96470 7590 96516 7642
rect 96540 7590 96586 7642
rect 96586 7590 96596 7642
rect 96620 7590 96650 7642
rect 96650 7590 96676 7642
rect 96380 7588 96436 7590
rect 96460 7588 96516 7590
rect 96540 7588 96596 7590
rect 96620 7588 96676 7590
rect 96380 6554 96436 6556
rect 96460 6554 96516 6556
rect 96540 6554 96596 6556
rect 96620 6554 96676 6556
rect 96380 6502 96406 6554
rect 96406 6502 96436 6554
rect 96460 6502 96470 6554
rect 96470 6502 96516 6554
rect 96540 6502 96586 6554
rect 96586 6502 96596 6554
rect 96620 6502 96650 6554
rect 96650 6502 96676 6554
rect 96380 6500 96436 6502
rect 96460 6500 96516 6502
rect 96540 6500 96596 6502
rect 96620 6500 96676 6502
rect 96380 5466 96436 5468
rect 96460 5466 96516 5468
rect 96540 5466 96596 5468
rect 96620 5466 96676 5468
rect 96380 5414 96406 5466
rect 96406 5414 96436 5466
rect 96460 5414 96470 5466
rect 96470 5414 96516 5466
rect 96540 5414 96586 5466
rect 96586 5414 96596 5466
rect 96620 5414 96650 5466
rect 96650 5414 96676 5466
rect 96380 5412 96436 5414
rect 96460 5412 96516 5414
rect 96540 5412 96596 5414
rect 96620 5412 96676 5414
rect 96380 4378 96436 4380
rect 96460 4378 96516 4380
rect 96540 4378 96596 4380
rect 96620 4378 96676 4380
rect 96380 4326 96406 4378
rect 96406 4326 96436 4378
rect 96460 4326 96470 4378
rect 96470 4326 96516 4378
rect 96540 4326 96586 4378
rect 96586 4326 96596 4378
rect 96620 4326 96650 4378
rect 96650 4326 96676 4378
rect 96380 4324 96436 4326
rect 96460 4324 96516 4326
rect 96540 4324 96596 4326
rect 96620 4324 96676 4326
rect 96380 3290 96436 3292
rect 96460 3290 96516 3292
rect 96540 3290 96596 3292
rect 96620 3290 96676 3292
rect 96380 3238 96406 3290
rect 96406 3238 96436 3290
rect 96460 3238 96470 3290
rect 96470 3238 96516 3290
rect 96540 3238 96586 3290
rect 96586 3238 96596 3290
rect 96620 3238 96650 3290
rect 96650 3238 96676 3290
rect 96380 3236 96436 3238
rect 96460 3236 96516 3238
rect 96540 3236 96596 3238
rect 96620 3236 96676 3238
rect 96380 2202 96436 2204
rect 96460 2202 96516 2204
rect 96540 2202 96596 2204
rect 96620 2202 96676 2204
rect 96380 2150 96406 2202
rect 96406 2150 96436 2202
rect 96460 2150 96470 2202
rect 96470 2150 96516 2202
rect 96540 2150 96586 2202
rect 96586 2150 96596 2202
rect 96620 2150 96650 2202
rect 96650 2150 96676 2202
rect 96380 2148 96436 2150
rect 96460 2148 96516 2150
rect 96540 2148 96596 2150
rect 96620 2148 96676 2150
<< metal3 >>
rect 19568 97408 19888 97409
rect 19568 97344 19576 97408
rect 19640 97344 19656 97408
rect 19720 97344 19736 97408
rect 19800 97344 19816 97408
rect 19880 97344 19888 97408
rect 19568 97343 19888 97344
rect 50288 97408 50608 97409
rect 50288 97344 50296 97408
rect 50360 97344 50376 97408
rect 50440 97344 50456 97408
rect 50520 97344 50536 97408
rect 50600 97344 50608 97408
rect 50288 97343 50608 97344
rect 81008 97408 81328 97409
rect 81008 97344 81016 97408
rect 81080 97344 81096 97408
rect 81160 97344 81176 97408
rect 81240 97344 81256 97408
rect 81320 97344 81328 97408
rect 81008 97343 81328 97344
rect 4208 96864 4528 96865
rect 4208 96800 4216 96864
rect 4280 96800 4296 96864
rect 4360 96800 4376 96864
rect 4440 96800 4456 96864
rect 4520 96800 4528 96864
rect 4208 96799 4528 96800
rect 34928 96864 35248 96865
rect 34928 96800 34936 96864
rect 35000 96800 35016 96864
rect 35080 96800 35096 96864
rect 35160 96800 35176 96864
rect 35240 96800 35248 96864
rect 34928 96799 35248 96800
rect 65648 96864 65968 96865
rect 65648 96800 65656 96864
rect 65720 96800 65736 96864
rect 65800 96800 65816 96864
rect 65880 96800 65896 96864
rect 65960 96800 65968 96864
rect 65648 96799 65968 96800
rect 96368 96864 96688 96865
rect 96368 96800 96376 96864
rect 96440 96800 96456 96864
rect 96520 96800 96536 96864
rect 96600 96800 96616 96864
rect 96680 96800 96688 96864
rect 96368 96799 96688 96800
rect 19568 96320 19888 96321
rect 19568 96256 19576 96320
rect 19640 96256 19656 96320
rect 19720 96256 19736 96320
rect 19800 96256 19816 96320
rect 19880 96256 19888 96320
rect 19568 96255 19888 96256
rect 50288 96320 50608 96321
rect 50288 96256 50296 96320
rect 50360 96256 50376 96320
rect 50440 96256 50456 96320
rect 50520 96256 50536 96320
rect 50600 96256 50608 96320
rect 50288 96255 50608 96256
rect 81008 96320 81328 96321
rect 81008 96256 81016 96320
rect 81080 96256 81096 96320
rect 81160 96256 81176 96320
rect 81240 96256 81256 96320
rect 81320 96256 81328 96320
rect 81008 96255 81328 96256
rect 4208 95776 4528 95777
rect 4208 95712 4216 95776
rect 4280 95712 4296 95776
rect 4360 95712 4376 95776
rect 4440 95712 4456 95776
rect 4520 95712 4528 95776
rect 4208 95711 4528 95712
rect 34928 95776 35248 95777
rect 34928 95712 34936 95776
rect 35000 95712 35016 95776
rect 35080 95712 35096 95776
rect 35160 95712 35176 95776
rect 35240 95712 35248 95776
rect 34928 95711 35248 95712
rect 65648 95776 65968 95777
rect 65648 95712 65656 95776
rect 65720 95712 65736 95776
rect 65800 95712 65816 95776
rect 65880 95712 65896 95776
rect 65960 95712 65968 95776
rect 65648 95711 65968 95712
rect 96368 95776 96688 95777
rect 96368 95712 96376 95776
rect 96440 95712 96456 95776
rect 96520 95712 96536 95776
rect 96600 95712 96616 95776
rect 96680 95712 96688 95776
rect 96368 95711 96688 95712
rect 19568 95232 19888 95233
rect 19568 95168 19576 95232
rect 19640 95168 19656 95232
rect 19720 95168 19736 95232
rect 19800 95168 19816 95232
rect 19880 95168 19888 95232
rect 19568 95167 19888 95168
rect 50288 95232 50608 95233
rect 50288 95168 50296 95232
rect 50360 95168 50376 95232
rect 50440 95168 50456 95232
rect 50520 95168 50536 95232
rect 50600 95168 50608 95232
rect 50288 95167 50608 95168
rect 81008 95232 81328 95233
rect 81008 95168 81016 95232
rect 81080 95168 81096 95232
rect 81160 95168 81176 95232
rect 81240 95168 81256 95232
rect 81320 95168 81328 95232
rect 81008 95167 81328 95168
rect 4208 94688 4528 94689
rect 4208 94624 4216 94688
rect 4280 94624 4296 94688
rect 4360 94624 4376 94688
rect 4440 94624 4456 94688
rect 4520 94624 4528 94688
rect 4208 94623 4528 94624
rect 34928 94688 35248 94689
rect 34928 94624 34936 94688
rect 35000 94624 35016 94688
rect 35080 94624 35096 94688
rect 35160 94624 35176 94688
rect 35240 94624 35248 94688
rect 34928 94623 35248 94624
rect 65648 94688 65968 94689
rect 65648 94624 65656 94688
rect 65720 94624 65736 94688
rect 65800 94624 65816 94688
rect 65880 94624 65896 94688
rect 65960 94624 65968 94688
rect 65648 94623 65968 94624
rect 96368 94688 96688 94689
rect 96368 94624 96376 94688
rect 96440 94624 96456 94688
rect 96520 94624 96536 94688
rect 96600 94624 96616 94688
rect 96680 94624 96688 94688
rect 96368 94623 96688 94624
rect 19568 94144 19888 94145
rect 19568 94080 19576 94144
rect 19640 94080 19656 94144
rect 19720 94080 19736 94144
rect 19800 94080 19816 94144
rect 19880 94080 19888 94144
rect 19568 94079 19888 94080
rect 50288 94144 50608 94145
rect 50288 94080 50296 94144
rect 50360 94080 50376 94144
rect 50440 94080 50456 94144
rect 50520 94080 50536 94144
rect 50600 94080 50608 94144
rect 50288 94079 50608 94080
rect 81008 94144 81328 94145
rect 81008 94080 81016 94144
rect 81080 94080 81096 94144
rect 81160 94080 81176 94144
rect 81240 94080 81256 94144
rect 81320 94080 81328 94144
rect 81008 94079 81328 94080
rect 4208 93600 4528 93601
rect 4208 93536 4216 93600
rect 4280 93536 4296 93600
rect 4360 93536 4376 93600
rect 4440 93536 4456 93600
rect 4520 93536 4528 93600
rect 4208 93535 4528 93536
rect 34928 93600 35248 93601
rect 34928 93536 34936 93600
rect 35000 93536 35016 93600
rect 35080 93536 35096 93600
rect 35160 93536 35176 93600
rect 35240 93536 35248 93600
rect 34928 93535 35248 93536
rect 65648 93600 65968 93601
rect 65648 93536 65656 93600
rect 65720 93536 65736 93600
rect 65800 93536 65816 93600
rect 65880 93536 65896 93600
rect 65960 93536 65968 93600
rect 65648 93535 65968 93536
rect 96368 93600 96688 93601
rect 96368 93536 96376 93600
rect 96440 93536 96456 93600
rect 96520 93536 96536 93600
rect 96600 93536 96616 93600
rect 96680 93536 96688 93600
rect 96368 93535 96688 93536
rect 19568 93056 19888 93057
rect 19568 92992 19576 93056
rect 19640 92992 19656 93056
rect 19720 92992 19736 93056
rect 19800 92992 19816 93056
rect 19880 92992 19888 93056
rect 19568 92991 19888 92992
rect 50288 93056 50608 93057
rect 50288 92992 50296 93056
rect 50360 92992 50376 93056
rect 50440 92992 50456 93056
rect 50520 92992 50536 93056
rect 50600 92992 50608 93056
rect 50288 92991 50608 92992
rect 81008 93056 81328 93057
rect 81008 92992 81016 93056
rect 81080 92992 81096 93056
rect 81160 92992 81176 93056
rect 81240 92992 81256 93056
rect 81320 92992 81328 93056
rect 81008 92991 81328 92992
rect 4208 92512 4528 92513
rect 4208 92448 4216 92512
rect 4280 92448 4296 92512
rect 4360 92448 4376 92512
rect 4440 92448 4456 92512
rect 4520 92448 4528 92512
rect 4208 92447 4528 92448
rect 34928 92512 35248 92513
rect 34928 92448 34936 92512
rect 35000 92448 35016 92512
rect 35080 92448 35096 92512
rect 35160 92448 35176 92512
rect 35240 92448 35248 92512
rect 34928 92447 35248 92448
rect 65648 92512 65968 92513
rect 65648 92448 65656 92512
rect 65720 92448 65736 92512
rect 65800 92448 65816 92512
rect 65880 92448 65896 92512
rect 65960 92448 65968 92512
rect 65648 92447 65968 92448
rect 96368 92512 96688 92513
rect 96368 92448 96376 92512
rect 96440 92448 96456 92512
rect 96520 92448 96536 92512
rect 96600 92448 96616 92512
rect 96680 92448 96688 92512
rect 96368 92447 96688 92448
rect 19568 91968 19888 91969
rect 19568 91904 19576 91968
rect 19640 91904 19656 91968
rect 19720 91904 19736 91968
rect 19800 91904 19816 91968
rect 19880 91904 19888 91968
rect 19568 91903 19888 91904
rect 50288 91968 50608 91969
rect 50288 91904 50296 91968
rect 50360 91904 50376 91968
rect 50440 91904 50456 91968
rect 50520 91904 50536 91968
rect 50600 91904 50608 91968
rect 50288 91903 50608 91904
rect 81008 91968 81328 91969
rect 81008 91904 81016 91968
rect 81080 91904 81096 91968
rect 81160 91904 81176 91968
rect 81240 91904 81256 91968
rect 81320 91904 81328 91968
rect 81008 91903 81328 91904
rect 4208 91424 4528 91425
rect 4208 91360 4216 91424
rect 4280 91360 4296 91424
rect 4360 91360 4376 91424
rect 4440 91360 4456 91424
rect 4520 91360 4528 91424
rect 4208 91359 4528 91360
rect 34928 91424 35248 91425
rect 34928 91360 34936 91424
rect 35000 91360 35016 91424
rect 35080 91360 35096 91424
rect 35160 91360 35176 91424
rect 35240 91360 35248 91424
rect 34928 91359 35248 91360
rect 65648 91424 65968 91425
rect 65648 91360 65656 91424
rect 65720 91360 65736 91424
rect 65800 91360 65816 91424
rect 65880 91360 65896 91424
rect 65960 91360 65968 91424
rect 65648 91359 65968 91360
rect 96368 91424 96688 91425
rect 96368 91360 96376 91424
rect 96440 91360 96456 91424
rect 96520 91360 96536 91424
rect 96600 91360 96616 91424
rect 96680 91360 96688 91424
rect 96368 91359 96688 91360
rect 19568 90880 19888 90881
rect 19568 90816 19576 90880
rect 19640 90816 19656 90880
rect 19720 90816 19736 90880
rect 19800 90816 19816 90880
rect 19880 90816 19888 90880
rect 19568 90815 19888 90816
rect 50288 90880 50608 90881
rect 50288 90816 50296 90880
rect 50360 90816 50376 90880
rect 50440 90816 50456 90880
rect 50520 90816 50536 90880
rect 50600 90816 50608 90880
rect 50288 90815 50608 90816
rect 81008 90880 81328 90881
rect 81008 90816 81016 90880
rect 81080 90816 81096 90880
rect 81160 90816 81176 90880
rect 81240 90816 81256 90880
rect 81320 90816 81328 90880
rect 81008 90815 81328 90816
rect 4208 90336 4528 90337
rect 4208 90272 4216 90336
rect 4280 90272 4296 90336
rect 4360 90272 4376 90336
rect 4440 90272 4456 90336
rect 4520 90272 4528 90336
rect 4208 90271 4528 90272
rect 34928 90336 35248 90337
rect 34928 90272 34936 90336
rect 35000 90272 35016 90336
rect 35080 90272 35096 90336
rect 35160 90272 35176 90336
rect 35240 90272 35248 90336
rect 34928 90271 35248 90272
rect 65648 90336 65968 90337
rect 65648 90272 65656 90336
rect 65720 90272 65736 90336
rect 65800 90272 65816 90336
rect 65880 90272 65896 90336
rect 65960 90272 65968 90336
rect 65648 90271 65968 90272
rect 96368 90336 96688 90337
rect 96368 90272 96376 90336
rect 96440 90272 96456 90336
rect 96520 90272 96536 90336
rect 96600 90272 96616 90336
rect 96680 90272 96688 90336
rect 96368 90271 96688 90272
rect 19568 89792 19888 89793
rect 19568 89728 19576 89792
rect 19640 89728 19656 89792
rect 19720 89728 19736 89792
rect 19800 89728 19816 89792
rect 19880 89728 19888 89792
rect 19568 89727 19888 89728
rect 50288 89792 50608 89793
rect 50288 89728 50296 89792
rect 50360 89728 50376 89792
rect 50440 89728 50456 89792
rect 50520 89728 50536 89792
rect 50600 89728 50608 89792
rect 50288 89727 50608 89728
rect 81008 89792 81328 89793
rect 81008 89728 81016 89792
rect 81080 89728 81096 89792
rect 81160 89728 81176 89792
rect 81240 89728 81256 89792
rect 81320 89728 81328 89792
rect 81008 89727 81328 89728
rect 4208 89248 4528 89249
rect 4208 89184 4216 89248
rect 4280 89184 4296 89248
rect 4360 89184 4376 89248
rect 4440 89184 4456 89248
rect 4520 89184 4528 89248
rect 4208 89183 4528 89184
rect 34928 89248 35248 89249
rect 34928 89184 34936 89248
rect 35000 89184 35016 89248
rect 35080 89184 35096 89248
rect 35160 89184 35176 89248
rect 35240 89184 35248 89248
rect 34928 89183 35248 89184
rect 65648 89248 65968 89249
rect 65648 89184 65656 89248
rect 65720 89184 65736 89248
rect 65800 89184 65816 89248
rect 65880 89184 65896 89248
rect 65960 89184 65968 89248
rect 65648 89183 65968 89184
rect 96368 89248 96688 89249
rect 96368 89184 96376 89248
rect 96440 89184 96456 89248
rect 96520 89184 96536 89248
rect 96600 89184 96616 89248
rect 96680 89184 96688 89248
rect 96368 89183 96688 89184
rect 19568 88704 19888 88705
rect 19568 88640 19576 88704
rect 19640 88640 19656 88704
rect 19720 88640 19736 88704
rect 19800 88640 19816 88704
rect 19880 88640 19888 88704
rect 19568 88639 19888 88640
rect 50288 88704 50608 88705
rect 50288 88640 50296 88704
rect 50360 88640 50376 88704
rect 50440 88640 50456 88704
rect 50520 88640 50536 88704
rect 50600 88640 50608 88704
rect 50288 88639 50608 88640
rect 81008 88704 81328 88705
rect 81008 88640 81016 88704
rect 81080 88640 81096 88704
rect 81160 88640 81176 88704
rect 81240 88640 81256 88704
rect 81320 88640 81328 88704
rect 81008 88639 81328 88640
rect 4208 88160 4528 88161
rect 4208 88096 4216 88160
rect 4280 88096 4296 88160
rect 4360 88096 4376 88160
rect 4440 88096 4456 88160
rect 4520 88096 4528 88160
rect 4208 88095 4528 88096
rect 34928 88160 35248 88161
rect 34928 88096 34936 88160
rect 35000 88096 35016 88160
rect 35080 88096 35096 88160
rect 35160 88096 35176 88160
rect 35240 88096 35248 88160
rect 34928 88095 35248 88096
rect 65648 88160 65968 88161
rect 65648 88096 65656 88160
rect 65720 88096 65736 88160
rect 65800 88096 65816 88160
rect 65880 88096 65896 88160
rect 65960 88096 65968 88160
rect 65648 88095 65968 88096
rect 96368 88160 96688 88161
rect 96368 88096 96376 88160
rect 96440 88096 96456 88160
rect 96520 88096 96536 88160
rect 96600 88096 96616 88160
rect 96680 88096 96688 88160
rect 96368 88095 96688 88096
rect 19568 87616 19888 87617
rect 19568 87552 19576 87616
rect 19640 87552 19656 87616
rect 19720 87552 19736 87616
rect 19800 87552 19816 87616
rect 19880 87552 19888 87616
rect 19568 87551 19888 87552
rect 50288 87616 50608 87617
rect 50288 87552 50296 87616
rect 50360 87552 50376 87616
rect 50440 87552 50456 87616
rect 50520 87552 50536 87616
rect 50600 87552 50608 87616
rect 50288 87551 50608 87552
rect 81008 87616 81328 87617
rect 81008 87552 81016 87616
rect 81080 87552 81096 87616
rect 81160 87552 81176 87616
rect 81240 87552 81256 87616
rect 81320 87552 81328 87616
rect 81008 87551 81328 87552
rect 4208 87072 4528 87073
rect 4208 87008 4216 87072
rect 4280 87008 4296 87072
rect 4360 87008 4376 87072
rect 4440 87008 4456 87072
rect 4520 87008 4528 87072
rect 4208 87007 4528 87008
rect 34928 87072 35248 87073
rect 34928 87008 34936 87072
rect 35000 87008 35016 87072
rect 35080 87008 35096 87072
rect 35160 87008 35176 87072
rect 35240 87008 35248 87072
rect 34928 87007 35248 87008
rect 65648 87072 65968 87073
rect 65648 87008 65656 87072
rect 65720 87008 65736 87072
rect 65800 87008 65816 87072
rect 65880 87008 65896 87072
rect 65960 87008 65968 87072
rect 65648 87007 65968 87008
rect 96368 87072 96688 87073
rect 96368 87008 96376 87072
rect 96440 87008 96456 87072
rect 96520 87008 96536 87072
rect 96600 87008 96616 87072
rect 96680 87008 96688 87072
rect 96368 87007 96688 87008
rect 19568 86528 19888 86529
rect 19568 86464 19576 86528
rect 19640 86464 19656 86528
rect 19720 86464 19736 86528
rect 19800 86464 19816 86528
rect 19880 86464 19888 86528
rect 19568 86463 19888 86464
rect 50288 86528 50608 86529
rect 50288 86464 50296 86528
rect 50360 86464 50376 86528
rect 50440 86464 50456 86528
rect 50520 86464 50536 86528
rect 50600 86464 50608 86528
rect 50288 86463 50608 86464
rect 81008 86528 81328 86529
rect 81008 86464 81016 86528
rect 81080 86464 81096 86528
rect 81160 86464 81176 86528
rect 81240 86464 81256 86528
rect 81320 86464 81328 86528
rect 81008 86463 81328 86464
rect 4208 85984 4528 85985
rect 4208 85920 4216 85984
rect 4280 85920 4296 85984
rect 4360 85920 4376 85984
rect 4440 85920 4456 85984
rect 4520 85920 4528 85984
rect 4208 85919 4528 85920
rect 34928 85984 35248 85985
rect 34928 85920 34936 85984
rect 35000 85920 35016 85984
rect 35080 85920 35096 85984
rect 35160 85920 35176 85984
rect 35240 85920 35248 85984
rect 34928 85919 35248 85920
rect 65648 85984 65968 85985
rect 65648 85920 65656 85984
rect 65720 85920 65736 85984
rect 65800 85920 65816 85984
rect 65880 85920 65896 85984
rect 65960 85920 65968 85984
rect 65648 85919 65968 85920
rect 96368 85984 96688 85985
rect 96368 85920 96376 85984
rect 96440 85920 96456 85984
rect 96520 85920 96536 85984
rect 96600 85920 96616 85984
rect 96680 85920 96688 85984
rect 96368 85919 96688 85920
rect 19568 85440 19888 85441
rect 19568 85376 19576 85440
rect 19640 85376 19656 85440
rect 19720 85376 19736 85440
rect 19800 85376 19816 85440
rect 19880 85376 19888 85440
rect 19568 85375 19888 85376
rect 50288 85440 50608 85441
rect 50288 85376 50296 85440
rect 50360 85376 50376 85440
rect 50440 85376 50456 85440
rect 50520 85376 50536 85440
rect 50600 85376 50608 85440
rect 50288 85375 50608 85376
rect 81008 85440 81328 85441
rect 81008 85376 81016 85440
rect 81080 85376 81096 85440
rect 81160 85376 81176 85440
rect 81240 85376 81256 85440
rect 81320 85376 81328 85440
rect 81008 85375 81328 85376
rect 10041 85234 10107 85237
rect 14641 85234 14707 85237
rect 10041 85232 14707 85234
rect 10041 85176 10046 85232
rect 10102 85176 14646 85232
rect 14702 85176 14707 85232
rect 10041 85174 14707 85176
rect 10041 85171 10107 85174
rect 14641 85171 14707 85174
rect 4208 84896 4528 84897
rect 4208 84832 4216 84896
rect 4280 84832 4296 84896
rect 4360 84832 4376 84896
rect 4440 84832 4456 84896
rect 4520 84832 4528 84896
rect 4208 84831 4528 84832
rect 34928 84896 35248 84897
rect 34928 84832 34936 84896
rect 35000 84832 35016 84896
rect 35080 84832 35096 84896
rect 35160 84832 35176 84896
rect 35240 84832 35248 84896
rect 34928 84831 35248 84832
rect 65648 84896 65968 84897
rect 65648 84832 65656 84896
rect 65720 84832 65736 84896
rect 65800 84832 65816 84896
rect 65880 84832 65896 84896
rect 65960 84832 65968 84896
rect 65648 84831 65968 84832
rect 96368 84896 96688 84897
rect 96368 84832 96376 84896
rect 96440 84832 96456 84896
rect 96520 84832 96536 84896
rect 96600 84832 96616 84896
rect 96680 84832 96688 84896
rect 96368 84831 96688 84832
rect 19568 84352 19888 84353
rect 19568 84288 19576 84352
rect 19640 84288 19656 84352
rect 19720 84288 19736 84352
rect 19800 84288 19816 84352
rect 19880 84288 19888 84352
rect 19568 84287 19888 84288
rect 50288 84352 50608 84353
rect 50288 84288 50296 84352
rect 50360 84288 50376 84352
rect 50440 84288 50456 84352
rect 50520 84288 50536 84352
rect 50600 84288 50608 84352
rect 50288 84287 50608 84288
rect 81008 84352 81328 84353
rect 81008 84288 81016 84352
rect 81080 84288 81096 84352
rect 81160 84288 81176 84352
rect 81240 84288 81256 84352
rect 81320 84288 81328 84352
rect 81008 84287 81328 84288
rect 4208 83808 4528 83809
rect 4208 83744 4216 83808
rect 4280 83744 4296 83808
rect 4360 83744 4376 83808
rect 4440 83744 4456 83808
rect 4520 83744 4528 83808
rect 4208 83743 4528 83744
rect 34928 83808 35248 83809
rect 34928 83744 34936 83808
rect 35000 83744 35016 83808
rect 35080 83744 35096 83808
rect 35160 83744 35176 83808
rect 35240 83744 35248 83808
rect 34928 83743 35248 83744
rect 65648 83808 65968 83809
rect 65648 83744 65656 83808
rect 65720 83744 65736 83808
rect 65800 83744 65816 83808
rect 65880 83744 65896 83808
rect 65960 83744 65968 83808
rect 65648 83743 65968 83744
rect 96368 83808 96688 83809
rect 96368 83744 96376 83808
rect 96440 83744 96456 83808
rect 96520 83744 96536 83808
rect 96600 83744 96616 83808
rect 96680 83744 96688 83808
rect 96368 83743 96688 83744
rect 19568 83264 19888 83265
rect 19568 83200 19576 83264
rect 19640 83200 19656 83264
rect 19720 83200 19736 83264
rect 19800 83200 19816 83264
rect 19880 83200 19888 83264
rect 19568 83199 19888 83200
rect 50288 83264 50608 83265
rect 50288 83200 50296 83264
rect 50360 83200 50376 83264
rect 50440 83200 50456 83264
rect 50520 83200 50536 83264
rect 50600 83200 50608 83264
rect 50288 83199 50608 83200
rect 81008 83264 81328 83265
rect 81008 83200 81016 83264
rect 81080 83200 81096 83264
rect 81160 83200 81176 83264
rect 81240 83200 81256 83264
rect 81320 83200 81328 83264
rect 81008 83199 81328 83200
rect 4208 82720 4528 82721
rect 4208 82656 4216 82720
rect 4280 82656 4296 82720
rect 4360 82656 4376 82720
rect 4440 82656 4456 82720
rect 4520 82656 4528 82720
rect 4208 82655 4528 82656
rect 34928 82720 35248 82721
rect 34928 82656 34936 82720
rect 35000 82656 35016 82720
rect 35080 82656 35096 82720
rect 35160 82656 35176 82720
rect 35240 82656 35248 82720
rect 34928 82655 35248 82656
rect 65648 82720 65968 82721
rect 65648 82656 65656 82720
rect 65720 82656 65736 82720
rect 65800 82656 65816 82720
rect 65880 82656 65896 82720
rect 65960 82656 65968 82720
rect 65648 82655 65968 82656
rect 96368 82720 96688 82721
rect 96368 82656 96376 82720
rect 96440 82656 96456 82720
rect 96520 82656 96536 82720
rect 96600 82656 96616 82720
rect 96680 82656 96688 82720
rect 96368 82655 96688 82656
rect 19568 82176 19888 82177
rect 19568 82112 19576 82176
rect 19640 82112 19656 82176
rect 19720 82112 19736 82176
rect 19800 82112 19816 82176
rect 19880 82112 19888 82176
rect 19568 82111 19888 82112
rect 50288 82176 50608 82177
rect 50288 82112 50296 82176
rect 50360 82112 50376 82176
rect 50440 82112 50456 82176
rect 50520 82112 50536 82176
rect 50600 82112 50608 82176
rect 50288 82111 50608 82112
rect 81008 82176 81328 82177
rect 81008 82112 81016 82176
rect 81080 82112 81096 82176
rect 81160 82112 81176 82176
rect 81240 82112 81256 82176
rect 81320 82112 81328 82176
rect 81008 82111 81328 82112
rect 4208 81632 4528 81633
rect 4208 81568 4216 81632
rect 4280 81568 4296 81632
rect 4360 81568 4376 81632
rect 4440 81568 4456 81632
rect 4520 81568 4528 81632
rect 4208 81567 4528 81568
rect 34928 81632 35248 81633
rect 34928 81568 34936 81632
rect 35000 81568 35016 81632
rect 35080 81568 35096 81632
rect 35160 81568 35176 81632
rect 35240 81568 35248 81632
rect 34928 81567 35248 81568
rect 65648 81632 65968 81633
rect 65648 81568 65656 81632
rect 65720 81568 65736 81632
rect 65800 81568 65816 81632
rect 65880 81568 65896 81632
rect 65960 81568 65968 81632
rect 65648 81567 65968 81568
rect 96368 81632 96688 81633
rect 96368 81568 96376 81632
rect 96440 81568 96456 81632
rect 96520 81568 96536 81632
rect 96600 81568 96616 81632
rect 96680 81568 96688 81632
rect 96368 81567 96688 81568
rect 19568 81088 19888 81089
rect 19568 81024 19576 81088
rect 19640 81024 19656 81088
rect 19720 81024 19736 81088
rect 19800 81024 19816 81088
rect 19880 81024 19888 81088
rect 19568 81023 19888 81024
rect 50288 81088 50608 81089
rect 50288 81024 50296 81088
rect 50360 81024 50376 81088
rect 50440 81024 50456 81088
rect 50520 81024 50536 81088
rect 50600 81024 50608 81088
rect 50288 81023 50608 81024
rect 81008 81088 81328 81089
rect 81008 81024 81016 81088
rect 81080 81024 81096 81088
rect 81160 81024 81176 81088
rect 81240 81024 81256 81088
rect 81320 81024 81328 81088
rect 81008 81023 81328 81024
rect 4208 80544 4528 80545
rect 4208 80480 4216 80544
rect 4280 80480 4296 80544
rect 4360 80480 4376 80544
rect 4440 80480 4456 80544
rect 4520 80480 4528 80544
rect 4208 80479 4528 80480
rect 34928 80544 35248 80545
rect 34928 80480 34936 80544
rect 35000 80480 35016 80544
rect 35080 80480 35096 80544
rect 35160 80480 35176 80544
rect 35240 80480 35248 80544
rect 34928 80479 35248 80480
rect 65648 80544 65968 80545
rect 65648 80480 65656 80544
rect 65720 80480 65736 80544
rect 65800 80480 65816 80544
rect 65880 80480 65896 80544
rect 65960 80480 65968 80544
rect 65648 80479 65968 80480
rect 96368 80544 96688 80545
rect 96368 80480 96376 80544
rect 96440 80480 96456 80544
rect 96520 80480 96536 80544
rect 96600 80480 96616 80544
rect 96680 80480 96688 80544
rect 96368 80479 96688 80480
rect 19568 80000 19888 80001
rect 19568 79936 19576 80000
rect 19640 79936 19656 80000
rect 19720 79936 19736 80000
rect 19800 79936 19816 80000
rect 19880 79936 19888 80000
rect 19568 79935 19888 79936
rect 50288 80000 50608 80001
rect 50288 79936 50296 80000
rect 50360 79936 50376 80000
rect 50440 79936 50456 80000
rect 50520 79936 50536 80000
rect 50600 79936 50608 80000
rect 50288 79935 50608 79936
rect 81008 80000 81328 80001
rect 81008 79936 81016 80000
rect 81080 79936 81096 80000
rect 81160 79936 81176 80000
rect 81240 79936 81256 80000
rect 81320 79936 81328 80000
rect 81008 79935 81328 79936
rect 42609 79658 42675 79661
rect 43437 79658 43503 79661
rect 42609 79656 43503 79658
rect 42609 79600 42614 79656
rect 42670 79600 43442 79656
rect 43498 79600 43503 79656
rect 42609 79598 43503 79600
rect 42609 79595 42675 79598
rect 43437 79595 43503 79598
rect 4208 79456 4528 79457
rect 4208 79392 4216 79456
rect 4280 79392 4296 79456
rect 4360 79392 4376 79456
rect 4440 79392 4456 79456
rect 4520 79392 4528 79456
rect 4208 79391 4528 79392
rect 34928 79456 35248 79457
rect 34928 79392 34936 79456
rect 35000 79392 35016 79456
rect 35080 79392 35096 79456
rect 35160 79392 35176 79456
rect 35240 79392 35248 79456
rect 34928 79391 35248 79392
rect 65648 79456 65968 79457
rect 65648 79392 65656 79456
rect 65720 79392 65736 79456
rect 65800 79392 65816 79456
rect 65880 79392 65896 79456
rect 65960 79392 65968 79456
rect 65648 79391 65968 79392
rect 96368 79456 96688 79457
rect 96368 79392 96376 79456
rect 96440 79392 96456 79456
rect 96520 79392 96536 79456
rect 96600 79392 96616 79456
rect 96680 79392 96688 79456
rect 96368 79391 96688 79392
rect 19568 78912 19888 78913
rect 19568 78848 19576 78912
rect 19640 78848 19656 78912
rect 19720 78848 19736 78912
rect 19800 78848 19816 78912
rect 19880 78848 19888 78912
rect 19568 78847 19888 78848
rect 50288 78912 50608 78913
rect 50288 78848 50296 78912
rect 50360 78848 50376 78912
rect 50440 78848 50456 78912
rect 50520 78848 50536 78912
rect 50600 78848 50608 78912
rect 50288 78847 50608 78848
rect 81008 78912 81328 78913
rect 81008 78848 81016 78912
rect 81080 78848 81096 78912
rect 81160 78848 81176 78912
rect 81240 78848 81256 78912
rect 81320 78848 81328 78912
rect 81008 78847 81328 78848
rect 4208 78368 4528 78369
rect 4208 78304 4216 78368
rect 4280 78304 4296 78368
rect 4360 78304 4376 78368
rect 4440 78304 4456 78368
rect 4520 78304 4528 78368
rect 4208 78303 4528 78304
rect 34928 78368 35248 78369
rect 34928 78304 34936 78368
rect 35000 78304 35016 78368
rect 35080 78304 35096 78368
rect 35160 78304 35176 78368
rect 35240 78304 35248 78368
rect 34928 78303 35248 78304
rect 65648 78368 65968 78369
rect 65648 78304 65656 78368
rect 65720 78304 65736 78368
rect 65800 78304 65816 78368
rect 65880 78304 65896 78368
rect 65960 78304 65968 78368
rect 65648 78303 65968 78304
rect 96368 78368 96688 78369
rect 96368 78304 96376 78368
rect 96440 78304 96456 78368
rect 96520 78304 96536 78368
rect 96600 78304 96616 78368
rect 96680 78304 96688 78368
rect 96368 78303 96688 78304
rect 19568 77824 19888 77825
rect 19568 77760 19576 77824
rect 19640 77760 19656 77824
rect 19720 77760 19736 77824
rect 19800 77760 19816 77824
rect 19880 77760 19888 77824
rect 19568 77759 19888 77760
rect 50288 77824 50608 77825
rect 50288 77760 50296 77824
rect 50360 77760 50376 77824
rect 50440 77760 50456 77824
rect 50520 77760 50536 77824
rect 50600 77760 50608 77824
rect 50288 77759 50608 77760
rect 81008 77824 81328 77825
rect 81008 77760 81016 77824
rect 81080 77760 81096 77824
rect 81160 77760 81176 77824
rect 81240 77760 81256 77824
rect 81320 77760 81328 77824
rect 81008 77759 81328 77760
rect 4208 77280 4528 77281
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 77215 4528 77216
rect 34928 77280 35248 77281
rect 34928 77216 34936 77280
rect 35000 77216 35016 77280
rect 35080 77216 35096 77280
rect 35160 77216 35176 77280
rect 35240 77216 35248 77280
rect 34928 77215 35248 77216
rect 65648 77280 65968 77281
rect 65648 77216 65656 77280
rect 65720 77216 65736 77280
rect 65800 77216 65816 77280
rect 65880 77216 65896 77280
rect 65960 77216 65968 77280
rect 65648 77215 65968 77216
rect 96368 77280 96688 77281
rect 96368 77216 96376 77280
rect 96440 77216 96456 77280
rect 96520 77216 96536 77280
rect 96600 77216 96616 77280
rect 96680 77216 96688 77280
rect 96368 77215 96688 77216
rect 19568 76736 19888 76737
rect 19568 76672 19576 76736
rect 19640 76672 19656 76736
rect 19720 76672 19736 76736
rect 19800 76672 19816 76736
rect 19880 76672 19888 76736
rect 19568 76671 19888 76672
rect 50288 76736 50608 76737
rect 50288 76672 50296 76736
rect 50360 76672 50376 76736
rect 50440 76672 50456 76736
rect 50520 76672 50536 76736
rect 50600 76672 50608 76736
rect 50288 76671 50608 76672
rect 81008 76736 81328 76737
rect 81008 76672 81016 76736
rect 81080 76672 81096 76736
rect 81160 76672 81176 76736
rect 81240 76672 81256 76736
rect 81320 76672 81328 76736
rect 81008 76671 81328 76672
rect 4208 76192 4528 76193
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 76127 4528 76128
rect 34928 76192 35248 76193
rect 34928 76128 34936 76192
rect 35000 76128 35016 76192
rect 35080 76128 35096 76192
rect 35160 76128 35176 76192
rect 35240 76128 35248 76192
rect 34928 76127 35248 76128
rect 65648 76192 65968 76193
rect 65648 76128 65656 76192
rect 65720 76128 65736 76192
rect 65800 76128 65816 76192
rect 65880 76128 65896 76192
rect 65960 76128 65968 76192
rect 65648 76127 65968 76128
rect 96368 76192 96688 76193
rect 96368 76128 96376 76192
rect 96440 76128 96456 76192
rect 96520 76128 96536 76192
rect 96600 76128 96616 76192
rect 96680 76128 96688 76192
rect 96368 76127 96688 76128
rect 19568 75648 19888 75649
rect 19568 75584 19576 75648
rect 19640 75584 19656 75648
rect 19720 75584 19736 75648
rect 19800 75584 19816 75648
rect 19880 75584 19888 75648
rect 19568 75583 19888 75584
rect 50288 75648 50608 75649
rect 50288 75584 50296 75648
rect 50360 75584 50376 75648
rect 50440 75584 50456 75648
rect 50520 75584 50536 75648
rect 50600 75584 50608 75648
rect 50288 75583 50608 75584
rect 81008 75648 81328 75649
rect 81008 75584 81016 75648
rect 81080 75584 81096 75648
rect 81160 75584 81176 75648
rect 81240 75584 81256 75648
rect 81320 75584 81328 75648
rect 81008 75583 81328 75584
rect 4208 75104 4528 75105
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 75039 4528 75040
rect 34928 75104 35248 75105
rect 34928 75040 34936 75104
rect 35000 75040 35016 75104
rect 35080 75040 35096 75104
rect 35160 75040 35176 75104
rect 35240 75040 35248 75104
rect 34928 75039 35248 75040
rect 65648 75104 65968 75105
rect 65648 75040 65656 75104
rect 65720 75040 65736 75104
rect 65800 75040 65816 75104
rect 65880 75040 65896 75104
rect 65960 75040 65968 75104
rect 65648 75039 65968 75040
rect 96368 75104 96688 75105
rect 96368 75040 96376 75104
rect 96440 75040 96456 75104
rect 96520 75040 96536 75104
rect 96600 75040 96616 75104
rect 96680 75040 96688 75104
rect 96368 75039 96688 75040
rect 19568 74560 19888 74561
rect 19568 74496 19576 74560
rect 19640 74496 19656 74560
rect 19720 74496 19736 74560
rect 19800 74496 19816 74560
rect 19880 74496 19888 74560
rect 19568 74495 19888 74496
rect 50288 74560 50608 74561
rect 50288 74496 50296 74560
rect 50360 74496 50376 74560
rect 50440 74496 50456 74560
rect 50520 74496 50536 74560
rect 50600 74496 50608 74560
rect 50288 74495 50608 74496
rect 81008 74560 81328 74561
rect 81008 74496 81016 74560
rect 81080 74496 81096 74560
rect 81160 74496 81176 74560
rect 81240 74496 81256 74560
rect 81320 74496 81328 74560
rect 81008 74495 81328 74496
rect 4208 74016 4528 74017
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 73951 4528 73952
rect 34928 74016 35248 74017
rect 34928 73952 34936 74016
rect 35000 73952 35016 74016
rect 35080 73952 35096 74016
rect 35160 73952 35176 74016
rect 35240 73952 35248 74016
rect 34928 73951 35248 73952
rect 65648 74016 65968 74017
rect 65648 73952 65656 74016
rect 65720 73952 65736 74016
rect 65800 73952 65816 74016
rect 65880 73952 65896 74016
rect 65960 73952 65968 74016
rect 65648 73951 65968 73952
rect 96368 74016 96688 74017
rect 96368 73952 96376 74016
rect 96440 73952 96456 74016
rect 96520 73952 96536 74016
rect 96600 73952 96616 74016
rect 96680 73952 96688 74016
rect 96368 73951 96688 73952
rect 19568 73472 19888 73473
rect 19568 73408 19576 73472
rect 19640 73408 19656 73472
rect 19720 73408 19736 73472
rect 19800 73408 19816 73472
rect 19880 73408 19888 73472
rect 19568 73407 19888 73408
rect 50288 73472 50608 73473
rect 50288 73408 50296 73472
rect 50360 73408 50376 73472
rect 50440 73408 50456 73472
rect 50520 73408 50536 73472
rect 50600 73408 50608 73472
rect 50288 73407 50608 73408
rect 81008 73472 81328 73473
rect 81008 73408 81016 73472
rect 81080 73408 81096 73472
rect 81160 73408 81176 73472
rect 81240 73408 81256 73472
rect 81320 73408 81328 73472
rect 81008 73407 81328 73408
rect 4208 72928 4528 72929
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 72863 4528 72864
rect 34928 72928 35248 72929
rect 34928 72864 34936 72928
rect 35000 72864 35016 72928
rect 35080 72864 35096 72928
rect 35160 72864 35176 72928
rect 35240 72864 35248 72928
rect 34928 72863 35248 72864
rect 65648 72928 65968 72929
rect 65648 72864 65656 72928
rect 65720 72864 65736 72928
rect 65800 72864 65816 72928
rect 65880 72864 65896 72928
rect 65960 72864 65968 72928
rect 65648 72863 65968 72864
rect 96368 72928 96688 72929
rect 96368 72864 96376 72928
rect 96440 72864 96456 72928
rect 96520 72864 96536 72928
rect 96600 72864 96616 72928
rect 96680 72864 96688 72928
rect 96368 72863 96688 72864
rect 19568 72384 19888 72385
rect 19568 72320 19576 72384
rect 19640 72320 19656 72384
rect 19720 72320 19736 72384
rect 19800 72320 19816 72384
rect 19880 72320 19888 72384
rect 19568 72319 19888 72320
rect 50288 72384 50608 72385
rect 50288 72320 50296 72384
rect 50360 72320 50376 72384
rect 50440 72320 50456 72384
rect 50520 72320 50536 72384
rect 50600 72320 50608 72384
rect 50288 72319 50608 72320
rect 81008 72384 81328 72385
rect 81008 72320 81016 72384
rect 81080 72320 81096 72384
rect 81160 72320 81176 72384
rect 81240 72320 81256 72384
rect 81320 72320 81328 72384
rect 81008 72319 81328 72320
rect 4208 71840 4528 71841
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 71775 4528 71776
rect 34928 71840 35248 71841
rect 34928 71776 34936 71840
rect 35000 71776 35016 71840
rect 35080 71776 35096 71840
rect 35160 71776 35176 71840
rect 35240 71776 35248 71840
rect 34928 71775 35248 71776
rect 65648 71840 65968 71841
rect 65648 71776 65656 71840
rect 65720 71776 65736 71840
rect 65800 71776 65816 71840
rect 65880 71776 65896 71840
rect 65960 71776 65968 71840
rect 65648 71775 65968 71776
rect 96368 71840 96688 71841
rect 96368 71776 96376 71840
rect 96440 71776 96456 71840
rect 96520 71776 96536 71840
rect 96600 71776 96616 71840
rect 96680 71776 96688 71840
rect 96368 71775 96688 71776
rect 19568 71296 19888 71297
rect 19568 71232 19576 71296
rect 19640 71232 19656 71296
rect 19720 71232 19736 71296
rect 19800 71232 19816 71296
rect 19880 71232 19888 71296
rect 19568 71231 19888 71232
rect 50288 71296 50608 71297
rect 50288 71232 50296 71296
rect 50360 71232 50376 71296
rect 50440 71232 50456 71296
rect 50520 71232 50536 71296
rect 50600 71232 50608 71296
rect 50288 71231 50608 71232
rect 81008 71296 81328 71297
rect 81008 71232 81016 71296
rect 81080 71232 81096 71296
rect 81160 71232 81176 71296
rect 81240 71232 81256 71296
rect 81320 71232 81328 71296
rect 81008 71231 81328 71232
rect 26417 71090 26483 71093
rect 26693 71090 26759 71093
rect 26417 71088 26759 71090
rect 26417 71032 26422 71088
rect 26478 71032 26698 71088
rect 26754 71032 26759 71088
rect 26417 71030 26759 71032
rect 26417 71027 26483 71030
rect 26693 71027 26759 71030
rect 4208 70752 4528 70753
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 70687 4528 70688
rect 34928 70752 35248 70753
rect 34928 70688 34936 70752
rect 35000 70688 35016 70752
rect 35080 70688 35096 70752
rect 35160 70688 35176 70752
rect 35240 70688 35248 70752
rect 34928 70687 35248 70688
rect 65648 70752 65968 70753
rect 65648 70688 65656 70752
rect 65720 70688 65736 70752
rect 65800 70688 65816 70752
rect 65880 70688 65896 70752
rect 65960 70688 65968 70752
rect 65648 70687 65968 70688
rect 96368 70752 96688 70753
rect 96368 70688 96376 70752
rect 96440 70688 96456 70752
rect 96520 70688 96536 70752
rect 96600 70688 96616 70752
rect 96680 70688 96688 70752
rect 96368 70687 96688 70688
rect 57421 70410 57487 70413
rect 57881 70410 57947 70413
rect 57421 70408 57947 70410
rect 57421 70352 57426 70408
rect 57482 70352 57886 70408
rect 57942 70352 57947 70408
rect 57421 70350 57947 70352
rect 57421 70347 57487 70350
rect 57881 70347 57947 70350
rect 19568 70208 19888 70209
rect 19568 70144 19576 70208
rect 19640 70144 19656 70208
rect 19720 70144 19736 70208
rect 19800 70144 19816 70208
rect 19880 70144 19888 70208
rect 19568 70143 19888 70144
rect 50288 70208 50608 70209
rect 50288 70144 50296 70208
rect 50360 70144 50376 70208
rect 50440 70144 50456 70208
rect 50520 70144 50536 70208
rect 50600 70144 50608 70208
rect 50288 70143 50608 70144
rect 81008 70208 81328 70209
rect 81008 70144 81016 70208
rect 81080 70144 81096 70208
rect 81160 70144 81176 70208
rect 81240 70144 81256 70208
rect 81320 70144 81328 70208
rect 81008 70143 81328 70144
rect 4208 69664 4528 69665
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 69599 4528 69600
rect 34928 69664 35248 69665
rect 34928 69600 34936 69664
rect 35000 69600 35016 69664
rect 35080 69600 35096 69664
rect 35160 69600 35176 69664
rect 35240 69600 35248 69664
rect 34928 69599 35248 69600
rect 65648 69664 65968 69665
rect 65648 69600 65656 69664
rect 65720 69600 65736 69664
rect 65800 69600 65816 69664
rect 65880 69600 65896 69664
rect 65960 69600 65968 69664
rect 65648 69599 65968 69600
rect 96368 69664 96688 69665
rect 96368 69600 96376 69664
rect 96440 69600 96456 69664
rect 96520 69600 96536 69664
rect 96600 69600 96616 69664
rect 96680 69600 96688 69664
rect 96368 69599 96688 69600
rect 19568 69120 19888 69121
rect 19568 69056 19576 69120
rect 19640 69056 19656 69120
rect 19720 69056 19736 69120
rect 19800 69056 19816 69120
rect 19880 69056 19888 69120
rect 19568 69055 19888 69056
rect 50288 69120 50608 69121
rect 50288 69056 50296 69120
rect 50360 69056 50376 69120
rect 50440 69056 50456 69120
rect 50520 69056 50536 69120
rect 50600 69056 50608 69120
rect 50288 69055 50608 69056
rect 81008 69120 81328 69121
rect 81008 69056 81016 69120
rect 81080 69056 81096 69120
rect 81160 69056 81176 69120
rect 81240 69056 81256 69120
rect 81320 69056 81328 69120
rect 81008 69055 81328 69056
rect 4208 68576 4528 68577
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 68511 4528 68512
rect 34928 68576 35248 68577
rect 34928 68512 34936 68576
rect 35000 68512 35016 68576
rect 35080 68512 35096 68576
rect 35160 68512 35176 68576
rect 35240 68512 35248 68576
rect 34928 68511 35248 68512
rect 65648 68576 65968 68577
rect 65648 68512 65656 68576
rect 65720 68512 65736 68576
rect 65800 68512 65816 68576
rect 65880 68512 65896 68576
rect 65960 68512 65968 68576
rect 65648 68511 65968 68512
rect 96368 68576 96688 68577
rect 96368 68512 96376 68576
rect 96440 68512 96456 68576
rect 96520 68512 96536 68576
rect 96600 68512 96616 68576
rect 96680 68512 96688 68576
rect 96368 68511 96688 68512
rect 19568 68032 19888 68033
rect 19568 67968 19576 68032
rect 19640 67968 19656 68032
rect 19720 67968 19736 68032
rect 19800 67968 19816 68032
rect 19880 67968 19888 68032
rect 19568 67967 19888 67968
rect 50288 68032 50608 68033
rect 50288 67968 50296 68032
rect 50360 67968 50376 68032
rect 50440 67968 50456 68032
rect 50520 67968 50536 68032
rect 50600 67968 50608 68032
rect 50288 67967 50608 67968
rect 81008 68032 81328 68033
rect 81008 67968 81016 68032
rect 81080 67968 81096 68032
rect 81160 67968 81176 68032
rect 81240 67968 81256 68032
rect 81320 67968 81328 68032
rect 81008 67967 81328 67968
rect 4208 67488 4528 67489
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 67423 4528 67424
rect 34928 67488 35248 67489
rect 34928 67424 34936 67488
rect 35000 67424 35016 67488
rect 35080 67424 35096 67488
rect 35160 67424 35176 67488
rect 35240 67424 35248 67488
rect 34928 67423 35248 67424
rect 65648 67488 65968 67489
rect 65648 67424 65656 67488
rect 65720 67424 65736 67488
rect 65800 67424 65816 67488
rect 65880 67424 65896 67488
rect 65960 67424 65968 67488
rect 65648 67423 65968 67424
rect 96368 67488 96688 67489
rect 96368 67424 96376 67488
rect 96440 67424 96456 67488
rect 96520 67424 96536 67488
rect 96600 67424 96616 67488
rect 96680 67424 96688 67488
rect 96368 67423 96688 67424
rect 3969 67146 4035 67149
rect 5165 67146 5231 67149
rect 3969 67144 5231 67146
rect 3969 67088 3974 67144
rect 4030 67088 5170 67144
rect 5226 67088 5231 67144
rect 3969 67086 5231 67088
rect 3969 67083 4035 67086
rect 5165 67083 5231 67086
rect 19568 66944 19888 66945
rect 19568 66880 19576 66944
rect 19640 66880 19656 66944
rect 19720 66880 19736 66944
rect 19800 66880 19816 66944
rect 19880 66880 19888 66944
rect 19568 66879 19888 66880
rect 50288 66944 50608 66945
rect 50288 66880 50296 66944
rect 50360 66880 50376 66944
rect 50440 66880 50456 66944
rect 50520 66880 50536 66944
rect 50600 66880 50608 66944
rect 50288 66879 50608 66880
rect 81008 66944 81328 66945
rect 81008 66880 81016 66944
rect 81080 66880 81096 66944
rect 81160 66880 81176 66944
rect 81240 66880 81256 66944
rect 81320 66880 81328 66944
rect 81008 66879 81328 66880
rect 4208 66400 4528 66401
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 66335 4528 66336
rect 34928 66400 35248 66401
rect 34928 66336 34936 66400
rect 35000 66336 35016 66400
rect 35080 66336 35096 66400
rect 35160 66336 35176 66400
rect 35240 66336 35248 66400
rect 34928 66335 35248 66336
rect 65648 66400 65968 66401
rect 65648 66336 65656 66400
rect 65720 66336 65736 66400
rect 65800 66336 65816 66400
rect 65880 66336 65896 66400
rect 65960 66336 65968 66400
rect 65648 66335 65968 66336
rect 96368 66400 96688 66401
rect 96368 66336 96376 66400
rect 96440 66336 96456 66400
rect 96520 66336 96536 66400
rect 96600 66336 96616 66400
rect 96680 66336 96688 66400
rect 96368 66335 96688 66336
rect 19568 65856 19888 65857
rect 19568 65792 19576 65856
rect 19640 65792 19656 65856
rect 19720 65792 19736 65856
rect 19800 65792 19816 65856
rect 19880 65792 19888 65856
rect 19568 65791 19888 65792
rect 50288 65856 50608 65857
rect 50288 65792 50296 65856
rect 50360 65792 50376 65856
rect 50440 65792 50456 65856
rect 50520 65792 50536 65856
rect 50600 65792 50608 65856
rect 50288 65791 50608 65792
rect 81008 65856 81328 65857
rect 81008 65792 81016 65856
rect 81080 65792 81096 65856
rect 81160 65792 81176 65856
rect 81240 65792 81256 65856
rect 81320 65792 81328 65856
rect 81008 65791 81328 65792
rect 4208 65312 4528 65313
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 65247 4528 65248
rect 34928 65312 35248 65313
rect 34928 65248 34936 65312
rect 35000 65248 35016 65312
rect 35080 65248 35096 65312
rect 35160 65248 35176 65312
rect 35240 65248 35248 65312
rect 34928 65247 35248 65248
rect 65648 65312 65968 65313
rect 65648 65248 65656 65312
rect 65720 65248 65736 65312
rect 65800 65248 65816 65312
rect 65880 65248 65896 65312
rect 65960 65248 65968 65312
rect 65648 65247 65968 65248
rect 96368 65312 96688 65313
rect 96368 65248 96376 65312
rect 96440 65248 96456 65312
rect 96520 65248 96536 65312
rect 96600 65248 96616 65312
rect 96680 65248 96688 65312
rect 96368 65247 96688 65248
rect 19568 64768 19888 64769
rect 19568 64704 19576 64768
rect 19640 64704 19656 64768
rect 19720 64704 19736 64768
rect 19800 64704 19816 64768
rect 19880 64704 19888 64768
rect 19568 64703 19888 64704
rect 50288 64768 50608 64769
rect 50288 64704 50296 64768
rect 50360 64704 50376 64768
rect 50440 64704 50456 64768
rect 50520 64704 50536 64768
rect 50600 64704 50608 64768
rect 50288 64703 50608 64704
rect 81008 64768 81328 64769
rect 81008 64704 81016 64768
rect 81080 64704 81096 64768
rect 81160 64704 81176 64768
rect 81240 64704 81256 64768
rect 81320 64704 81328 64768
rect 81008 64703 81328 64704
rect 49417 64562 49483 64565
rect 50337 64562 50403 64565
rect 49417 64560 50403 64562
rect 49417 64504 49422 64560
rect 49478 64504 50342 64560
rect 50398 64504 50403 64560
rect 49417 64502 50403 64504
rect 49417 64499 49483 64502
rect 50337 64499 50403 64502
rect 49877 64426 49943 64429
rect 50245 64426 50311 64429
rect 49877 64424 50311 64426
rect 49877 64368 49882 64424
rect 49938 64368 50250 64424
rect 50306 64368 50311 64424
rect 49877 64366 50311 64368
rect 49877 64363 49943 64366
rect 50245 64363 50311 64366
rect 4208 64224 4528 64225
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 64159 4528 64160
rect 34928 64224 35248 64225
rect 34928 64160 34936 64224
rect 35000 64160 35016 64224
rect 35080 64160 35096 64224
rect 35160 64160 35176 64224
rect 35240 64160 35248 64224
rect 34928 64159 35248 64160
rect 65648 64224 65968 64225
rect 65648 64160 65656 64224
rect 65720 64160 65736 64224
rect 65800 64160 65816 64224
rect 65880 64160 65896 64224
rect 65960 64160 65968 64224
rect 65648 64159 65968 64160
rect 96368 64224 96688 64225
rect 96368 64160 96376 64224
rect 96440 64160 96456 64224
rect 96520 64160 96536 64224
rect 96600 64160 96616 64224
rect 96680 64160 96688 64224
rect 96368 64159 96688 64160
rect 66345 64018 66411 64021
rect 66989 64018 67055 64021
rect 67449 64018 67515 64021
rect 66345 64016 67515 64018
rect 66345 63960 66350 64016
rect 66406 63960 66994 64016
rect 67050 63960 67454 64016
rect 67510 63960 67515 64016
rect 66345 63958 67515 63960
rect 66345 63955 66411 63958
rect 66989 63955 67055 63958
rect 67449 63955 67515 63958
rect 62665 63882 62731 63885
rect 67265 63882 67331 63885
rect 62665 63880 67331 63882
rect 62665 63824 62670 63880
rect 62726 63824 67270 63880
rect 67326 63824 67331 63880
rect 62665 63822 67331 63824
rect 62665 63819 62731 63822
rect 67265 63819 67331 63822
rect 19568 63680 19888 63681
rect 19568 63616 19576 63680
rect 19640 63616 19656 63680
rect 19720 63616 19736 63680
rect 19800 63616 19816 63680
rect 19880 63616 19888 63680
rect 19568 63615 19888 63616
rect 50288 63680 50608 63681
rect 50288 63616 50296 63680
rect 50360 63616 50376 63680
rect 50440 63616 50456 63680
rect 50520 63616 50536 63680
rect 50600 63616 50608 63680
rect 50288 63615 50608 63616
rect 81008 63680 81328 63681
rect 81008 63616 81016 63680
rect 81080 63616 81096 63680
rect 81160 63616 81176 63680
rect 81240 63616 81256 63680
rect 81320 63616 81328 63680
rect 81008 63615 81328 63616
rect 4208 63136 4528 63137
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 63071 4528 63072
rect 34928 63136 35248 63137
rect 34928 63072 34936 63136
rect 35000 63072 35016 63136
rect 35080 63072 35096 63136
rect 35160 63072 35176 63136
rect 35240 63072 35248 63136
rect 34928 63071 35248 63072
rect 65648 63136 65968 63137
rect 65648 63072 65656 63136
rect 65720 63072 65736 63136
rect 65800 63072 65816 63136
rect 65880 63072 65896 63136
rect 65960 63072 65968 63136
rect 65648 63071 65968 63072
rect 96368 63136 96688 63137
rect 96368 63072 96376 63136
rect 96440 63072 96456 63136
rect 96520 63072 96536 63136
rect 96600 63072 96616 63136
rect 96680 63072 96688 63136
rect 96368 63071 96688 63072
rect 19568 62592 19888 62593
rect 19568 62528 19576 62592
rect 19640 62528 19656 62592
rect 19720 62528 19736 62592
rect 19800 62528 19816 62592
rect 19880 62528 19888 62592
rect 19568 62527 19888 62528
rect 50288 62592 50608 62593
rect 50288 62528 50296 62592
rect 50360 62528 50376 62592
rect 50440 62528 50456 62592
rect 50520 62528 50536 62592
rect 50600 62528 50608 62592
rect 50288 62527 50608 62528
rect 81008 62592 81328 62593
rect 81008 62528 81016 62592
rect 81080 62528 81096 62592
rect 81160 62528 81176 62592
rect 81240 62528 81256 62592
rect 81320 62528 81328 62592
rect 81008 62527 81328 62528
rect 4208 62048 4528 62049
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 61983 4528 61984
rect 34928 62048 35248 62049
rect 34928 61984 34936 62048
rect 35000 61984 35016 62048
rect 35080 61984 35096 62048
rect 35160 61984 35176 62048
rect 35240 61984 35248 62048
rect 34928 61983 35248 61984
rect 65648 62048 65968 62049
rect 65648 61984 65656 62048
rect 65720 61984 65736 62048
rect 65800 61984 65816 62048
rect 65880 61984 65896 62048
rect 65960 61984 65968 62048
rect 65648 61983 65968 61984
rect 96368 62048 96688 62049
rect 96368 61984 96376 62048
rect 96440 61984 96456 62048
rect 96520 61984 96536 62048
rect 96600 61984 96616 62048
rect 96680 61984 96688 62048
rect 96368 61983 96688 61984
rect 19568 61504 19888 61505
rect 19568 61440 19576 61504
rect 19640 61440 19656 61504
rect 19720 61440 19736 61504
rect 19800 61440 19816 61504
rect 19880 61440 19888 61504
rect 19568 61439 19888 61440
rect 50288 61504 50608 61505
rect 50288 61440 50296 61504
rect 50360 61440 50376 61504
rect 50440 61440 50456 61504
rect 50520 61440 50536 61504
rect 50600 61440 50608 61504
rect 50288 61439 50608 61440
rect 81008 61504 81328 61505
rect 81008 61440 81016 61504
rect 81080 61440 81096 61504
rect 81160 61440 81176 61504
rect 81240 61440 81256 61504
rect 81320 61440 81328 61504
rect 81008 61439 81328 61440
rect 4208 60960 4528 60961
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 60895 4528 60896
rect 34928 60960 35248 60961
rect 34928 60896 34936 60960
rect 35000 60896 35016 60960
rect 35080 60896 35096 60960
rect 35160 60896 35176 60960
rect 35240 60896 35248 60960
rect 34928 60895 35248 60896
rect 65648 60960 65968 60961
rect 65648 60896 65656 60960
rect 65720 60896 65736 60960
rect 65800 60896 65816 60960
rect 65880 60896 65896 60960
rect 65960 60896 65968 60960
rect 65648 60895 65968 60896
rect 96368 60960 96688 60961
rect 96368 60896 96376 60960
rect 96440 60896 96456 60960
rect 96520 60896 96536 60960
rect 96600 60896 96616 60960
rect 96680 60896 96688 60960
rect 96368 60895 96688 60896
rect 19568 60416 19888 60417
rect 19568 60352 19576 60416
rect 19640 60352 19656 60416
rect 19720 60352 19736 60416
rect 19800 60352 19816 60416
rect 19880 60352 19888 60416
rect 19568 60351 19888 60352
rect 50288 60416 50608 60417
rect 50288 60352 50296 60416
rect 50360 60352 50376 60416
rect 50440 60352 50456 60416
rect 50520 60352 50536 60416
rect 50600 60352 50608 60416
rect 50288 60351 50608 60352
rect 81008 60416 81328 60417
rect 81008 60352 81016 60416
rect 81080 60352 81096 60416
rect 81160 60352 81176 60416
rect 81240 60352 81256 60416
rect 81320 60352 81328 60416
rect 81008 60351 81328 60352
rect 4208 59872 4528 59873
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 59807 4528 59808
rect 34928 59872 35248 59873
rect 34928 59808 34936 59872
rect 35000 59808 35016 59872
rect 35080 59808 35096 59872
rect 35160 59808 35176 59872
rect 35240 59808 35248 59872
rect 34928 59807 35248 59808
rect 65648 59872 65968 59873
rect 65648 59808 65656 59872
rect 65720 59808 65736 59872
rect 65800 59808 65816 59872
rect 65880 59808 65896 59872
rect 65960 59808 65968 59872
rect 65648 59807 65968 59808
rect 96368 59872 96688 59873
rect 96368 59808 96376 59872
rect 96440 59808 96456 59872
rect 96520 59808 96536 59872
rect 96600 59808 96616 59872
rect 96680 59808 96688 59872
rect 96368 59807 96688 59808
rect 19568 59328 19888 59329
rect 19568 59264 19576 59328
rect 19640 59264 19656 59328
rect 19720 59264 19736 59328
rect 19800 59264 19816 59328
rect 19880 59264 19888 59328
rect 19568 59263 19888 59264
rect 50288 59328 50608 59329
rect 50288 59264 50296 59328
rect 50360 59264 50376 59328
rect 50440 59264 50456 59328
rect 50520 59264 50536 59328
rect 50600 59264 50608 59328
rect 50288 59263 50608 59264
rect 81008 59328 81328 59329
rect 81008 59264 81016 59328
rect 81080 59264 81096 59328
rect 81160 59264 81176 59328
rect 81240 59264 81256 59328
rect 81320 59264 81328 59328
rect 81008 59263 81328 59264
rect 4208 58784 4528 58785
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 58719 4528 58720
rect 34928 58784 35248 58785
rect 34928 58720 34936 58784
rect 35000 58720 35016 58784
rect 35080 58720 35096 58784
rect 35160 58720 35176 58784
rect 35240 58720 35248 58784
rect 34928 58719 35248 58720
rect 65648 58784 65968 58785
rect 65648 58720 65656 58784
rect 65720 58720 65736 58784
rect 65800 58720 65816 58784
rect 65880 58720 65896 58784
rect 65960 58720 65968 58784
rect 65648 58719 65968 58720
rect 96368 58784 96688 58785
rect 96368 58720 96376 58784
rect 96440 58720 96456 58784
rect 96520 58720 96536 58784
rect 96600 58720 96616 58784
rect 96680 58720 96688 58784
rect 96368 58719 96688 58720
rect 19568 58240 19888 58241
rect 19568 58176 19576 58240
rect 19640 58176 19656 58240
rect 19720 58176 19736 58240
rect 19800 58176 19816 58240
rect 19880 58176 19888 58240
rect 19568 58175 19888 58176
rect 50288 58240 50608 58241
rect 50288 58176 50296 58240
rect 50360 58176 50376 58240
rect 50440 58176 50456 58240
rect 50520 58176 50536 58240
rect 50600 58176 50608 58240
rect 50288 58175 50608 58176
rect 81008 58240 81328 58241
rect 81008 58176 81016 58240
rect 81080 58176 81096 58240
rect 81160 58176 81176 58240
rect 81240 58176 81256 58240
rect 81320 58176 81328 58240
rect 81008 58175 81328 58176
rect 4208 57696 4528 57697
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 57631 4528 57632
rect 34928 57696 35248 57697
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 57631 35248 57632
rect 65648 57696 65968 57697
rect 65648 57632 65656 57696
rect 65720 57632 65736 57696
rect 65800 57632 65816 57696
rect 65880 57632 65896 57696
rect 65960 57632 65968 57696
rect 65648 57631 65968 57632
rect 96368 57696 96688 57697
rect 96368 57632 96376 57696
rect 96440 57632 96456 57696
rect 96520 57632 96536 57696
rect 96600 57632 96616 57696
rect 96680 57632 96688 57696
rect 96368 57631 96688 57632
rect 19568 57152 19888 57153
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 57087 19888 57088
rect 50288 57152 50608 57153
rect 50288 57088 50296 57152
rect 50360 57088 50376 57152
rect 50440 57088 50456 57152
rect 50520 57088 50536 57152
rect 50600 57088 50608 57152
rect 50288 57087 50608 57088
rect 81008 57152 81328 57153
rect 81008 57088 81016 57152
rect 81080 57088 81096 57152
rect 81160 57088 81176 57152
rect 81240 57088 81256 57152
rect 81320 57088 81328 57152
rect 81008 57087 81328 57088
rect 4208 56608 4528 56609
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 56543 4528 56544
rect 34928 56608 35248 56609
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 56543 35248 56544
rect 65648 56608 65968 56609
rect 65648 56544 65656 56608
rect 65720 56544 65736 56608
rect 65800 56544 65816 56608
rect 65880 56544 65896 56608
rect 65960 56544 65968 56608
rect 65648 56543 65968 56544
rect 96368 56608 96688 56609
rect 96368 56544 96376 56608
rect 96440 56544 96456 56608
rect 96520 56544 96536 56608
rect 96600 56544 96616 56608
rect 96680 56544 96688 56608
rect 96368 56543 96688 56544
rect 19568 56064 19888 56065
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 55999 19888 56000
rect 50288 56064 50608 56065
rect 50288 56000 50296 56064
rect 50360 56000 50376 56064
rect 50440 56000 50456 56064
rect 50520 56000 50536 56064
rect 50600 56000 50608 56064
rect 50288 55999 50608 56000
rect 81008 56064 81328 56065
rect 81008 56000 81016 56064
rect 81080 56000 81096 56064
rect 81160 56000 81176 56064
rect 81240 56000 81256 56064
rect 81320 56000 81328 56064
rect 81008 55999 81328 56000
rect 4208 55520 4528 55521
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 55455 4528 55456
rect 34928 55520 35248 55521
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 55455 35248 55456
rect 65648 55520 65968 55521
rect 65648 55456 65656 55520
rect 65720 55456 65736 55520
rect 65800 55456 65816 55520
rect 65880 55456 65896 55520
rect 65960 55456 65968 55520
rect 65648 55455 65968 55456
rect 96368 55520 96688 55521
rect 96368 55456 96376 55520
rect 96440 55456 96456 55520
rect 96520 55456 96536 55520
rect 96600 55456 96616 55520
rect 96680 55456 96688 55520
rect 96368 55455 96688 55456
rect 19568 54976 19888 54977
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 54911 19888 54912
rect 50288 54976 50608 54977
rect 50288 54912 50296 54976
rect 50360 54912 50376 54976
rect 50440 54912 50456 54976
rect 50520 54912 50536 54976
rect 50600 54912 50608 54976
rect 50288 54911 50608 54912
rect 81008 54976 81328 54977
rect 81008 54912 81016 54976
rect 81080 54912 81096 54976
rect 81160 54912 81176 54976
rect 81240 54912 81256 54976
rect 81320 54912 81328 54976
rect 81008 54911 81328 54912
rect 4208 54432 4528 54433
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 54367 4528 54368
rect 34928 54432 35248 54433
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 54367 35248 54368
rect 65648 54432 65968 54433
rect 65648 54368 65656 54432
rect 65720 54368 65736 54432
rect 65800 54368 65816 54432
rect 65880 54368 65896 54432
rect 65960 54368 65968 54432
rect 65648 54367 65968 54368
rect 96368 54432 96688 54433
rect 96368 54368 96376 54432
rect 96440 54368 96456 54432
rect 96520 54368 96536 54432
rect 96600 54368 96616 54432
rect 96680 54368 96688 54432
rect 96368 54367 96688 54368
rect 19568 53888 19888 53889
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 53823 19888 53824
rect 50288 53888 50608 53889
rect 50288 53824 50296 53888
rect 50360 53824 50376 53888
rect 50440 53824 50456 53888
rect 50520 53824 50536 53888
rect 50600 53824 50608 53888
rect 50288 53823 50608 53824
rect 81008 53888 81328 53889
rect 81008 53824 81016 53888
rect 81080 53824 81096 53888
rect 81160 53824 81176 53888
rect 81240 53824 81256 53888
rect 81320 53824 81328 53888
rect 81008 53823 81328 53824
rect 4208 53344 4528 53345
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 53279 4528 53280
rect 34928 53344 35248 53345
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 53279 35248 53280
rect 65648 53344 65968 53345
rect 65648 53280 65656 53344
rect 65720 53280 65736 53344
rect 65800 53280 65816 53344
rect 65880 53280 65896 53344
rect 65960 53280 65968 53344
rect 65648 53279 65968 53280
rect 96368 53344 96688 53345
rect 96368 53280 96376 53344
rect 96440 53280 96456 53344
rect 96520 53280 96536 53344
rect 96600 53280 96616 53344
rect 96680 53280 96688 53344
rect 96368 53279 96688 53280
rect 19568 52800 19888 52801
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 52735 19888 52736
rect 50288 52800 50608 52801
rect 50288 52736 50296 52800
rect 50360 52736 50376 52800
rect 50440 52736 50456 52800
rect 50520 52736 50536 52800
rect 50600 52736 50608 52800
rect 50288 52735 50608 52736
rect 81008 52800 81328 52801
rect 81008 52736 81016 52800
rect 81080 52736 81096 52800
rect 81160 52736 81176 52800
rect 81240 52736 81256 52800
rect 81320 52736 81328 52800
rect 81008 52735 81328 52736
rect 4208 52256 4528 52257
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 52191 4528 52192
rect 34928 52256 35248 52257
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 52191 35248 52192
rect 65648 52256 65968 52257
rect 65648 52192 65656 52256
rect 65720 52192 65736 52256
rect 65800 52192 65816 52256
rect 65880 52192 65896 52256
rect 65960 52192 65968 52256
rect 65648 52191 65968 52192
rect 96368 52256 96688 52257
rect 96368 52192 96376 52256
rect 96440 52192 96456 52256
rect 96520 52192 96536 52256
rect 96600 52192 96616 52256
rect 96680 52192 96688 52256
rect 96368 52191 96688 52192
rect 19568 51712 19888 51713
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 51647 19888 51648
rect 50288 51712 50608 51713
rect 50288 51648 50296 51712
rect 50360 51648 50376 51712
rect 50440 51648 50456 51712
rect 50520 51648 50536 51712
rect 50600 51648 50608 51712
rect 50288 51647 50608 51648
rect 81008 51712 81328 51713
rect 81008 51648 81016 51712
rect 81080 51648 81096 51712
rect 81160 51648 81176 51712
rect 81240 51648 81256 51712
rect 81320 51648 81328 51712
rect 81008 51647 81328 51648
rect 4208 51168 4528 51169
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 51103 4528 51104
rect 34928 51168 35248 51169
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 51103 35248 51104
rect 65648 51168 65968 51169
rect 65648 51104 65656 51168
rect 65720 51104 65736 51168
rect 65800 51104 65816 51168
rect 65880 51104 65896 51168
rect 65960 51104 65968 51168
rect 65648 51103 65968 51104
rect 96368 51168 96688 51169
rect 96368 51104 96376 51168
rect 96440 51104 96456 51168
rect 96520 51104 96536 51168
rect 96600 51104 96616 51168
rect 96680 51104 96688 51168
rect 96368 51103 96688 51104
rect 19568 50624 19888 50625
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 50559 19888 50560
rect 50288 50624 50608 50625
rect 50288 50560 50296 50624
rect 50360 50560 50376 50624
rect 50440 50560 50456 50624
rect 50520 50560 50536 50624
rect 50600 50560 50608 50624
rect 50288 50559 50608 50560
rect 81008 50624 81328 50625
rect 81008 50560 81016 50624
rect 81080 50560 81096 50624
rect 81160 50560 81176 50624
rect 81240 50560 81256 50624
rect 81320 50560 81328 50624
rect 81008 50559 81328 50560
rect 4208 50080 4528 50081
rect 0 50010 800 50040
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 50015 4528 50016
rect 34928 50080 35248 50081
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 50015 35248 50016
rect 65648 50080 65968 50081
rect 65648 50016 65656 50080
rect 65720 50016 65736 50080
rect 65800 50016 65816 50080
rect 65880 50016 65896 50080
rect 65960 50016 65968 50080
rect 65648 50015 65968 50016
rect 96368 50080 96688 50081
rect 96368 50016 96376 50080
rect 96440 50016 96456 50080
rect 96520 50016 96536 50080
rect 96600 50016 96616 50080
rect 96680 50016 96688 50080
rect 96368 50015 96688 50016
rect 1393 50010 1459 50013
rect 0 50008 1459 50010
rect 0 49952 1398 50008
rect 1454 49952 1459 50008
rect 0 49950 1459 49952
rect 0 49920 800 49950
rect 1393 49947 1459 49950
rect 19568 49536 19888 49537
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 49471 19888 49472
rect 50288 49536 50608 49537
rect 50288 49472 50296 49536
rect 50360 49472 50376 49536
rect 50440 49472 50456 49536
rect 50520 49472 50536 49536
rect 50600 49472 50608 49536
rect 50288 49471 50608 49472
rect 81008 49536 81328 49537
rect 81008 49472 81016 49536
rect 81080 49472 81096 49536
rect 81160 49472 81176 49536
rect 81240 49472 81256 49536
rect 81320 49472 81328 49536
rect 81008 49471 81328 49472
rect 4208 48992 4528 48993
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 48927 4528 48928
rect 34928 48992 35248 48993
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 48927 35248 48928
rect 65648 48992 65968 48993
rect 65648 48928 65656 48992
rect 65720 48928 65736 48992
rect 65800 48928 65816 48992
rect 65880 48928 65896 48992
rect 65960 48928 65968 48992
rect 65648 48927 65968 48928
rect 96368 48992 96688 48993
rect 96368 48928 96376 48992
rect 96440 48928 96456 48992
rect 96520 48928 96536 48992
rect 96600 48928 96616 48992
rect 96680 48928 96688 48992
rect 96368 48927 96688 48928
rect 19568 48448 19888 48449
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 48383 19888 48384
rect 50288 48448 50608 48449
rect 50288 48384 50296 48448
rect 50360 48384 50376 48448
rect 50440 48384 50456 48448
rect 50520 48384 50536 48448
rect 50600 48384 50608 48448
rect 50288 48383 50608 48384
rect 81008 48448 81328 48449
rect 81008 48384 81016 48448
rect 81080 48384 81096 48448
rect 81160 48384 81176 48448
rect 81240 48384 81256 48448
rect 81320 48384 81328 48448
rect 81008 48383 81328 48384
rect 4208 47904 4528 47905
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 34928 47904 35248 47905
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 47839 35248 47840
rect 65648 47904 65968 47905
rect 65648 47840 65656 47904
rect 65720 47840 65736 47904
rect 65800 47840 65816 47904
rect 65880 47840 65896 47904
rect 65960 47840 65968 47904
rect 65648 47839 65968 47840
rect 96368 47904 96688 47905
rect 96368 47840 96376 47904
rect 96440 47840 96456 47904
rect 96520 47840 96536 47904
rect 96600 47840 96616 47904
rect 96680 47840 96688 47904
rect 96368 47839 96688 47840
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 50288 47360 50608 47361
rect 50288 47296 50296 47360
rect 50360 47296 50376 47360
rect 50440 47296 50456 47360
rect 50520 47296 50536 47360
rect 50600 47296 50608 47360
rect 50288 47295 50608 47296
rect 81008 47360 81328 47361
rect 81008 47296 81016 47360
rect 81080 47296 81096 47360
rect 81160 47296 81176 47360
rect 81240 47296 81256 47360
rect 81320 47296 81328 47360
rect 81008 47295 81328 47296
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 65648 46816 65968 46817
rect 65648 46752 65656 46816
rect 65720 46752 65736 46816
rect 65800 46752 65816 46816
rect 65880 46752 65896 46816
rect 65960 46752 65968 46816
rect 65648 46751 65968 46752
rect 96368 46816 96688 46817
rect 96368 46752 96376 46816
rect 96440 46752 96456 46816
rect 96520 46752 96536 46816
rect 96600 46752 96616 46816
rect 96680 46752 96688 46816
rect 96368 46751 96688 46752
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 50288 46272 50608 46273
rect 50288 46208 50296 46272
rect 50360 46208 50376 46272
rect 50440 46208 50456 46272
rect 50520 46208 50536 46272
rect 50600 46208 50608 46272
rect 50288 46207 50608 46208
rect 81008 46272 81328 46273
rect 81008 46208 81016 46272
rect 81080 46208 81096 46272
rect 81160 46208 81176 46272
rect 81240 46208 81256 46272
rect 81320 46208 81328 46272
rect 81008 46207 81328 46208
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 65648 45728 65968 45729
rect 65648 45664 65656 45728
rect 65720 45664 65736 45728
rect 65800 45664 65816 45728
rect 65880 45664 65896 45728
rect 65960 45664 65968 45728
rect 65648 45663 65968 45664
rect 96368 45728 96688 45729
rect 96368 45664 96376 45728
rect 96440 45664 96456 45728
rect 96520 45664 96536 45728
rect 96600 45664 96616 45728
rect 96680 45664 96688 45728
rect 96368 45663 96688 45664
rect 19568 45184 19888 45185
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 50288 45184 50608 45185
rect 50288 45120 50296 45184
rect 50360 45120 50376 45184
rect 50440 45120 50456 45184
rect 50520 45120 50536 45184
rect 50600 45120 50608 45184
rect 50288 45119 50608 45120
rect 81008 45184 81328 45185
rect 81008 45120 81016 45184
rect 81080 45120 81096 45184
rect 81160 45120 81176 45184
rect 81240 45120 81256 45184
rect 81320 45120 81328 45184
rect 81008 45119 81328 45120
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 65648 44640 65968 44641
rect 65648 44576 65656 44640
rect 65720 44576 65736 44640
rect 65800 44576 65816 44640
rect 65880 44576 65896 44640
rect 65960 44576 65968 44640
rect 65648 44575 65968 44576
rect 96368 44640 96688 44641
rect 96368 44576 96376 44640
rect 96440 44576 96456 44640
rect 96520 44576 96536 44640
rect 96600 44576 96616 44640
rect 96680 44576 96688 44640
rect 96368 44575 96688 44576
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 50288 44096 50608 44097
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 44031 50608 44032
rect 81008 44096 81328 44097
rect 81008 44032 81016 44096
rect 81080 44032 81096 44096
rect 81160 44032 81176 44096
rect 81240 44032 81256 44096
rect 81320 44032 81328 44096
rect 81008 44031 81328 44032
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 65648 43552 65968 43553
rect 65648 43488 65656 43552
rect 65720 43488 65736 43552
rect 65800 43488 65816 43552
rect 65880 43488 65896 43552
rect 65960 43488 65968 43552
rect 65648 43487 65968 43488
rect 96368 43552 96688 43553
rect 96368 43488 96376 43552
rect 96440 43488 96456 43552
rect 96520 43488 96536 43552
rect 96600 43488 96616 43552
rect 96680 43488 96688 43552
rect 96368 43487 96688 43488
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 50288 43008 50608 43009
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 42943 50608 42944
rect 81008 43008 81328 43009
rect 81008 42944 81016 43008
rect 81080 42944 81096 43008
rect 81160 42944 81176 43008
rect 81240 42944 81256 43008
rect 81320 42944 81328 43008
rect 81008 42943 81328 42944
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 65648 42464 65968 42465
rect 65648 42400 65656 42464
rect 65720 42400 65736 42464
rect 65800 42400 65816 42464
rect 65880 42400 65896 42464
rect 65960 42400 65968 42464
rect 65648 42399 65968 42400
rect 96368 42464 96688 42465
rect 96368 42400 96376 42464
rect 96440 42400 96456 42464
rect 96520 42400 96536 42464
rect 96600 42400 96616 42464
rect 96680 42400 96688 42464
rect 96368 42399 96688 42400
rect 19568 41920 19888 41921
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 50288 41920 50608 41921
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 41855 50608 41856
rect 81008 41920 81328 41921
rect 81008 41856 81016 41920
rect 81080 41856 81096 41920
rect 81160 41856 81176 41920
rect 81240 41856 81256 41920
rect 81320 41856 81328 41920
rect 81008 41855 81328 41856
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 65648 41376 65968 41377
rect 65648 41312 65656 41376
rect 65720 41312 65736 41376
rect 65800 41312 65816 41376
rect 65880 41312 65896 41376
rect 65960 41312 65968 41376
rect 65648 41311 65968 41312
rect 96368 41376 96688 41377
rect 96368 41312 96376 41376
rect 96440 41312 96456 41376
rect 96520 41312 96536 41376
rect 96600 41312 96616 41376
rect 96680 41312 96688 41376
rect 96368 41311 96688 41312
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 50288 40832 50608 40833
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 40767 50608 40768
rect 81008 40832 81328 40833
rect 81008 40768 81016 40832
rect 81080 40768 81096 40832
rect 81160 40768 81176 40832
rect 81240 40768 81256 40832
rect 81320 40768 81328 40832
rect 81008 40767 81328 40768
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 65648 40288 65968 40289
rect 65648 40224 65656 40288
rect 65720 40224 65736 40288
rect 65800 40224 65816 40288
rect 65880 40224 65896 40288
rect 65960 40224 65968 40288
rect 65648 40223 65968 40224
rect 96368 40288 96688 40289
rect 96368 40224 96376 40288
rect 96440 40224 96456 40288
rect 96520 40224 96536 40288
rect 96600 40224 96616 40288
rect 96680 40224 96688 40288
rect 96368 40223 96688 40224
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 50288 39744 50608 39745
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 39679 50608 39680
rect 81008 39744 81328 39745
rect 81008 39680 81016 39744
rect 81080 39680 81096 39744
rect 81160 39680 81176 39744
rect 81240 39680 81256 39744
rect 81320 39680 81328 39744
rect 81008 39679 81328 39680
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 65648 39200 65968 39201
rect 65648 39136 65656 39200
rect 65720 39136 65736 39200
rect 65800 39136 65816 39200
rect 65880 39136 65896 39200
rect 65960 39136 65968 39200
rect 65648 39135 65968 39136
rect 96368 39200 96688 39201
rect 96368 39136 96376 39200
rect 96440 39136 96456 39200
rect 96520 39136 96536 39200
rect 96600 39136 96616 39200
rect 96680 39136 96688 39200
rect 96368 39135 96688 39136
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 50288 38656 50608 38657
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 38591 50608 38592
rect 81008 38656 81328 38657
rect 81008 38592 81016 38656
rect 81080 38592 81096 38656
rect 81160 38592 81176 38656
rect 81240 38592 81256 38656
rect 81320 38592 81328 38656
rect 81008 38591 81328 38592
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 65648 38112 65968 38113
rect 65648 38048 65656 38112
rect 65720 38048 65736 38112
rect 65800 38048 65816 38112
rect 65880 38048 65896 38112
rect 65960 38048 65968 38112
rect 65648 38047 65968 38048
rect 96368 38112 96688 38113
rect 96368 38048 96376 38112
rect 96440 38048 96456 38112
rect 96520 38048 96536 38112
rect 96600 38048 96616 38112
rect 96680 38048 96688 38112
rect 96368 38047 96688 38048
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 50288 37568 50608 37569
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 37503 50608 37504
rect 81008 37568 81328 37569
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 37503 81328 37504
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 65648 37024 65968 37025
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 36959 65968 36960
rect 96368 37024 96688 37025
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 36959 96688 36960
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 50288 36480 50608 36481
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 36415 50608 36416
rect 81008 36480 81328 36481
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 36415 81328 36416
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 65648 35936 65968 35937
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 35871 65968 35872
rect 96368 35936 96688 35937
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 35871 96688 35872
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 50288 35392 50608 35393
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 35327 50608 35328
rect 81008 35392 81328 35393
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 35327 81328 35328
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 65648 34848 65968 34849
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 34783 65968 34784
rect 96368 34848 96688 34849
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 34783 96688 34784
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 50288 34304 50608 34305
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 34239 50608 34240
rect 81008 34304 81328 34305
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 34239 81328 34240
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 65648 33760 65968 33761
rect 65648 33696 65656 33760
rect 65720 33696 65736 33760
rect 65800 33696 65816 33760
rect 65880 33696 65896 33760
rect 65960 33696 65968 33760
rect 65648 33695 65968 33696
rect 96368 33760 96688 33761
rect 96368 33696 96376 33760
rect 96440 33696 96456 33760
rect 96520 33696 96536 33760
rect 96600 33696 96616 33760
rect 96680 33696 96688 33760
rect 96368 33695 96688 33696
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 50288 33216 50608 33217
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 33151 50608 33152
rect 81008 33216 81328 33217
rect 81008 33152 81016 33216
rect 81080 33152 81096 33216
rect 81160 33152 81176 33216
rect 81240 33152 81256 33216
rect 81320 33152 81328 33216
rect 81008 33151 81328 33152
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 65648 32672 65968 32673
rect 65648 32608 65656 32672
rect 65720 32608 65736 32672
rect 65800 32608 65816 32672
rect 65880 32608 65896 32672
rect 65960 32608 65968 32672
rect 65648 32607 65968 32608
rect 96368 32672 96688 32673
rect 96368 32608 96376 32672
rect 96440 32608 96456 32672
rect 96520 32608 96536 32672
rect 96600 32608 96616 32672
rect 96680 32608 96688 32672
rect 96368 32607 96688 32608
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 50288 32128 50608 32129
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 32063 50608 32064
rect 81008 32128 81328 32129
rect 81008 32064 81016 32128
rect 81080 32064 81096 32128
rect 81160 32064 81176 32128
rect 81240 32064 81256 32128
rect 81320 32064 81328 32128
rect 81008 32063 81328 32064
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 65648 31584 65968 31585
rect 65648 31520 65656 31584
rect 65720 31520 65736 31584
rect 65800 31520 65816 31584
rect 65880 31520 65896 31584
rect 65960 31520 65968 31584
rect 65648 31519 65968 31520
rect 96368 31584 96688 31585
rect 96368 31520 96376 31584
rect 96440 31520 96456 31584
rect 96520 31520 96536 31584
rect 96600 31520 96616 31584
rect 96680 31520 96688 31584
rect 96368 31519 96688 31520
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 50288 31040 50608 31041
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 30975 50608 30976
rect 81008 31040 81328 31041
rect 81008 30976 81016 31040
rect 81080 30976 81096 31040
rect 81160 30976 81176 31040
rect 81240 30976 81256 31040
rect 81320 30976 81328 31040
rect 81008 30975 81328 30976
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 65648 30496 65968 30497
rect 65648 30432 65656 30496
rect 65720 30432 65736 30496
rect 65800 30432 65816 30496
rect 65880 30432 65896 30496
rect 65960 30432 65968 30496
rect 65648 30431 65968 30432
rect 96368 30496 96688 30497
rect 96368 30432 96376 30496
rect 96440 30432 96456 30496
rect 96520 30432 96536 30496
rect 96600 30432 96616 30496
rect 96680 30432 96688 30496
rect 96368 30431 96688 30432
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 50288 29952 50608 29953
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 29887 50608 29888
rect 81008 29952 81328 29953
rect 81008 29888 81016 29952
rect 81080 29888 81096 29952
rect 81160 29888 81176 29952
rect 81240 29888 81256 29952
rect 81320 29888 81328 29952
rect 81008 29887 81328 29888
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 65648 29408 65968 29409
rect 65648 29344 65656 29408
rect 65720 29344 65736 29408
rect 65800 29344 65816 29408
rect 65880 29344 65896 29408
rect 65960 29344 65968 29408
rect 65648 29343 65968 29344
rect 96368 29408 96688 29409
rect 96368 29344 96376 29408
rect 96440 29344 96456 29408
rect 96520 29344 96536 29408
rect 96600 29344 96616 29408
rect 96680 29344 96688 29408
rect 96368 29343 96688 29344
rect 25681 29066 25747 29069
rect 26509 29066 26575 29069
rect 25681 29064 26575 29066
rect 25681 29008 25686 29064
rect 25742 29008 26514 29064
rect 26570 29008 26575 29064
rect 25681 29006 26575 29008
rect 25681 29003 25747 29006
rect 26509 29003 26575 29006
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 50288 28864 50608 28865
rect 50288 28800 50296 28864
rect 50360 28800 50376 28864
rect 50440 28800 50456 28864
rect 50520 28800 50536 28864
rect 50600 28800 50608 28864
rect 50288 28799 50608 28800
rect 81008 28864 81328 28865
rect 81008 28800 81016 28864
rect 81080 28800 81096 28864
rect 81160 28800 81176 28864
rect 81240 28800 81256 28864
rect 81320 28800 81328 28864
rect 81008 28799 81328 28800
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 65648 28320 65968 28321
rect 65648 28256 65656 28320
rect 65720 28256 65736 28320
rect 65800 28256 65816 28320
rect 65880 28256 65896 28320
rect 65960 28256 65968 28320
rect 65648 28255 65968 28256
rect 96368 28320 96688 28321
rect 96368 28256 96376 28320
rect 96440 28256 96456 28320
rect 96520 28256 96536 28320
rect 96600 28256 96616 28320
rect 96680 28256 96688 28320
rect 96368 28255 96688 28256
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 50288 27776 50608 27777
rect 50288 27712 50296 27776
rect 50360 27712 50376 27776
rect 50440 27712 50456 27776
rect 50520 27712 50536 27776
rect 50600 27712 50608 27776
rect 50288 27711 50608 27712
rect 81008 27776 81328 27777
rect 81008 27712 81016 27776
rect 81080 27712 81096 27776
rect 81160 27712 81176 27776
rect 81240 27712 81256 27776
rect 81320 27712 81328 27776
rect 81008 27711 81328 27712
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 65648 27232 65968 27233
rect 65648 27168 65656 27232
rect 65720 27168 65736 27232
rect 65800 27168 65816 27232
rect 65880 27168 65896 27232
rect 65960 27168 65968 27232
rect 65648 27167 65968 27168
rect 96368 27232 96688 27233
rect 96368 27168 96376 27232
rect 96440 27168 96456 27232
rect 96520 27168 96536 27232
rect 96600 27168 96616 27232
rect 96680 27168 96688 27232
rect 96368 27167 96688 27168
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 50288 26688 50608 26689
rect 50288 26624 50296 26688
rect 50360 26624 50376 26688
rect 50440 26624 50456 26688
rect 50520 26624 50536 26688
rect 50600 26624 50608 26688
rect 50288 26623 50608 26624
rect 81008 26688 81328 26689
rect 81008 26624 81016 26688
rect 81080 26624 81096 26688
rect 81160 26624 81176 26688
rect 81240 26624 81256 26688
rect 81320 26624 81328 26688
rect 81008 26623 81328 26624
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 65648 26144 65968 26145
rect 65648 26080 65656 26144
rect 65720 26080 65736 26144
rect 65800 26080 65816 26144
rect 65880 26080 65896 26144
rect 65960 26080 65968 26144
rect 65648 26079 65968 26080
rect 96368 26144 96688 26145
rect 96368 26080 96376 26144
rect 96440 26080 96456 26144
rect 96520 26080 96536 26144
rect 96600 26080 96616 26144
rect 96680 26080 96688 26144
rect 96368 26079 96688 26080
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 50288 25600 50608 25601
rect 50288 25536 50296 25600
rect 50360 25536 50376 25600
rect 50440 25536 50456 25600
rect 50520 25536 50536 25600
rect 50600 25536 50608 25600
rect 50288 25535 50608 25536
rect 81008 25600 81328 25601
rect 81008 25536 81016 25600
rect 81080 25536 81096 25600
rect 81160 25536 81176 25600
rect 81240 25536 81256 25600
rect 81320 25536 81328 25600
rect 81008 25535 81328 25536
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 65648 25056 65968 25057
rect 65648 24992 65656 25056
rect 65720 24992 65736 25056
rect 65800 24992 65816 25056
rect 65880 24992 65896 25056
rect 65960 24992 65968 25056
rect 65648 24991 65968 24992
rect 96368 25056 96688 25057
rect 96368 24992 96376 25056
rect 96440 24992 96456 25056
rect 96520 24992 96536 25056
rect 96600 24992 96616 25056
rect 96680 24992 96688 25056
rect 96368 24991 96688 24992
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 50288 24512 50608 24513
rect 50288 24448 50296 24512
rect 50360 24448 50376 24512
rect 50440 24448 50456 24512
rect 50520 24448 50536 24512
rect 50600 24448 50608 24512
rect 50288 24447 50608 24448
rect 81008 24512 81328 24513
rect 81008 24448 81016 24512
rect 81080 24448 81096 24512
rect 81160 24448 81176 24512
rect 81240 24448 81256 24512
rect 81320 24448 81328 24512
rect 81008 24447 81328 24448
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 65648 23968 65968 23969
rect 65648 23904 65656 23968
rect 65720 23904 65736 23968
rect 65800 23904 65816 23968
rect 65880 23904 65896 23968
rect 65960 23904 65968 23968
rect 65648 23903 65968 23904
rect 96368 23968 96688 23969
rect 96368 23904 96376 23968
rect 96440 23904 96456 23968
rect 96520 23904 96536 23968
rect 96600 23904 96616 23968
rect 96680 23904 96688 23968
rect 96368 23903 96688 23904
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 50288 23424 50608 23425
rect 50288 23360 50296 23424
rect 50360 23360 50376 23424
rect 50440 23360 50456 23424
rect 50520 23360 50536 23424
rect 50600 23360 50608 23424
rect 50288 23359 50608 23360
rect 81008 23424 81328 23425
rect 81008 23360 81016 23424
rect 81080 23360 81096 23424
rect 81160 23360 81176 23424
rect 81240 23360 81256 23424
rect 81320 23360 81328 23424
rect 81008 23359 81328 23360
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 65648 22880 65968 22881
rect 65648 22816 65656 22880
rect 65720 22816 65736 22880
rect 65800 22816 65816 22880
rect 65880 22816 65896 22880
rect 65960 22816 65968 22880
rect 65648 22815 65968 22816
rect 96368 22880 96688 22881
rect 96368 22816 96376 22880
rect 96440 22816 96456 22880
rect 96520 22816 96536 22880
rect 96600 22816 96616 22880
rect 96680 22816 96688 22880
rect 96368 22815 96688 22816
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 50288 22336 50608 22337
rect 50288 22272 50296 22336
rect 50360 22272 50376 22336
rect 50440 22272 50456 22336
rect 50520 22272 50536 22336
rect 50600 22272 50608 22336
rect 50288 22271 50608 22272
rect 81008 22336 81328 22337
rect 81008 22272 81016 22336
rect 81080 22272 81096 22336
rect 81160 22272 81176 22336
rect 81240 22272 81256 22336
rect 81320 22272 81328 22336
rect 81008 22271 81328 22272
rect 43069 21994 43135 21997
rect 47945 21994 48011 21997
rect 43069 21992 48011 21994
rect 43069 21936 43074 21992
rect 43130 21936 47950 21992
rect 48006 21936 48011 21992
rect 43069 21934 48011 21936
rect 43069 21931 43135 21934
rect 47945 21931 48011 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 65648 21792 65968 21793
rect 65648 21728 65656 21792
rect 65720 21728 65736 21792
rect 65800 21728 65816 21792
rect 65880 21728 65896 21792
rect 65960 21728 65968 21792
rect 65648 21727 65968 21728
rect 96368 21792 96688 21793
rect 96368 21728 96376 21792
rect 96440 21728 96456 21792
rect 96520 21728 96536 21792
rect 96600 21728 96616 21792
rect 96680 21728 96688 21792
rect 96368 21727 96688 21728
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 50288 21248 50608 21249
rect 50288 21184 50296 21248
rect 50360 21184 50376 21248
rect 50440 21184 50456 21248
rect 50520 21184 50536 21248
rect 50600 21184 50608 21248
rect 50288 21183 50608 21184
rect 81008 21248 81328 21249
rect 81008 21184 81016 21248
rect 81080 21184 81096 21248
rect 81160 21184 81176 21248
rect 81240 21184 81256 21248
rect 81320 21184 81328 21248
rect 81008 21183 81328 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 65648 20704 65968 20705
rect 65648 20640 65656 20704
rect 65720 20640 65736 20704
rect 65800 20640 65816 20704
rect 65880 20640 65896 20704
rect 65960 20640 65968 20704
rect 65648 20639 65968 20640
rect 96368 20704 96688 20705
rect 96368 20640 96376 20704
rect 96440 20640 96456 20704
rect 96520 20640 96536 20704
rect 96600 20640 96616 20704
rect 96680 20640 96688 20704
rect 96368 20639 96688 20640
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 50288 20160 50608 20161
rect 50288 20096 50296 20160
rect 50360 20096 50376 20160
rect 50440 20096 50456 20160
rect 50520 20096 50536 20160
rect 50600 20096 50608 20160
rect 50288 20095 50608 20096
rect 81008 20160 81328 20161
rect 81008 20096 81016 20160
rect 81080 20096 81096 20160
rect 81160 20096 81176 20160
rect 81240 20096 81256 20160
rect 81320 20096 81328 20160
rect 81008 20095 81328 20096
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 65648 19616 65968 19617
rect 65648 19552 65656 19616
rect 65720 19552 65736 19616
rect 65800 19552 65816 19616
rect 65880 19552 65896 19616
rect 65960 19552 65968 19616
rect 65648 19551 65968 19552
rect 96368 19616 96688 19617
rect 96368 19552 96376 19616
rect 96440 19552 96456 19616
rect 96520 19552 96536 19616
rect 96600 19552 96616 19616
rect 96680 19552 96688 19616
rect 96368 19551 96688 19552
rect 44449 19546 44515 19549
rect 45093 19546 45159 19549
rect 44449 19544 45159 19546
rect 44449 19488 44454 19544
rect 44510 19488 45098 19544
rect 45154 19488 45159 19544
rect 44449 19486 45159 19488
rect 44449 19483 44515 19486
rect 45093 19483 45159 19486
rect 44541 19410 44607 19413
rect 45369 19410 45435 19413
rect 44541 19408 45435 19410
rect 44541 19352 44546 19408
rect 44602 19352 45374 19408
rect 45430 19352 45435 19408
rect 44541 19350 45435 19352
rect 44541 19347 44607 19350
rect 45369 19347 45435 19350
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 50288 19072 50608 19073
rect 50288 19008 50296 19072
rect 50360 19008 50376 19072
rect 50440 19008 50456 19072
rect 50520 19008 50536 19072
rect 50600 19008 50608 19072
rect 50288 19007 50608 19008
rect 81008 19072 81328 19073
rect 81008 19008 81016 19072
rect 81080 19008 81096 19072
rect 81160 19008 81176 19072
rect 81240 19008 81256 19072
rect 81320 19008 81328 19072
rect 81008 19007 81328 19008
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 65648 18528 65968 18529
rect 65648 18464 65656 18528
rect 65720 18464 65736 18528
rect 65800 18464 65816 18528
rect 65880 18464 65896 18528
rect 65960 18464 65968 18528
rect 65648 18463 65968 18464
rect 96368 18528 96688 18529
rect 96368 18464 96376 18528
rect 96440 18464 96456 18528
rect 96520 18464 96536 18528
rect 96600 18464 96616 18528
rect 96680 18464 96688 18528
rect 96368 18463 96688 18464
rect 67725 18322 67791 18325
rect 71129 18322 71195 18325
rect 67725 18320 71195 18322
rect 67725 18264 67730 18320
rect 67786 18264 71134 18320
rect 71190 18264 71195 18320
rect 67725 18262 71195 18264
rect 67725 18259 67791 18262
rect 71129 18259 71195 18262
rect 70485 18186 70551 18189
rect 71313 18186 71379 18189
rect 70485 18184 71379 18186
rect 70485 18128 70490 18184
rect 70546 18128 71318 18184
rect 71374 18128 71379 18184
rect 70485 18126 71379 18128
rect 70485 18123 70551 18126
rect 71313 18123 71379 18126
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 50288 17984 50608 17985
rect 50288 17920 50296 17984
rect 50360 17920 50376 17984
rect 50440 17920 50456 17984
rect 50520 17920 50536 17984
rect 50600 17920 50608 17984
rect 50288 17919 50608 17920
rect 81008 17984 81328 17985
rect 81008 17920 81016 17984
rect 81080 17920 81096 17984
rect 81160 17920 81176 17984
rect 81240 17920 81256 17984
rect 81320 17920 81328 17984
rect 81008 17919 81328 17920
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 65648 17440 65968 17441
rect 65648 17376 65656 17440
rect 65720 17376 65736 17440
rect 65800 17376 65816 17440
rect 65880 17376 65896 17440
rect 65960 17376 65968 17440
rect 65648 17375 65968 17376
rect 96368 17440 96688 17441
rect 96368 17376 96376 17440
rect 96440 17376 96456 17440
rect 96520 17376 96536 17440
rect 96600 17376 96616 17440
rect 96680 17376 96688 17440
rect 96368 17375 96688 17376
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 50288 16896 50608 16897
rect 50288 16832 50296 16896
rect 50360 16832 50376 16896
rect 50440 16832 50456 16896
rect 50520 16832 50536 16896
rect 50600 16832 50608 16896
rect 50288 16831 50608 16832
rect 81008 16896 81328 16897
rect 81008 16832 81016 16896
rect 81080 16832 81096 16896
rect 81160 16832 81176 16896
rect 81240 16832 81256 16896
rect 81320 16832 81328 16896
rect 81008 16831 81328 16832
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 65648 16352 65968 16353
rect 65648 16288 65656 16352
rect 65720 16288 65736 16352
rect 65800 16288 65816 16352
rect 65880 16288 65896 16352
rect 65960 16288 65968 16352
rect 65648 16287 65968 16288
rect 96368 16352 96688 16353
rect 96368 16288 96376 16352
rect 96440 16288 96456 16352
rect 96520 16288 96536 16352
rect 96600 16288 96616 16352
rect 96680 16288 96688 16352
rect 96368 16287 96688 16288
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 50288 15808 50608 15809
rect 50288 15744 50296 15808
rect 50360 15744 50376 15808
rect 50440 15744 50456 15808
rect 50520 15744 50536 15808
rect 50600 15744 50608 15808
rect 50288 15743 50608 15744
rect 81008 15808 81328 15809
rect 81008 15744 81016 15808
rect 81080 15744 81096 15808
rect 81160 15744 81176 15808
rect 81240 15744 81256 15808
rect 81320 15744 81328 15808
rect 81008 15743 81328 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 65648 15264 65968 15265
rect 65648 15200 65656 15264
rect 65720 15200 65736 15264
rect 65800 15200 65816 15264
rect 65880 15200 65896 15264
rect 65960 15200 65968 15264
rect 65648 15199 65968 15200
rect 96368 15264 96688 15265
rect 96368 15200 96376 15264
rect 96440 15200 96456 15264
rect 96520 15200 96536 15264
rect 96600 15200 96616 15264
rect 96680 15200 96688 15264
rect 96368 15199 96688 15200
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 50288 14720 50608 14721
rect 50288 14656 50296 14720
rect 50360 14656 50376 14720
rect 50440 14656 50456 14720
rect 50520 14656 50536 14720
rect 50600 14656 50608 14720
rect 50288 14655 50608 14656
rect 81008 14720 81328 14721
rect 81008 14656 81016 14720
rect 81080 14656 81096 14720
rect 81160 14656 81176 14720
rect 81240 14656 81256 14720
rect 81320 14656 81328 14720
rect 81008 14655 81328 14656
rect 44541 14378 44607 14381
rect 45369 14378 45435 14381
rect 44541 14376 45435 14378
rect 44541 14320 44546 14376
rect 44602 14320 45374 14376
rect 45430 14320 45435 14376
rect 44541 14318 45435 14320
rect 44541 14315 44607 14318
rect 45369 14315 45435 14318
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 65648 14176 65968 14177
rect 65648 14112 65656 14176
rect 65720 14112 65736 14176
rect 65800 14112 65816 14176
rect 65880 14112 65896 14176
rect 65960 14112 65968 14176
rect 65648 14111 65968 14112
rect 96368 14176 96688 14177
rect 96368 14112 96376 14176
rect 96440 14112 96456 14176
rect 96520 14112 96536 14176
rect 96600 14112 96616 14176
rect 96680 14112 96688 14176
rect 96368 14111 96688 14112
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 50288 13632 50608 13633
rect 50288 13568 50296 13632
rect 50360 13568 50376 13632
rect 50440 13568 50456 13632
rect 50520 13568 50536 13632
rect 50600 13568 50608 13632
rect 50288 13567 50608 13568
rect 81008 13632 81328 13633
rect 81008 13568 81016 13632
rect 81080 13568 81096 13632
rect 81160 13568 81176 13632
rect 81240 13568 81256 13632
rect 81320 13568 81328 13632
rect 81008 13567 81328 13568
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 65648 13088 65968 13089
rect 65648 13024 65656 13088
rect 65720 13024 65736 13088
rect 65800 13024 65816 13088
rect 65880 13024 65896 13088
rect 65960 13024 65968 13088
rect 65648 13023 65968 13024
rect 96368 13088 96688 13089
rect 96368 13024 96376 13088
rect 96440 13024 96456 13088
rect 96520 13024 96536 13088
rect 96600 13024 96616 13088
rect 96680 13024 96688 13088
rect 96368 13023 96688 13024
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 50288 12544 50608 12545
rect 50288 12480 50296 12544
rect 50360 12480 50376 12544
rect 50440 12480 50456 12544
rect 50520 12480 50536 12544
rect 50600 12480 50608 12544
rect 50288 12479 50608 12480
rect 81008 12544 81328 12545
rect 81008 12480 81016 12544
rect 81080 12480 81096 12544
rect 81160 12480 81176 12544
rect 81240 12480 81256 12544
rect 81320 12480 81328 12544
rect 81008 12479 81328 12480
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 65648 12000 65968 12001
rect 65648 11936 65656 12000
rect 65720 11936 65736 12000
rect 65800 11936 65816 12000
rect 65880 11936 65896 12000
rect 65960 11936 65968 12000
rect 65648 11935 65968 11936
rect 96368 12000 96688 12001
rect 96368 11936 96376 12000
rect 96440 11936 96456 12000
rect 96520 11936 96536 12000
rect 96600 11936 96616 12000
rect 96680 11936 96688 12000
rect 96368 11935 96688 11936
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 50288 11456 50608 11457
rect 50288 11392 50296 11456
rect 50360 11392 50376 11456
rect 50440 11392 50456 11456
rect 50520 11392 50536 11456
rect 50600 11392 50608 11456
rect 50288 11391 50608 11392
rect 81008 11456 81328 11457
rect 81008 11392 81016 11456
rect 81080 11392 81096 11456
rect 81160 11392 81176 11456
rect 81240 11392 81256 11456
rect 81320 11392 81328 11456
rect 81008 11391 81328 11392
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 65648 10912 65968 10913
rect 65648 10848 65656 10912
rect 65720 10848 65736 10912
rect 65800 10848 65816 10912
rect 65880 10848 65896 10912
rect 65960 10848 65968 10912
rect 65648 10847 65968 10848
rect 96368 10912 96688 10913
rect 96368 10848 96376 10912
rect 96440 10848 96456 10912
rect 96520 10848 96536 10912
rect 96600 10848 96616 10912
rect 96680 10848 96688 10912
rect 96368 10847 96688 10848
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 50288 10368 50608 10369
rect 50288 10304 50296 10368
rect 50360 10304 50376 10368
rect 50440 10304 50456 10368
rect 50520 10304 50536 10368
rect 50600 10304 50608 10368
rect 50288 10303 50608 10304
rect 81008 10368 81328 10369
rect 81008 10304 81016 10368
rect 81080 10304 81096 10368
rect 81160 10304 81176 10368
rect 81240 10304 81256 10368
rect 81320 10304 81328 10368
rect 81008 10303 81328 10304
rect 62941 10026 63007 10029
rect 63861 10026 63927 10029
rect 62941 10024 63927 10026
rect 62941 9968 62946 10024
rect 63002 9968 63866 10024
rect 63922 9968 63927 10024
rect 62941 9966 63927 9968
rect 62941 9963 63007 9966
rect 63861 9963 63927 9966
rect 62757 9890 62823 9893
rect 63585 9890 63651 9893
rect 62757 9888 63651 9890
rect 62757 9832 62762 9888
rect 62818 9832 63590 9888
rect 63646 9832 63651 9888
rect 62757 9830 63651 9832
rect 62757 9827 62823 9830
rect 63585 9827 63651 9830
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 65648 9824 65968 9825
rect 65648 9760 65656 9824
rect 65720 9760 65736 9824
rect 65800 9760 65816 9824
rect 65880 9760 65896 9824
rect 65960 9760 65968 9824
rect 65648 9759 65968 9760
rect 96368 9824 96688 9825
rect 96368 9760 96376 9824
rect 96440 9760 96456 9824
rect 96520 9760 96536 9824
rect 96600 9760 96616 9824
rect 96680 9760 96688 9824
rect 96368 9759 96688 9760
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 50288 9280 50608 9281
rect 50288 9216 50296 9280
rect 50360 9216 50376 9280
rect 50440 9216 50456 9280
rect 50520 9216 50536 9280
rect 50600 9216 50608 9280
rect 50288 9215 50608 9216
rect 81008 9280 81328 9281
rect 81008 9216 81016 9280
rect 81080 9216 81096 9280
rect 81160 9216 81176 9280
rect 81240 9216 81256 9280
rect 81320 9216 81328 9280
rect 81008 9215 81328 9216
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 65648 8736 65968 8737
rect 65648 8672 65656 8736
rect 65720 8672 65736 8736
rect 65800 8672 65816 8736
rect 65880 8672 65896 8736
rect 65960 8672 65968 8736
rect 65648 8671 65968 8672
rect 96368 8736 96688 8737
rect 96368 8672 96376 8736
rect 96440 8672 96456 8736
rect 96520 8672 96536 8736
rect 96600 8672 96616 8736
rect 96680 8672 96688 8736
rect 96368 8671 96688 8672
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 50288 8192 50608 8193
rect 50288 8128 50296 8192
rect 50360 8128 50376 8192
rect 50440 8128 50456 8192
rect 50520 8128 50536 8192
rect 50600 8128 50608 8192
rect 50288 8127 50608 8128
rect 81008 8192 81328 8193
rect 81008 8128 81016 8192
rect 81080 8128 81096 8192
rect 81160 8128 81176 8192
rect 81240 8128 81256 8192
rect 81320 8128 81328 8192
rect 81008 8127 81328 8128
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 65648 7648 65968 7649
rect 65648 7584 65656 7648
rect 65720 7584 65736 7648
rect 65800 7584 65816 7648
rect 65880 7584 65896 7648
rect 65960 7584 65968 7648
rect 65648 7583 65968 7584
rect 96368 7648 96688 7649
rect 96368 7584 96376 7648
rect 96440 7584 96456 7648
rect 96520 7584 96536 7648
rect 96600 7584 96616 7648
rect 96680 7584 96688 7648
rect 96368 7583 96688 7584
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 50288 7104 50608 7105
rect 50288 7040 50296 7104
rect 50360 7040 50376 7104
rect 50440 7040 50456 7104
rect 50520 7040 50536 7104
rect 50600 7040 50608 7104
rect 50288 7039 50608 7040
rect 81008 7104 81328 7105
rect 81008 7040 81016 7104
rect 81080 7040 81096 7104
rect 81160 7040 81176 7104
rect 81240 7040 81256 7104
rect 81320 7040 81328 7104
rect 81008 7039 81328 7040
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 65648 6560 65968 6561
rect 65648 6496 65656 6560
rect 65720 6496 65736 6560
rect 65800 6496 65816 6560
rect 65880 6496 65896 6560
rect 65960 6496 65968 6560
rect 65648 6495 65968 6496
rect 96368 6560 96688 6561
rect 96368 6496 96376 6560
rect 96440 6496 96456 6560
rect 96520 6496 96536 6560
rect 96600 6496 96616 6560
rect 96680 6496 96688 6560
rect 96368 6495 96688 6496
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 50288 6016 50608 6017
rect 50288 5952 50296 6016
rect 50360 5952 50376 6016
rect 50440 5952 50456 6016
rect 50520 5952 50536 6016
rect 50600 5952 50608 6016
rect 50288 5951 50608 5952
rect 81008 6016 81328 6017
rect 81008 5952 81016 6016
rect 81080 5952 81096 6016
rect 81160 5952 81176 6016
rect 81240 5952 81256 6016
rect 81320 5952 81328 6016
rect 81008 5951 81328 5952
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 65648 5472 65968 5473
rect 65648 5408 65656 5472
rect 65720 5408 65736 5472
rect 65800 5408 65816 5472
rect 65880 5408 65896 5472
rect 65960 5408 65968 5472
rect 65648 5407 65968 5408
rect 96368 5472 96688 5473
rect 96368 5408 96376 5472
rect 96440 5408 96456 5472
rect 96520 5408 96536 5472
rect 96600 5408 96616 5472
rect 96680 5408 96688 5472
rect 96368 5407 96688 5408
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 50288 4928 50608 4929
rect 50288 4864 50296 4928
rect 50360 4864 50376 4928
rect 50440 4864 50456 4928
rect 50520 4864 50536 4928
rect 50600 4864 50608 4928
rect 50288 4863 50608 4864
rect 81008 4928 81328 4929
rect 81008 4864 81016 4928
rect 81080 4864 81096 4928
rect 81160 4864 81176 4928
rect 81240 4864 81256 4928
rect 81320 4864 81328 4928
rect 81008 4863 81328 4864
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 65648 4384 65968 4385
rect 65648 4320 65656 4384
rect 65720 4320 65736 4384
rect 65800 4320 65816 4384
rect 65880 4320 65896 4384
rect 65960 4320 65968 4384
rect 65648 4319 65968 4320
rect 96368 4384 96688 4385
rect 96368 4320 96376 4384
rect 96440 4320 96456 4384
rect 96520 4320 96536 4384
rect 96600 4320 96616 4384
rect 96680 4320 96688 4384
rect 96368 4319 96688 4320
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 50288 3840 50608 3841
rect 50288 3776 50296 3840
rect 50360 3776 50376 3840
rect 50440 3776 50456 3840
rect 50520 3776 50536 3840
rect 50600 3776 50608 3840
rect 50288 3775 50608 3776
rect 81008 3840 81328 3841
rect 81008 3776 81016 3840
rect 81080 3776 81096 3840
rect 81160 3776 81176 3840
rect 81240 3776 81256 3840
rect 81320 3776 81328 3840
rect 81008 3775 81328 3776
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 65648 3296 65968 3297
rect 65648 3232 65656 3296
rect 65720 3232 65736 3296
rect 65800 3232 65816 3296
rect 65880 3232 65896 3296
rect 65960 3232 65968 3296
rect 65648 3231 65968 3232
rect 96368 3296 96688 3297
rect 96368 3232 96376 3296
rect 96440 3232 96456 3296
rect 96520 3232 96536 3296
rect 96600 3232 96616 3296
rect 96680 3232 96688 3296
rect 96368 3231 96688 3232
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 50288 2752 50608 2753
rect 50288 2688 50296 2752
rect 50360 2688 50376 2752
rect 50440 2688 50456 2752
rect 50520 2688 50536 2752
rect 50600 2688 50608 2752
rect 50288 2687 50608 2688
rect 81008 2752 81328 2753
rect 81008 2688 81016 2752
rect 81080 2688 81096 2752
rect 81160 2688 81176 2752
rect 81240 2688 81256 2752
rect 81320 2688 81328 2752
rect 81008 2687 81328 2688
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 65648 2208 65968 2209
rect 65648 2144 65656 2208
rect 65720 2144 65736 2208
rect 65800 2144 65816 2208
rect 65880 2144 65896 2208
rect 65960 2144 65968 2208
rect 65648 2143 65968 2144
rect 96368 2208 96688 2209
rect 96368 2144 96376 2208
rect 96440 2144 96456 2208
rect 96520 2144 96536 2208
rect 96600 2144 96616 2208
rect 96680 2144 96688 2208
rect 96368 2143 96688 2144
<< via3 >>
rect 19576 97404 19640 97408
rect 19576 97348 19580 97404
rect 19580 97348 19636 97404
rect 19636 97348 19640 97404
rect 19576 97344 19640 97348
rect 19656 97404 19720 97408
rect 19656 97348 19660 97404
rect 19660 97348 19716 97404
rect 19716 97348 19720 97404
rect 19656 97344 19720 97348
rect 19736 97404 19800 97408
rect 19736 97348 19740 97404
rect 19740 97348 19796 97404
rect 19796 97348 19800 97404
rect 19736 97344 19800 97348
rect 19816 97404 19880 97408
rect 19816 97348 19820 97404
rect 19820 97348 19876 97404
rect 19876 97348 19880 97404
rect 19816 97344 19880 97348
rect 50296 97404 50360 97408
rect 50296 97348 50300 97404
rect 50300 97348 50356 97404
rect 50356 97348 50360 97404
rect 50296 97344 50360 97348
rect 50376 97404 50440 97408
rect 50376 97348 50380 97404
rect 50380 97348 50436 97404
rect 50436 97348 50440 97404
rect 50376 97344 50440 97348
rect 50456 97404 50520 97408
rect 50456 97348 50460 97404
rect 50460 97348 50516 97404
rect 50516 97348 50520 97404
rect 50456 97344 50520 97348
rect 50536 97404 50600 97408
rect 50536 97348 50540 97404
rect 50540 97348 50596 97404
rect 50596 97348 50600 97404
rect 50536 97344 50600 97348
rect 81016 97404 81080 97408
rect 81016 97348 81020 97404
rect 81020 97348 81076 97404
rect 81076 97348 81080 97404
rect 81016 97344 81080 97348
rect 81096 97404 81160 97408
rect 81096 97348 81100 97404
rect 81100 97348 81156 97404
rect 81156 97348 81160 97404
rect 81096 97344 81160 97348
rect 81176 97404 81240 97408
rect 81176 97348 81180 97404
rect 81180 97348 81236 97404
rect 81236 97348 81240 97404
rect 81176 97344 81240 97348
rect 81256 97404 81320 97408
rect 81256 97348 81260 97404
rect 81260 97348 81316 97404
rect 81316 97348 81320 97404
rect 81256 97344 81320 97348
rect 4216 96860 4280 96864
rect 4216 96804 4220 96860
rect 4220 96804 4276 96860
rect 4276 96804 4280 96860
rect 4216 96800 4280 96804
rect 4296 96860 4360 96864
rect 4296 96804 4300 96860
rect 4300 96804 4356 96860
rect 4356 96804 4360 96860
rect 4296 96800 4360 96804
rect 4376 96860 4440 96864
rect 4376 96804 4380 96860
rect 4380 96804 4436 96860
rect 4436 96804 4440 96860
rect 4376 96800 4440 96804
rect 4456 96860 4520 96864
rect 4456 96804 4460 96860
rect 4460 96804 4516 96860
rect 4516 96804 4520 96860
rect 4456 96800 4520 96804
rect 34936 96860 35000 96864
rect 34936 96804 34940 96860
rect 34940 96804 34996 96860
rect 34996 96804 35000 96860
rect 34936 96800 35000 96804
rect 35016 96860 35080 96864
rect 35016 96804 35020 96860
rect 35020 96804 35076 96860
rect 35076 96804 35080 96860
rect 35016 96800 35080 96804
rect 35096 96860 35160 96864
rect 35096 96804 35100 96860
rect 35100 96804 35156 96860
rect 35156 96804 35160 96860
rect 35096 96800 35160 96804
rect 35176 96860 35240 96864
rect 35176 96804 35180 96860
rect 35180 96804 35236 96860
rect 35236 96804 35240 96860
rect 35176 96800 35240 96804
rect 65656 96860 65720 96864
rect 65656 96804 65660 96860
rect 65660 96804 65716 96860
rect 65716 96804 65720 96860
rect 65656 96800 65720 96804
rect 65736 96860 65800 96864
rect 65736 96804 65740 96860
rect 65740 96804 65796 96860
rect 65796 96804 65800 96860
rect 65736 96800 65800 96804
rect 65816 96860 65880 96864
rect 65816 96804 65820 96860
rect 65820 96804 65876 96860
rect 65876 96804 65880 96860
rect 65816 96800 65880 96804
rect 65896 96860 65960 96864
rect 65896 96804 65900 96860
rect 65900 96804 65956 96860
rect 65956 96804 65960 96860
rect 65896 96800 65960 96804
rect 96376 96860 96440 96864
rect 96376 96804 96380 96860
rect 96380 96804 96436 96860
rect 96436 96804 96440 96860
rect 96376 96800 96440 96804
rect 96456 96860 96520 96864
rect 96456 96804 96460 96860
rect 96460 96804 96516 96860
rect 96516 96804 96520 96860
rect 96456 96800 96520 96804
rect 96536 96860 96600 96864
rect 96536 96804 96540 96860
rect 96540 96804 96596 96860
rect 96596 96804 96600 96860
rect 96536 96800 96600 96804
rect 96616 96860 96680 96864
rect 96616 96804 96620 96860
rect 96620 96804 96676 96860
rect 96676 96804 96680 96860
rect 96616 96800 96680 96804
rect 19576 96316 19640 96320
rect 19576 96260 19580 96316
rect 19580 96260 19636 96316
rect 19636 96260 19640 96316
rect 19576 96256 19640 96260
rect 19656 96316 19720 96320
rect 19656 96260 19660 96316
rect 19660 96260 19716 96316
rect 19716 96260 19720 96316
rect 19656 96256 19720 96260
rect 19736 96316 19800 96320
rect 19736 96260 19740 96316
rect 19740 96260 19796 96316
rect 19796 96260 19800 96316
rect 19736 96256 19800 96260
rect 19816 96316 19880 96320
rect 19816 96260 19820 96316
rect 19820 96260 19876 96316
rect 19876 96260 19880 96316
rect 19816 96256 19880 96260
rect 50296 96316 50360 96320
rect 50296 96260 50300 96316
rect 50300 96260 50356 96316
rect 50356 96260 50360 96316
rect 50296 96256 50360 96260
rect 50376 96316 50440 96320
rect 50376 96260 50380 96316
rect 50380 96260 50436 96316
rect 50436 96260 50440 96316
rect 50376 96256 50440 96260
rect 50456 96316 50520 96320
rect 50456 96260 50460 96316
rect 50460 96260 50516 96316
rect 50516 96260 50520 96316
rect 50456 96256 50520 96260
rect 50536 96316 50600 96320
rect 50536 96260 50540 96316
rect 50540 96260 50596 96316
rect 50596 96260 50600 96316
rect 50536 96256 50600 96260
rect 81016 96316 81080 96320
rect 81016 96260 81020 96316
rect 81020 96260 81076 96316
rect 81076 96260 81080 96316
rect 81016 96256 81080 96260
rect 81096 96316 81160 96320
rect 81096 96260 81100 96316
rect 81100 96260 81156 96316
rect 81156 96260 81160 96316
rect 81096 96256 81160 96260
rect 81176 96316 81240 96320
rect 81176 96260 81180 96316
rect 81180 96260 81236 96316
rect 81236 96260 81240 96316
rect 81176 96256 81240 96260
rect 81256 96316 81320 96320
rect 81256 96260 81260 96316
rect 81260 96260 81316 96316
rect 81316 96260 81320 96316
rect 81256 96256 81320 96260
rect 4216 95772 4280 95776
rect 4216 95716 4220 95772
rect 4220 95716 4276 95772
rect 4276 95716 4280 95772
rect 4216 95712 4280 95716
rect 4296 95772 4360 95776
rect 4296 95716 4300 95772
rect 4300 95716 4356 95772
rect 4356 95716 4360 95772
rect 4296 95712 4360 95716
rect 4376 95772 4440 95776
rect 4376 95716 4380 95772
rect 4380 95716 4436 95772
rect 4436 95716 4440 95772
rect 4376 95712 4440 95716
rect 4456 95772 4520 95776
rect 4456 95716 4460 95772
rect 4460 95716 4516 95772
rect 4516 95716 4520 95772
rect 4456 95712 4520 95716
rect 34936 95772 35000 95776
rect 34936 95716 34940 95772
rect 34940 95716 34996 95772
rect 34996 95716 35000 95772
rect 34936 95712 35000 95716
rect 35016 95772 35080 95776
rect 35016 95716 35020 95772
rect 35020 95716 35076 95772
rect 35076 95716 35080 95772
rect 35016 95712 35080 95716
rect 35096 95772 35160 95776
rect 35096 95716 35100 95772
rect 35100 95716 35156 95772
rect 35156 95716 35160 95772
rect 35096 95712 35160 95716
rect 35176 95772 35240 95776
rect 35176 95716 35180 95772
rect 35180 95716 35236 95772
rect 35236 95716 35240 95772
rect 35176 95712 35240 95716
rect 65656 95772 65720 95776
rect 65656 95716 65660 95772
rect 65660 95716 65716 95772
rect 65716 95716 65720 95772
rect 65656 95712 65720 95716
rect 65736 95772 65800 95776
rect 65736 95716 65740 95772
rect 65740 95716 65796 95772
rect 65796 95716 65800 95772
rect 65736 95712 65800 95716
rect 65816 95772 65880 95776
rect 65816 95716 65820 95772
rect 65820 95716 65876 95772
rect 65876 95716 65880 95772
rect 65816 95712 65880 95716
rect 65896 95772 65960 95776
rect 65896 95716 65900 95772
rect 65900 95716 65956 95772
rect 65956 95716 65960 95772
rect 65896 95712 65960 95716
rect 96376 95772 96440 95776
rect 96376 95716 96380 95772
rect 96380 95716 96436 95772
rect 96436 95716 96440 95772
rect 96376 95712 96440 95716
rect 96456 95772 96520 95776
rect 96456 95716 96460 95772
rect 96460 95716 96516 95772
rect 96516 95716 96520 95772
rect 96456 95712 96520 95716
rect 96536 95772 96600 95776
rect 96536 95716 96540 95772
rect 96540 95716 96596 95772
rect 96596 95716 96600 95772
rect 96536 95712 96600 95716
rect 96616 95772 96680 95776
rect 96616 95716 96620 95772
rect 96620 95716 96676 95772
rect 96676 95716 96680 95772
rect 96616 95712 96680 95716
rect 19576 95228 19640 95232
rect 19576 95172 19580 95228
rect 19580 95172 19636 95228
rect 19636 95172 19640 95228
rect 19576 95168 19640 95172
rect 19656 95228 19720 95232
rect 19656 95172 19660 95228
rect 19660 95172 19716 95228
rect 19716 95172 19720 95228
rect 19656 95168 19720 95172
rect 19736 95228 19800 95232
rect 19736 95172 19740 95228
rect 19740 95172 19796 95228
rect 19796 95172 19800 95228
rect 19736 95168 19800 95172
rect 19816 95228 19880 95232
rect 19816 95172 19820 95228
rect 19820 95172 19876 95228
rect 19876 95172 19880 95228
rect 19816 95168 19880 95172
rect 50296 95228 50360 95232
rect 50296 95172 50300 95228
rect 50300 95172 50356 95228
rect 50356 95172 50360 95228
rect 50296 95168 50360 95172
rect 50376 95228 50440 95232
rect 50376 95172 50380 95228
rect 50380 95172 50436 95228
rect 50436 95172 50440 95228
rect 50376 95168 50440 95172
rect 50456 95228 50520 95232
rect 50456 95172 50460 95228
rect 50460 95172 50516 95228
rect 50516 95172 50520 95228
rect 50456 95168 50520 95172
rect 50536 95228 50600 95232
rect 50536 95172 50540 95228
rect 50540 95172 50596 95228
rect 50596 95172 50600 95228
rect 50536 95168 50600 95172
rect 81016 95228 81080 95232
rect 81016 95172 81020 95228
rect 81020 95172 81076 95228
rect 81076 95172 81080 95228
rect 81016 95168 81080 95172
rect 81096 95228 81160 95232
rect 81096 95172 81100 95228
rect 81100 95172 81156 95228
rect 81156 95172 81160 95228
rect 81096 95168 81160 95172
rect 81176 95228 81240 95232
rect 81176 95172 81180 95228
rect 81180 95172 81236 95228
rect 81236 95172 81240 95228
rect 81176 95168 81240 95172
rect 81256 95228 81320 95232
rect 81256 95172 81260 95228
rect 81260 95172 81316 95228
rect 81316 95172 81320 95228
rect 81256 95168 81320 95172
rect 4216 94684 4280 94688
rect 4216 94628 4220 94684
rect 4220 94628 4276 94684
rect 4276 94628 4280 94684
rect 4216 94624 4280 94628
rect 4296 94684 4360 94688
rect 4296 94628 4300 94684
rect 4300 94628 4356 94684
rect 4356 94628 4360 94684
rect 4296 94624 4360 94628
rect 4376 94684 4440 94688
rect 4376 94628 4380 94684
rect 4380 94628 4436 94684
rect 4436 94628 4440 94684
rect 4376 94624 4440 94628
rect 4456 94684 4520 94688
rect 4456 94628 4460 94684
rect 4460 94628 4516 94684
rect 4516 94628 4520 94684
rect 4456 94624 4520 94628
rect 34936 94684 35000 94688
rect 34936 94628 34940 94684
rect 34940 94628 34996 94684
rect 34996 94628 35000 94684
rect 34936 94624 35000 94628
rect 35016 94684 35080 94688
rect 35016 94628 35020 94684
rect 35020 94628 35076 94684
rect 35076 94628 35080 94684
rect 35016 94624 35080 94628
rect 35096 94684 35160 94688
rect 35096 94628 35100 94684
rect 35100 94628 35156 94684
rect 35156 94628 35160 94684
rect 35096 94624 35160 94628
rect 35176 94684 35240 94688
rect 35176 94628 35180 94684
rect 35180 94628 35236 94684
rect 35236 94628 35240 94684
rect 35176 94624 35240 94628
rect 65656 94684 65720 94688
rect 65656 94628 65660 94684
rect 65660 94628 65716 94684
rect 65716 94628 65720 94684
rect 65656 94624 65720 94628
rect 65736 94684 65800 94688
rect 65736 94628 65740 94684
rect 65740 94628 65796 94684
rect 65796 94628 65800 94684
rect 65736 94624 65800 94628
rect 65816 94684 65880 94688
rect 65816 94628 65820 94684
rect 65820 94628 65876 94684
rect 65876 94628 65880 94684
rect 65816 94624 65880 94628
rect 65896 94684 65960 94688
rect 65896 94628 65900 94684
rect 65900 94628 65956 94684
rect 65956 94628 65960 94684
rect 65896 94624 65960 94628
rect 96376 94684 96440 94688
rect 96376 94628 96380 94684
rect 96380 94628 96436 94684
rect 96436 94628 96440 94684
rect 96376 94624 96440 94628
rect 96456 94684 96520 94688
rect 96456 94628 96460 94684
rect 96460 94628 96516 94684
rect 96516 94628 96520 94684
rect 96456 94624 96520 94628
rect 96536 94684 96600 94688
rect 96536 94628 96540 94684
rect 96540 94628 96596 94684
rect 96596 94628 96600 94684
rect 96536 94624 96600 94628
rect 96616 94684 96680 94688
rect 96616 94628 96620 94684
rect 96620 94628 96676 94684
rect 96676 94628 96680 94684
rect 96616 94624 96680 94628
rect 19576 94140 19640 94144
rect 19576 94084 19580 94140
rect 19580 94084 19636 94140
rect 19636 94084 19640 94140
rect 19576 94080 19640 94084
rect 19656 94140 19720 94144
rect 19656 94084 19660 94140
rect 19660 94084 19716 94140
rect 19716 94084 19720 94140
rect 19656 94080 19720 94084
rect 19736 94140 19800 94144
rect 19736 94084 19740 94140
rect 19740 94084 19796 94140
rect 19796 94084 19800 94140
rect 19736 94080 19800 94084
rect 19816 94140 19880 94144
rect 19816 94084 19820 94140
rect 19820 94084 19876 94140
rect 19876 94084 19880 94140
rect 19816 94080 19880 94084
rect 50296 94140 50360 94144
rect 50296 94084 50300 94140
rect 50300 94084 50356 94140
rect 50356 94084 50360 94140
rect 50296 94080 50360 94084
rect 50376 94140 50440 94144
rect 50376 94084 50380 94140
rect 50380 94084 50436 94140
rect 50436 94084 50440 94140
rect 50376 94080 50440 94084
rect 50456 94140 50520 94144
rect 50456 94084 50460 94140
rect 50460 94084 50516 94140
rect 50516 94084 50520 94140
rect 50456 94080 50520 94084
rect 50536 94140 50600 94144
rect 50536 94084 50540 94140
rect 50540 94084 50596 94140
rect 50596 94084 50600 94140
rect 50536 94080 50600 94084
rect 81016 94140 81080 94144
rect 81016 94084 81020 94140
rect 81020 94084 81076 94140
rect 81076 94084 81080 94140
rect 81016 94080 81080 94084
rect 81096 94140 81160 94144
rect 81096 94084 81100 94140
rect 81100 94084 81156 94140
rect 81156 94084 81160 94140
rect 81096 94080 81160 94084
rect 81176 94140 81240 94144
rect 81176 94084 81180 94140
rect 81180 94084 81236 94140
rect 81236 94084 81240 94140
rect 81176 94080 81240 94084
rect 81256 94140 81320 94144
rect 81256 94084 81260 94140
rect 81260 94084 81316 94140
rect 81316 94084 81320 94140
rect 81256 94080 81320 94084
rect 4216 93596 4280 93600
rect 4216 93540 4220 93596
rect 4220 93540 4276 93596
rect 4276 93540 4280 93596
rect 4216 93536 4280 93540
rect 4296 93596 4360 93600
rect 4296 93540 4300 93596
rect 4300 93540 4356 93596
rect 4356 93540 4360 93596
rect 4296 93536 4360 93540
rect 4376 93596 4440 93600
rect 4376 93540 4380 93596
rect 4380 93540 4436 93596
rect 4436 93540 4440 93596
rect 4376 93536 4440 93540
rect 4456 93596 4520 93600
rect 4456 93540 4460 93596
rect 4460 93540 4516 93596
rect 4516 93540 4520 93596
rect 4456 93536 4520 93540
rect 34936 93596 35000 93600
rect 34936 93540 34940 93596
rect 34940 93540 34996 93596
rect 34996 93540 35000 93596
rect 34936 93536 35000 93540
rect 35016 93596 35080 93600
rect 35016 93540 35020 93596
rect 35020 93540 35076 93596
rect 35076 93540 35080 93596
rect 35016 93536 35080 93540
rect 35096 93596 35160 93600
rect 35096 93540 35100 93596
rect 35100 93540 35156 93596
rect 35156 93540 35160 93596
rect 35096 93536 35160 93540
rect 35176 93596 35240 93600
rect 35176 93540 35180 93596
rect 35180 93540 35236 93596
rect 35236 93540 35240 93596
rect 35176 93536 35240 93540
rect 65656 93596 65720 93600
rect 65656 93540 65660 93596
rect 65660 93540 65716 93596
rect 65716 93540 65720 93596
rect 65656 93536 65720 93540
rect 65736 93596 65800 93600
rect 65736 93540 65740 93596
rect 65740 93540 65796 93596
rect 65796 93540 65800 93596
rect 65736 93536 65800 93540
rect 65816 93596 65880 93600
rect 65816 93540 65820 93596
rect 65820 93540 65876 93596
rect 65876 93540 65880 93596
rect 65816 93536 65880 93540
rect 65896 93596 65960 93600
rect 65896 93540 65900 93596
rect 65900 93540 65956 93596
rect 65956 93540 65960 93596
rect 65896 93536 65960 93540
rect 96376 93596 96440 93600
rect 96376 93540 96380 93596
rect 96380 93540 96436 93596
rect 96436 93540 96440 93596
rect 96376 93536 96440 93540
rect 96456 93596 96520 93600
rect 96456 93540 96460 93596
rect 96460 93540 96516 93596
rect 96516 93540 96520 93596
rect 96456 93536 96520 93540
rect 96536 93596 96600 93600
rect 96536 93540 96540 93596
rect 96540 93540 96596 93596
rect 96596 93540 96600 93596
rect 96536 93536 96600 93540
rect 96616 93596 96680 93600
rect 96616 93540 96620 93596
rect 96620 93540 96676 93596
rect 96676 93540 96680 93596
rect 96616 93536 96680 93540
rect 19576 93052 19640 93056
rect 19576 92996 19580 93052
rect 19580 92996 19636 93052
rect 19636 92996 19640 93052
rect 19576 92992 19640 92996
rect 19656 93052 19720 93056
rect 19656 92996 19660 93052
rect 19660 92996 19716 93052
rect 19716 92996 19720 93052
rect 19656 92992 19720 92996
rect 19736 93052 19800 93056
rect 19736 92996 19740 93052
rect 19740 92996 19796 93052
rect 19796 92996 19800 93052
rect 19736 92992 19800 92996
rect 19816 93052 19880 93056
rect 19816 92996 19820 93052
rect 19820 92996 19876 93052
rect 19876 92996 19880 93052
rect 19816 92992 19880 92996
rect 50296 93052 50360 93056
rect 50296 92996 50300 93052
rect 50300 92996 50356 93052
rect 50356 92996 50360 93052
rect 50296 92992 50360 92996
rect 50376 93052 50440 93056
rect 50376 92996 50380 93052
rect 50380 92996 50436 93052
rect 50436 92996 50440 93052
rect 50376 92992 50440 92996
rect 50456 93052 50520 93056
rect 50456 92996 50460 93052
rect 50460 92996 50516 93052
rect 50516 92996 50520 93052
rect 50456 92992 50520 92996
rect 50536 93052 50600 93056
rect 50536 92996 50540 93052
rect 50540 92996 50596 93052
rect 50596 92996 50600 93052
rect 50536 92992 50600 92996
rect 81016 93052 81080 93056
rect 81016 92996 81020 93052
rect 81020 92996 81076 93052
rect 81076 92996 81080 93052
rect 81016 92992 81080 92996
rect 81096 93052 81160 93056
rect 81096 92996 81100 93052
rect 81100 92996 81156 93052
rect 81156 92996 81160 93052
rect 81096 92992 81160 92996
rect 81176 93052 81240 93056
rect 81176 92996 81180 93052
rect 81180 92996 81236 93052
rect 81236 92996 81240 93052
rect 81176 92992 81240 92996
rect 81256 93052 81320 93056
rect 81256 92996 81260 93052
rect 81260 92996 81316 93052
rect 81316 92996 81320 93052
rect 81256 92992 81320 92996
rect 4216 92508 4280 92512
rect 4216 92452 4220 92508
rect 4220 92452 4276 92508
rect 4276 92452 4280 92508
rect 4216 92448 4280 92452
rect 4296 92508 4360 92512
rect 4296 92452 4300 92508
rect 4300 92452 4356 92508
rect 4356 92452 4360 92508
rect 4296 92448 4360 92452
rect 4376 92508 4440 92512
rect 4376 92452 4380 92508
rect 4380 92452 4436 92508
rect 4436 92452 4440 92508
rect 4376 92448 4440 92452
rect 4456 92508 4520 92512
rect 4456 92452 4460 92508
rect 4460 92452 4516 92508
rect 4516 92452 4520 92508
rect 4456 92448 4520 92452
rect 34936 92508 35000 92512
rect 34936 92452 34940 92508
rect 34940 92452 34996 92508
rect 34996 92452 35000 92508
rect 34936 92448 35000 92452
rect 35016 92508 35080 92512
rect 35016 92452 35020 92508
rect 35020 92452 35076 92508
rect 35076 92452 35080 92508
rect 35016 92448 35080 92452
rect 35096 92508 35160 92512
rect 35096 92452 35100 92508
rect 35100 92452 35156 92508
rect 35156 92452 35160 92508
rect 35096 92448 35160 92452
rect 35176 92508 35240 92512
rect 35176 92452 35180 92508
rect 35180 92452 35236 92508
rect 35236 92452 35240 92508
rect 35176 92448 35240 92452
rect 65656 92508 65720 92512
rect 65656 92452 65660 92508
rect 65660 92452 65716 92508
rect 65716 92452 65720 92508
rect 65656 92448 65720 92452
rect 65736 92508 65800 92512
rect 65736 92452 65740 92508
rect 65740 92452 65796 92508
rect 65796 92452 65800 92508
rect 65736 92448 65800 92452
rect 65816 92508 65880 92512
rect 65816 92452 65820 92508
rect 65820 92452 65876 92508
rect 65876 92452 65880 92508
rect 65816 92448 65880 92452
rect 65896 92508 65960 92512
rect 65896 92452 65900 92508
rect 65900 92452 65956 92508
rect 65956 92452 65960 92508
rect 65896 92448 65960 92452
rect 96376 92508 96440 92512
rect 96376 92452 96380 92508
rect 96380 92452 96436 92508
rect 96436 92452 96440 92508
rect 96376 92448 96440 92452
rect 96456 92508 96520 92512
rect 96456 92452 96460 92508
rect 96460 92452 96516 92508
rect 96516 92452 96520 92508
rect 96456 92448 96520 92452
rect 96536 92508 96600 92512
rect 96536 92452 96540 92508
rect 96540 92452 96596 92508
rect 96596 92452 96600 92508
rect 96536 92448 96600 92452
rect 96616 92508 96680 92512
rect 96616 92452 96620 92508
rect 96620 92452 96676 92508
rect 96676 92452 96680 92508
rect 96616 92448 96680 92452
rect 19576 91964 19640 91968
rect 19576 91908 19580 91964
rect 19580 91908 19636 91964
rect 19636 91908 19640 91964
rect 19576 91904 19640 91908
rect 19656 91964 19720 91968
rect 19656 91908 19660 91964
rect 19660 91908 19716 91964
rect 19716 91908 19720 91964
rect 19656 91904 19720 91908
rect 19736 91964 19800 91968
rect 19736 91908 19740 91964
rect 19740 91908 19796 91964
rect 19796 91908 19800 91964
rect 19736 91904 19800 91908
rect 19816 91964 19880 91968
rect 19816 91908 19820 91964
rect 19820 91908 19876 91964
rect 19876 91908 19880 91964
rect 19816 91904 19880 91908
rect 50296 91964 50360 91968
rect 50296 91908 50300 91964
rect 50300 91908 50356 91964
rect 50356 91908 50360 91964
rect 50296 91904 50360 91908
rect 50376 91964 50440 91968
rect 50376 91908 50380 91964
rect 50380 91908 50436 91964
rect 50436 91908 50440 91964
rect 50376 91904 50440 91908
rect 50456 91964 50520 91968
rect 50456 91908 50460 91964
rect 50460 91908 50516 91964
rect 50516 91908 50520 91964
rect 50456 91904 50520 91908
rect 50536 91964 50600 91968
rect 50536 91908 50540 91964
rect 50540 91908 50596 91964
rect 50596 91908 50600 91964
rect 50536 91904 50600 91908
rect 81016 91964 81080 91968
rect 81016 91908 81020 91964
rect 81020 91908 81076 91964
rect 81076 91908 81080 91964
rect 81016 91904 81080 91908
rect 81096 91964 81160 91968
rect 81096 91908 81100 91964
rect 81100 91908 81156 91964
rect 81156 91908 81160 91964
rect 81096 91904 81160 91908
rect 81176 91964 81240 91968
rect 81176 91908 81180 91964
rect 81180 91908 81236 91964
rect 81236 91908 81240 91964
rect 81176 91904 81240 91908
rect 81256 91964 81320 91968
rect 81256 91908 81260 91964
rect 81260 91908 81316 91964
rect 81316 91908 81320 91964
rect 81256 91904 81320 91908
rect 4216 91420 4280 91424
rect 4216 91364 4220 91420
rect 4220 91364 4276 91420
rect 4276 91364 4280 91420
rect 4216 91360 4280 91364
rect 4296 91420 4360 91424
rect 4296 91364 4300 91420
rect 4300 91364 4356 91420
rect 4356 91364 4360 91420
rect 4296 91360 4360 91364
rect 4376 91420 4440 91424
rect 4376 91364 4380 91420
rect 4380 91364 4436 91420
rect 4436 91364 4440 91420
rect 4376 91360 4440 91364
rect 4456 91420 4520 91424
rect 4456 91364 4460 91420
rect 4460 91364 4516 91420
rect 4516 91364 4520 91420
rect 4456 91360 4520 91364
rect 34936 91420 35000 91424
rect 34936 91364 34940 91420
rect 34940 91364 34996 91420
rect 34996 91364 35000 91420
rect 34936 91360 35000 91364
rect 35016 91420 35080 91424
rect 35016 91364 35020 91420
rect 35020 91364 35076 91420
rect 35076 91364 35080 91420
rect 35016 91360 35080 91364
rect 35096 91420 35160 91424
rect 35096 91364 35100 91420
rect 35100 91364 35156 91420
rect 35156 91364 35160 91420
rect 35096 91360 35160 91364
rect 35176 91420 35240 91424
rect 35176 91364 35180 91420
rect 35180 91364 35236 91420
rect 35236 91364 35240 91420
rect 35176 91360 35240 91364
rect 65656 91420 65720 91424
rect 65656 91364 65660 91420
rect 65660 91364 65716 91420
rect 65716 91364 65720 91420
rect 65656 91360 65720 91364
rect 65736 91420 65800 91424
rect 65736 91364 65740 91420
rect 65740 91364 65796 91420
rect 65796 91364 65800 91420
rect 65736 91360 65800 91364
rect 65816 91420 65880 91424
rect 65816 91364 65820 91420
rect 65820 91364 65876 91420
rect 65876 91364 65880 91420
rect 65816 91360 65880 91364
rect 65896 91420 65960 91424
rect 65896 91364 65900 91420
rect 65900 91364 65956 91420
rect 65956 91364 65960 91420
rect 65896 91360 65960 91364
rect 96376 91420 96440 91424
rect 96376 91364 96380 91420
rect 96380 91364 96436 91420
rect 96436 91364 96440 91420
rect 96376 91360 96440 91364
rect 96456 91420 96520 91424
rect 96456 91364 96460 91420
rect 96460 91364 96516 91420
rect 96516 91364 96520 91420
rect 96456 91360 96520 91364
rect 96536 91420 96600 91424
rect 96536 91364 96540 91420
rect 96540 91364 96596 91420
rect 96596 91364 96600 91420
rect 96536 91360 96600 91364
rect 96616 91420 96680 91424
rect 96616 91364 96620 91420
rect 96620 91364 96676 91420
rect 96676 91364 96680 91420
rect 96616 91360 96680 91364
rect 19576 90876 19640 90880
rect 19576 90820 19580 90876
rect 19580 90820 19636 90876
rect 19636 90820 19640 90876
rect 19576 90816 19640 90820
rect 19656 90876 19720 90880
rect 19656 90820 19660 90876
rect 19660 90820 19716 90876
rect 19716 90820 19720 90876
rect 19656 90816 19720 90820
rect 19736 90876 19800 90880
rect 19736 90820 19740 90876
rect 19740 90820 19796 90876
rect 19796 90820 19800 90876
rect 19736 90816 19800 90820
rect 19816 90876 19880 90880
rect 19816 90820 19820 90876
rect 19820 90820 19876 90876
rect 19876 90820 19880 90876
rect 19816 90816 19880 90820
rect 50296 90876 50360 90880
rect 50296 90820 50300 90876
rect 50300 90820 50356 90876
rect 50356 90820 50360 90876
rect 50296 90816 50360 90820
rect 50376 90876 50440 90880
rect 50376 90820 50380 90876
rect 50380 90820 50436 90876
rect 50436 90820 50440 90876
rect 50376 90816 50440 90820
rect 50456 90876 50520 90880
rect 50456 90820 50460 90876
rect 50460 90820 50516 90876
rect 50516 90820 50520 90876
rect 50456 90816 50520 90820
rect 50536 90876 50600 90880
rect 50536 90820 50540 90876
rect 50540 90820 50596 90876
rect 50596 90820 50600 90876
rect 50536 90816 50600 90820
rect 81016 90876 81080 90880
rect 81016 90820 81020 90876
rect 81020 90820 81076 90876
rect 81076 90820 81080 90876
rect 81016 90816 81080 90820
rect 81096 90876 81160 90880
rect 81096 90820 81100 90876
rect 81100 90820 81156 90876
rect 81156 90820 81160 90876
rect 81096 90816 81160 90820
rect 81176 90876 81240 90880
rect 81176 90820 81180 90876
rect 81180 90820 81236 90876
rect 81236 90820 81240 90876
rect 81176 90816 81240 90820
rect 81256 90876 81320 90880
rect 81256 90820 81260 90876
rect 81260 90820 81316 90876
rect 81316 90820 81320 90876
rect 81256 90816 81320 90820
rect 4216 90332 4280 90336
rect 4216 90276 4220 90332
rect 4220 90276 4276 90332
rect 4276 90276 4280 90332
rect 4216 90272 4280 90276
rect 4296 90332 4360 90336
rect 4296 90276 4300 90332
rect 4300 90276 4356 90332
rect 4356 90276 4360 90332
rect 4296 90272 4360 90276
rect 4376 90332 4440 90336
rect 4376 90276 4380 90332
rect 4380 90276 4436 90332
rect 4436 90276 4440 90332
rect 4376 90272 4440 90276
rect 4456 90332 4520 90336
rect 4456 90276 4460 90332
rect 4460 90276 4516 90332
rect 4516 90276 4520 90332
rect 4456 90272 4520 90276
rect 34936 90332 35000 90336
rect 34936 90276 34940 90332
rect 34940 90276 34996 90332
rect 34996 90276 35000 90332
rect 34936 90272 35000 90276
rect 35016 90332 35080 90336
rect 35016 90276 35020 90332
rect 35020 90276 35076 90332
rect 35076 90276 35080 90332
rect 35016 90272 35080 90276
rect 35096 90332 35160 90336
rect 35096 90276 35100 90332
rect 35100 90276 35156 90332
rect 35156 90276 35160 90332
rect 35096 90272 35160 90276
rect 35176 90332 35240 90336
rect 35176 90276 35180 90332
rect 35180 90276 35236 90332
rect 35236 90276 35240 90332
rect 35176 90272 35240 90276
rect 65656 90332 65720 90336
rect 65656 90276 65660 90332
rect 65660 90276 65716 90332
rect 65716 90276 65720 90332
rect 65656 90272 65720 90276
rect 65736 90332 65800 90336
rect 65736 90276 65740 90332
rect 65740 90276 65796 90332
rect 65796 90276 65800 90332
rect 65736 90272 65800 90276
rect 65816 90332 65880 90336
rect 65816 90276 65820 90332
rect 65820 90276 65876 90332
rect 65876 90276 65880 90332
rect 65816 90272 65880 90276
rect 65896 90332 65960 90336
rect 65896 90276 65900 90332
rect 65900 90276 65956 90332
rect 65956 90276 65960 90332
rect 65896 90272 65960 90276
rect 96376 90332 96440 90336
rect 96376 90276 96380 90332
rect 96380 90276 96436 90332
rect 96436 90276 96440 90332
rect 96376 90272 96440 90276
rect 96456 90332 96520 90336
rect 96456 90276 96460 90332
rect 96460 90276 96516 90332
rect 96516 90276 96520 90332
rect 96456 90272 96520 90276
rect 96536 90332 96600 90336
rect 96536 90276 96540 90332
rect 96540 90276 96596 90332
rect 96596 90276 96600 90332
rect 96536 90272 96600 90276
rect 96616 90332 96680 90336
rect 96616 90276 96620 90332
rect 96620 90276 96676 90332
rect 96676 90276 96680 90332
rect 96616 90272 96680 90276
rect 19576 89788 19640 89792
rect 19576 89732 19580 89788
rect 19580 89732 19636 89788
rect 19636 89732 19640 89788
rect 19576 89728 19640 89732
rect 19656 89788 19720 89792
rect 19656 89732 19660 89788
rect 19660 89732 19716 89788
rect 19716 89732 19720 89788
rect 19656 89728 19720 89732
rect 19736 89788 19800 89792
rect 19736 89732 19740 89788
rect 19740 89732 19796 89788
rect 19796 89732 19800 89788
rect 19736 89728 19800 89732
rect 19816 89788 19880 89792
rect 19816 89732 19820 89788
rect 19820 89732 19876 89788
rect 19876 89732 19880 89788
rect 19816 89728 19880 89732
rect 50296 89788 50360 89792
rect 50296 89732 50300 89788
rect 50300 89732 50356 89788
rect 50356 89732 50360 89788
rect 50296 89728 50360 89732
rect 50376 89788 50440 89792
rect 50376 89732 50380 89788
rect 50380 89732 50436 89788
rect 50436 89732 50440 89788
rect 50376 89728 50440 89732
rect 50456 89788 50520 89792
rect 50456 89732 50460 89788
rect 50460 89732 50516 89788
rect 50516 89732 50520 89788
rect 50456 89728 50520 89732
rect 50536 89788 50600 89792
rect 50536 89732 50540 89788
rect 50540 89732 50596 89788
rect 50596 89732 50600 89788
rect 50536 89728 50600 89732
rect 81016 89788 81080 89792
rect 81016 89732 81020 89788
rect 81020 89732 81076 89788
rect 81076 89732 81080 89788
rect 81016 89728 81080 89732
rect 81096 89788 81160 89792
rect 81096 89732 81100 89788
rect 81100 89732 81156 89788
rect 81156 89732 81160 89788
rect 81096 89728 81160 89732
rect 81176 89788 81240 89792
rect 81176 89732 81180 89788
rect 81180 89732 81236 89788
rect 81236 89732 81240 89788
rect 81176 89728 81240 89732
rect 81256 89788 81320 89792
rect 81256 89732 81260 89788
rect 81260 89732 81316 89788
rect 81316 89732 81320 89788
rect 81256 89728 81320 89732
rect 4216 89244 4280 89248
rect 4216 89188 4220 89244
rect 4220 89188 4276 89244
rect 4276 89188 4280 89244
rect 4216 89184 4280 89188
rect 4296 89244 4360 89248
rect 4296 89188 4300 89244
rect 4300 89188 4356 89244
rect 4356 89188 4360 89244
rect 4296 89184 4360 89188
rect 4376 89244 4440 89248
rect 4376 89188 4380 89244
rect 4380 89188 4436 89244
rect 4436 89188 4440 89244
rect 4376 89184 4440 89188
rect 4456 89244 4520 89248
rect 4456 89188 4460 89244
rect 4460 89188 4516 89244
rect 4516 89188 4520 89244
rect 4456 89184 4520 89188
rect 34936 89244 35000 89248
rect 34936 89188 34940 89244
rect 34940 89188 34996 89244
rect 34996 89188 35000 89244
rect 34936 89184 35000 89188
rect 35016 89244 35080 89248
rect 35016 89188 35020 89244
rect 35020 89188 35076 89244
rect 35076 89188 35080 89244
rect 35016 89184 35080 89188
rect 35096 89244 35160 89248
rect 35096 89188 35100 89244
rect 35100 89188 35156 89244
rect 35156 89188 35160 89244
rect 35096 89184 35160 89188
rect 35176 89244 35240 89248
rect 35176 89188 35180 89244
rect 35180 89188 35236 89244
rect 35236 89188 35240 89244
rect 35176 89184 35240 89188
rect 65656 89244 65720 89248
rect 65656 89188 65660 89244
rect 65660 89188 65716 89244
rect 65716 89188 65720 89244
rect 65656 89184 65720 89188
rect 65736 89244 65800 89248
rect 65736 89188 65740 89244
rect 65740 89188 65796 89244
rect 65796 89188 65800 89244
rect 65736 89184 65800 89188
rect 65816 89244 65880 89248
rect 65816 89188 65820 89244
rect 65820 89188 65876 89244
rect 65876 89188 65880 89244
rect 65816 89184 65880 89188
rect 65896 89244 65960 89248
rect 65896 89188 65900 89244
rect 65900 89188 65956 89244
rect 65956 89188 65960 89244
rect 65896 89184 65960 89188
rect 96376 89244 96440 89248
rect 96376 89188 96380 89244
rect 96380 89188 96436 89244
rect 96436 89188 96440 89244
rect 96376 89184 96440 89188
rect 96456 89244 96520 89248
rect 96456 89188 96460 89244
rect 96460 89188 96516 89244
rect 96516 89188 96520 89244
rect 96456 89184 96520 89188
rect 96536 89244 96600 89248
rect 96536 89188 96540 89244
rect 96540 89188 96596 89244
rect 96596 89188 96600 89244
rect 96536 89184 96600 89188
rect 96616 89244 96680 89248
rect 96616 89188 96620 89244
rect 96620 89188 96676 89244
rect 96676 89188 96680 89244
rect 96616 89184 96680 89188
rect 19576 88700 19640 88704
rect 19576 88644 19580 88700
rect 19580 88644 19636 88700
rect 19636 88644 19640 88700
rect 19576 88640 19640 88644
rect 19656 88700 19720 88704
rect 19656 88644 19660 88700
rect 19660 88644 19716 88700
rect 19716 88644 19720 88700
rect 19656 88640 19720 88644
rect 19736 88700 19800 88704
rect 19736 88644 19740 88700
rect 19740 88644 19796 88700
rect 19796 88644 19800 88700
rect 19736 88640 19800 88644
rect 19816 88700 19880 88704
rect 19816 88644 19820 88700
rect 19820 88644 19876 88700
rect 19876 88644 19880 88700
rect 19816 88640 19880 88644
rect 50296 88700 50360 88704
rect 50296 88644 50300 88700
rect 50300 88644 50356 88700
rect 50356 88644 50360 88700
rect 50296 88640 50360 88644
rect 50376 88700 50440 88704
rect 50376 88644 50380 88700
rect 50380 88644 50436 88700
rect 50436 88644 50440 88700
rect 50376 88640 50440 88644
rect 50456 88700 50520 88704
rect 50456 88644 50460 88700
rect 50460 88644 50516 88700
rect 50516 88644 50520 88700
rect 50456 88640 50520 88644
rect 50536 88700 50600 88704
rect 50536 88644 50540 88700
rect 50540 88644 50596 88700
rect 50596 88644 50600 88700
rect 50536 88640 50600 88644
rect 81016 88700 81080 88704
rect 81016 88644 81020 88700
rect 81020 88644 81076 88700
rect 81076 88644 81080 88700
rect 81016 88640 81080 88644
rect 81096 88700 81160 88704
rect 81096 88644 81100 88700
rect 81100 88644 81156 88700
rect 81156 88644 81160 88700
rect 81096 88640 81160 88644
rect 81176 88700 81240 88704
rect 81176 88644 81180 88700
rect 81180 88644 81236 88700
rect 81236 88644 81240 88700
rect 81176 88640 81240 88644
rect 81256 88700 81320 88704
rect 81256 88644 81260 88700
rect 81260 88644 81316 88700
rect 81316 88644 81320 88700
rect 81256 88640 81320 88644
rect 4216 88156 4280 88160
rect 4216 88100 4220 88156
rect 4220 88100 4276 88156
rect 4276 88100 4280 88156
rect 4216 88096 4280 88100
rect 4296 88156 4360 88160
rect 4296 88100 4300 88156
rect 4300 88100 4356 88156
rect 4356 88100 4360 88156
rect 4296 88096 4360 88100
rect 4376 88156 4440 88160
rect 4376 88100 4380 88156
rect 4380 88100 4436 88156
rect 4436 88100 4440 88156
rect 4376 88096 4440 88100
rect 4456 88156 4520 88160
rect 4456 88100 4460 88156
rect 4460 88100 4516 88156
rect 4516 88100 4520 88156
rect 4456 88096 4520 88100
rect 34936 88156 35000 88160
rect 34936 88100 34940 88156
rect 34940 88100 34996 88156
rect 34996 88100 35000 88156
rect 34936 88096 35000 88100
rect 35016 88156 35080 88160
rect 35016 88100 35020 88156
rect 35020 88100 35076 88156
rect 35076 88100 35080 88156
rect 35016 88096 35080 88100
rect 35096 88156 35160 88160
rect 35096 88100 35100 88156
rect 35100 88100 35156 88156
rect 35156 88100 35160 88156
rect 35096 88096 35160 88100
rect 35176 88156 35240 88160
rect 35176 88100 35180 88156
rect 35180 88100 35236 88156
rect 35236 88100 35240 88156
rect 35176 88096 35240 88100
rect 65656 88156 65720 88160
rect 65656 88100 65660 88156
rect 65660 88100 65716 88156
rect 65716 88100 65720 88156
rect 65656 88096 65720 88100
rect 65736 88156 65800 88160
rect 65736 88100 65740 88156
rect 65740 88100 65796 88156
rect 65796 88100 65800 88156
rect 65736 88096 65800 88100
rect 65816 88156 65880 88160
rect 65816 88100 65820 88156
rect 65820 88100 65876 88156
rect 65876 88100 65880 88156
rect 65816 88096 65880 88100
rect 65896 88156 65960 88160
rect 65896 88100 65900 88156
rect 65900 88100 65956 88156
rect 65956 88100 65960 88156
rect 65896 88096 65960 88100
rect 96376 88156 96440 88160
rect 96376 88100 96380 88156
rect 96380 88100 96436 88156
rect 96436 88100 96440 88156
rect 96376 88096 96440 88100
rect 96456 88156 96520 88160
rect 96456 88100 96460 88156
rect 96460 88100 96516 88156
rect 96516 88100 96520 88156
rect 96456 88096 96520 88100
rect 96536 88156 96600 88160
rect 96536 88100 96540 88156
rect 96540 88100 96596 88156
rect 96596 88100 96600 88156
rect 96536 88096 96600 88100
rect 96616 88156 96680 88160
rect 96616 88100 96620 88156
rect 96620 88100 96676 88156
rect 96676 88100 96680 88156
rect 96616 88096 96680 88100
rect 19576 87612 19640 87616
rect 19576 87556 19580 87612
rect 19580 87556 19636 87612
rect 19636 87556 19640 87612
rect 19576 87552 19640 87556
rect 19656 87612 19720 87616
rect 19656 87556 19660 87612
rect 19660 87556 19716 87612
rect 19716 87556 19720 87612
rect 19656 87552 19720 87556
rect 19736 87612 19800 87616
rect 19736 87556 19740 87612
rect 19740 87556 19796 87612
rect 19796 87556 19800 87612
rect 19736 87552 19800 87556
rect 19816 87612 19880 87616
rect 19816 87556 19820 87612
rect 19820 87556 19876 87612
rect 19876 87556 19880 87612
rect 19816 87552 19880 87556
rect 50296 87612 50360 87616
rect 50296 87556 50300 87612
rect 50300 87556 50356 87612
rect 50356 87556 50360 87612
rect 50296 87552 50360 87556
rect 50376 87612 50440 87616
rect 50376 87556 50380 87612
rect 50380 87556 50436 87612
rect 50436 87556 50440 87612
rect 50376 87552 50440 87556
rect 50456 87612 50520 87616
rect 50456 87556 50460 87612
rect 50460 87556 50516 87612
rect 50516 87556 50520 87612
rect 50456 87552 50520 87556
rect 50536 87612 50600 87616
rect 50536 87556 50540 87612
rect 50540 87556 50596 87612
rect 50596 87556 50600 87612
rect 50536 87552 50600 87556
rect 81016 87612 81080 87616
rect 81016 87556 81020 87612
rect 81020 87556 81076 87612
rect 81076 87556 81080 87612
rect 81016 87552 81080 87556
rect 81096 87612 81160 87616
rect 81096 87556 81100 87612
rect 81100 87556 81156 87612
rect 81156 87556 81160 87612
rect 81096 87552 81160 87556
rect 81176 87612 81240 87616
rect 81176 87556 81180 87612
rect 81180 87556 81236 87612
rect 81236 87556 81240 87612
rect 81176 87552 81240 87556
rect 81256 87612 81320 87616
rect 81256 87556 81260 87612
rect 81260 87556 81316 87612
rect 81316 87556 81320 87612
rect 81256 87552 81320 87556
rect 4216 87068 4280 87072
rect 4216 87012 4220 87068
rect 4220 87012 4276 87068
rect 4276 87012 4280 87068
rect 4216 87008 4280 87012
rect 4296 87068 4360 87072
rect 4296 87012 4300 87068
rect 4300 87012 4356 87068
rect 4356 87012 4360 87068
rect 4296 87008 4360 87012
rect 4376 87068 4440 87072
rect 4376 87012 4380 87068
rect 4380 87012 4436 87068
rect 4436 87012 4440 87068
rect 4376 87008 4440 87012
rect 4456 87068 4520 87072
rect 4456 87012 4460 87068
rect 4460 87012 4516 87068
rect 4516 87012 4520 87068
rect 4456 87008 4520 87012
rect 34936 87068 35000 87072
rect 34936 87012 34940 87068
rect 34940 87012 34996 87068
rect 34996 87012 35000 87068
rect 34936 87008 35000 87012
rect 35016 87068 35080 87072
rect 35016 87012 35020 87068
rect 35020 87012 35076 87068
rect 35076 87012 35080 87068
rect 35016 87008 35080 87012
rect 35096 87068 35160 87072
rect 35096 87012 35100 87068
rect 35100 87012 35156 87068
rect 35156 87012 35160 87068
rect 35096 87008 35160 87012
rect 35176 87068 35240 87072
rect 35176 87012 35180 87068
rect 35180 87012 35236 87068
rect 35236 87012 35240 87068
rect 35176 87008 35240 87012
rect 65656 87068 65720 87072
rect 65656 87012 65660 87068
rect 65660 87012 65716 87068
rect 65716 87012 65720 87068
rect 65656 87008 65720 87012
rect 65736 87068 65800 87072
rect 65736 87012 65740 87068
rect 65740 87012 65796 87068
rect 65796 87012 65800 87068
rect 65736 87008 65800 87012
rect 65816 87068 65880 87072
rect 65816 87012 65820 87068
rect 65820 87012 65876 87068
rect 65876 87012 65880 87068
rect 65816 87008 65880 87012
rect 65896 87068 65960 87072
rect 65896 87012 65900 87068
rect 65900 87012 65956 87068
rect 65956 87012 65960 87068
rect 65896 87008 65960 87012
rect 96376 87068 96440 87072
rect 96376 87012 96380 87068
rect 96380 87012 96436 87068
rect 96436 87012 96440 87068
rect 96376 87008 96440 87012
rect 96456 87068 96520 87072
rect 96456 87012 96460 87068
rect 96460 87012 96516 87068
rect 96516 87012 96520 87068
rect 96456 87008 96520 87012
rect 96536 87068 96600 87072
rect 96536 87012 96540 87068
rect 96540 87012 96596 87068
rect 96596 87012 96600 87068
rect 96536 87008 96600 87012
rect 96616 87068 96680 87072
rect 96616 87012 96620 87068
rect 96620 87012 96676 87068
rect 96676 87012 96680 87068
rect 96616 87008 96680 87012
rect 19576 86524 19640 86528
rect 19576 86468 19580 86524
rect 19580 86468 19636 86524
rect 19636 86468 19640 86524
rect 19576 86464 19640 86468
rect 19656 86524 19720 86528
rect 19656 86468 19660 86524
rect 19660 86468 19716 86524
rect 19716 86468 19720 86524
rect 19656 86464 19720 86468
rect 19736 86524 19800 86528
rect 19736 86468 19740 86524
rect 19740 86468 19796 86524
rect 19796 86468 19800 86524
rect 19736 86464 19800 86468
rect 19816 86524 19880 86528
rect 19816 86468 19820 86524
rect 19820 86468 19876 86524
rect 19876 86468 19880 86524
rect 19816 86464 19880 86468
rect 50296 86524 50360 86528
rect 50296 86468 50300 86524
rect 50300 86468 50356 86524
rect 50356 86468 50360 86524
rect 50296 86464 50360 86468
rect 50376 86524 50440 86528
rect 50376 86468 50380 86524
rect 50380 86468 50436 86524
rect 50436 86468 50440 86524
rect 50376 86464 50440 86468
rect 50456 86524 50520 86528
rect 50456 86468 50460 86524
rect 50460 86468 50516 86524
rect 50516 86468 50520 86524
rect 50456 86464 50520 86468
rect 50536 86524 50600 86528
rect 50536 86468 50540 86524
rect 50540 86468 50596 86524
rect 50596 86468 50600 86524
rect 50536 86464 50600 86468
rect 81016 86524 81080 86528
rect 81016 86468 81020 86524
rect 81020 86468 81076 86524
rect 81076 86468 81080 86524
rect 81016 86464 81080 86468
rect 81096 86524 81160 86528
rect 81096 86468 81100 86524
rect 81100 86468 81156 86524
rect 81156 86468 81160 86524
rect 81096 86464 81160 86468
rect 81176 86524 81240 86528
rect 81176 86468 81180 86524
rect 81180 86468 81236 86524
rect 81236 86468 81240 86524
rect 81176 86464 81240 86468
rect 81256 86524 81320 86528
rect 81256 86468 81260 86524
rect 81260 86468 81316 86524
rect 81316 86468 81320 86524
rect 81256 86464 81320 86468
rect 4216 85980 4280 85984
rect 4216 85924 4220 85980
rect 4220 85924 4276 85980
rect 4276 85924 4280 85980
rect 4216 85920 4280 85924
rect 4296 85980 4360 85984
rect 4296 85924 4300 85980
rect 4300 85924 4356 85980
rect 4356 85924 4360 85980
rect 4296 85920 4360 85924
rect 4376 85980 4440 85984
rect 4376 85924 4380 85980
rect 4380 85924 4436 85980
rect 4436 85924 4440 85980
rect 4376 85920 4440 85924
rect 4456 85980 4520 85984
rect 4456 85924 4460 85980
rect 4460 85924 4516 85980
rect 4516 85924 4520 85980
rect 4456 85920 4520 85924
rect 34936 85980 35000 85984
rect 34936 85924 34940 85980
rect 34940 85924 34996 85980
rect 34996 85924 35000 85980
rect 34936 85920 35000 85924
rect 35016 85980 35080 85984
rect 35016 85924 35020 85980
rect 35020 85924 35076 85980
rect 35076 85924 35080 85980
rect 35016 85920 35080 85924
rect 35096 85980 35160 85984
rect 35096 85924 35100 85980
rect 35100 85924 35156 85980
rect 35156 85924 35160 85980
rect 35096 85920 35160 85924
rect 35176 85980 35240 85984
rect 35176 85924 35180 85980
rect 35180 85924 35236 85980
rect 35236 85924 35240 85980
rect 35176 85920 35240 85924
rect 65656 85980 65720 85984
rect 65656 85924 65660 85980
rect 65660 85924 65716 85980
rect 65716 85924 65720 85980
rect 65656 85920 65720 85924
rect 65736 85980 65800 85984
rect 65736 85924 65740 85980
rect 65740 85924 65796 85980
rect 65796 85924 65800 85980
rect 65736 85920 65800 85924
rect 65816 85980 65880 85984
rect 65816 85924 65820 85980
rect 65820 85924 65876 85980
rect 65876 85924 65880 85980
rect 65816 85920 65880 85924
rect 65896 85980 65960 85984
rect 65896 85924 65900 85980
rect 65900 85924 65956 85980
rect 65956 85924 65960 85980
rect 65896 85920 65960 85924
rect 96376 85980 96440 85984
rect 96376 85924 96380 85980
rect 96380 85924 96436 85980
rect 96436 85924 96440 85980
rect 96376 85920 96440 85924
rect 96456 85980 96520 85984
rect 96456 85924 96460 85980
rect 96460 85924 96516 85980
rect 96516 85924 96520 85980
rect 96456 85920 96520 85924
rect 96536 85980 96600 85984
rect 96536 85924 96540 85980
rect 96540 85924 96596 85980
rect 96596 85924 96600 85980
rect 96536 85920 96600 85924
rect 96616 85980 96680 85984
rect 96616 85924 96620 85980
rect 96620 85924 96676 85980
rect 96676 85924 96680 85980
rect 96616 85920 96680 85924
rect 19576 85436 19640 85440
rect 19576 85380 19580 85436
rect 19580 85380 19636 85436
rect 19636 85380 19640 85436
rect 19576 85376 19640 85380
rect 19656 85436 19720 85440
rect 19656 85380 19660 85436
rect 19660 85380 19716 85436
rect 19716 85380 19720 85436
rect 19656 85376 19720 85380
rect 19736 85436 19800 85440
rect 19736 85380 19740 85436
rect 19740 85380 19796 85436
rect 19796 85380 19800 85436
rect 19736 85376 19800 85380
rect 19816 85436 19880 85440
rect 19816 85380 19820 85436
rect 19820 85380 19876 85436
rect 19876 85380 19880 85436
rect 19816 85376 19880 85380
rect 50296 85436 50360 85440
rect 50296 85380 50300 85436
rect 50300 85380 50356 85436
rect 50356 85380 50360 85436
rect 50296 85376 50360 85380
rect 50376 85436 50440 85440
rect 50376 85380 50380 85436
rect 50380 85380 50436 85436
rect 50436 85380 50440 85436
rect 50376 85376 50440 85380
rect 50456 85436 50520 85440
rect 50456 85380 50460 85436
rect 50460 85380 50516 85436
rect 50516 85380 50520 85436
rect 50456 85376 50520 85380
rect 50536 85436 50600 85440
rect 50536 85380 50540 85436
rect 50540 85380 50596 85436
rect 50596 85380 50600 85436
rect 50536 85376 50600 85380
rect 81016 85436 81080 85440
rect 81016 85380 81020 85436
rect 81020 85380 81076 85436
rect 81076 85380 81080 85436
rect 81016 85376 81080 85380
rect 81096 85436 81160 85440
rect 81096 85380 81100 85436
rect 81100 85380 81156 85436
rect 81156 85380 81160 85436
rect 81096 85376 81160 85380
rect 81176 85436 81240 85440
rect 81176 85380 81180 85436
rect 81180 85380 81236 85436
rect 81236 85380 81240 85436
rect 81176 85376 81240 85380
rect 81256 85436 81320 85440
rect 81256 85380 81260 85436
rect 81260 85380 81316 85436
rect 81316 85380 81320 85436
rect 81256 85376 81320 85380
rect 4216 84892 4280 84896
rect 4216 84836 4220 84892
rect 4220 84836 4276 84892
rect 4276 84836 4280 84892
rect 4216 84832 4280 84836
rect 4296 84892 4360 84896
rect 4296 84836 4300 84892
rect 4300 84836 4356 84892
rect 4356 84836 4360 84892
rect 4296 84832 4360 84836
rect 4376 84892 4440 84896
rect 4376 84836 4380 84892
rect 4380 84836 4436 84892
rect 4436 84836 4440 84892
rect 4376 84832 4440 84836
rect 4456 84892 4520 84896
rect 4456 84836 4460 84892
rect 4460 84836 4516 84892
rect 4516 84836 4520 84892
rect 4456 84832 4520 84836
rect 34936 84892 35000 84896
rect 34936 84836 34940 84892
rect 34940 84836 34996 84892
rect 34996 84836 35000 84892
rect 34936 84832 35000 84836
rect 35016 84892 35080 84896
rect 35016 84836 35020 84892
rect 35020 84836 35076 84892
rect 35076 84836 35080 84892
rect 35016 84832 35080 84836
rect 35096 84892 35160 84896
rect 35096 84836 35100 84892
rect 35100 84836 35156 84892
rect 35156 84836 35160 84892
rect 35096 84832 35160 84836
rect 35176 84892 35240 84896
rect 35176 84836 35180 84892
rect 35180 84836 35236 84892
rect 35236 84836 35240 84892
rect 35176 84832 35240 84836
rect 65656 84892 65720 84896
rect 65656 84836 65660 84892
rect 65660 84836 65716 84892
rect 65716 84836 65720 84892
rect 65656 84832 65720 84836
rect 65736 84892 65800 84896
rect 65736 84836 65740 84892
rect 65740 84836 65796 84892
rect 65796 84836 65800 84892
rect 65736 84832 65800 84836
rect 65816 84892 65880 84896
rect 65816 84836 65820 84892
rect 65820 84836 65876 84892
rect 65876 84836 65880 84892
rect 65816 84832 65880 84836
rect 65896 84892 65960 84896
rect 65896 84836 65900 84892
rect 65900 84836 65956 84892
rect 65956 84836 65960 84892
rect 65896 84832 65960 84836
rect 96376 84892 96440 84896
rect 96376 84836 96380 84892
rect 96380 84836 96436 84892
rect 96436 84836 96440 84892
rect 96376 84832 96440 84836
rect 96456 84892 96520 84896
rect 96456 84836 96460 84892
rect 96460 84836 96516 84892
rect 96516 84836 96520 84892
rect 96456 84832 96520 84836
rect 96536 84892 96600 84896
rect 96536 84836 96540 84892
rect 96540 84836 96596 84892
rect 96596 84836 96600 84892
rect 96536 84832 96600 84836
rect 96616 84892 96680 84896
rect 96616 84836 96620 84892
rect 96620 84836 96676 84892
rect 96676 84836 96680 84892
rect 96616 84832 96680 84836
rect 19576 84348 19640 84352
rect 19576 84292 19580 84348
rect 19580 84292 19636 84348
rect 19636 84292 19640 84348
rect 19576 84288 19640 84292
rect 19656 84348 19720 84352
rect 19656 84292 19660 84348
rect 19660 84292 19716 84348
rect 19716 84292 19720 84348
rect 19656 84288 19720 84292
rect 19736 84348 19800 84352
rect 19736 84292 19740 84348
rect 19740 84292 19796 84348
rect 19796 84292 19800 84348
rect 19736 84288 19800 84292
rect 19816 84348 19880 84352
rect 19816 84292 19820 84348
rect 19820 84292 19876 84348
rect 19876 84292 19880 84348
rect 19816 84288 19880 84292
rect 50296 84348 50360 84352
rect 50296 84292 50300 84348
rect 50300 84292 50356 84348
rect 50356 84292 50360 84348
rect 50296 84288 50360 84292
rect 50376 84348 50440 84352
rect 50376 84292 50380 84348
rect 50380 84292 50436 84348
rect 50436 84292 50440 84348
rect 50376 84288 50440 84292
rect 50456 84348 50520 84352
rect 50456 84292 50460 84348
rect 50460 84292 50516 84348
rect 50516 84292 50520 84348
rect 50456 84288 50520 84292
rect 50536 84348 50600 84352
rect 50536 84292 50540 84348
rect 50540 84292 50596 84348
rect 50596 84292 50600 84348
rect 50536 84288 50600 84292
rect 81016 84348 81080 84352
rect 81016 84292 81020 84348
rect 81020 84292 81076 84348
rect 81076 84292 81080 84348
rect 81016 84288 81080 84292
rect 81096 84348 81160 84352
rect 81096 84292 81100 84348
rect 81100 84292 81156 84348
rect 81156 84292 81160 84348
rect 81096 84288 81160 84292
rect 81176 84348 81240 84352
rect 81176 84292 81180 84348
rect 81180 84292 81236 84348
rect 81236 84292 81240 84348
rect 81176 84288 81240 84292
rect 81256 84348 81320 84352
rect 81256 84292 81260 84348
rect 81260 84292 81316 84348
rect 81316 84292 81320 84348
rect 81256 84288 81320 84292
rect 4216 83804 4280 83808
rect 4216 83748 4220 83804
rect 4220 83748 4276 83804
rect 4276 83748 4280 83804
rect 4216 83744 4280 83748
rect 4296 83804 4360 83808
rect 4296 83748 4300 83804
rect 4300 83748 4356 83804
rect 4356 83748 4360 83804
rect 4296 83744 4360 83748
rect 4376 83804 4440 83808
rect 4376 83748 4380 83804
rect 4380 83748 4436 83804
rect 4436 83748 4440 83804
rect 4376 83744 4440 83748
rect 4456 83804 4520 83808
rect 4456 83748 4460 83804
rect 4460 83748 4516 83804
rect 4516 83748 4520 83804
rect 4456 83744 4520 83748
rect 34936 83804 35000 83808
rect 34936 83748 34940 83804
rect 34940 83748 34996 83804
rect 34996 83748 35000 83804
rect 34936 83744 35000 83748
rect 35016 83804 35080 83808
rect 35016 83748 35020 83804
rect 35020 83748 35076 83804
rect 35076 83748 35080 83804
rect 35016 83744 35080 83748
rect 35096 83804 35160 83808
rect 35096 83748 35100 83804
rect 35100 83748 35156 83804
rect 35156 83748 35160 83804
rect 35096 83744 35160 83748
rect 35176 83804 35240 83808
rect 35176 83748 35180 83804
rect 35180 83748 35236 83804
rect 35236 83748 35240 83804
rect 35176 83744 35240 83748
rect 65656 83804 65720 83808
rect 65656 83748 65660 83804
rect 65660 83748 65716 83804
rect 65716 83748 65720 83804
rect 65656 83744 65720 83748
rect 65736 83804 65800 83808
rect 65736 83748 65740 83804
rect 65740 83748 65796 83804
rect 65796 83748 65800 83804
rect 65736 83744 65800 83748
rect 65816 83804 65880 83808
rect 65816 83748 65820 83804
rect 65820 83748 65876 83804
rect 65876 83748 65880 83804
rect 65816 83744 65880 83748
rect 65896 83804 65960 83808
rect 65896 83748 65900 83804
rect 65900 83748 65956 83804
rect 65956 83748 65960 83804
rect 65896 83744 65960 83748
rect 96376 83804 96440 83808
rect 96376 83748 96380 83804
rect 96380 83748 96436 83804
rect 96436 83748 96440 83804
rect 96376 83744 96440 83748
rect 96456 83804 96520 83808
rect 96456 83748 96460 83804
rect 96460 83748 96516 83804
rect 96516 83748 96520 83804
rect 96456 83744 96520 83748
rect 96536 83804 96600 83808
rect 96536 83748 96540 83804
rect 96540 83748 96596 83804
rect 96596 83748 96600 83804
rect 96536 83744 96600 83748
rect 96616 83804 96680 83808
rect 96616 83748 96620 83804
rect 96620 83748 96676 83804
rect 96676 83748 96680 83804
rect 96616 83744 96680 83748
rect 19576 83260 19640 83264
rect 19576 83204 19580 83260
rect 19580 83204 19636 83260
rect 19636 83204 19640 83260
rect 19576 83200 19640 83204
rect 19656 83260 19720 83264
rect 19656 83204 19660 83260
rect 19660 83204 19716 83260
rect 19716 83204 19720 83260
rect 19656 83200 19720 83204
rect 19736 83260 19800 83264
rect 19736 83204 19740 83260
rect 19740 83204 19796 83260
rect 19796 83204 19800 83260
rect 19736 83200 19800 83204
rect 19816 83260 19880 83264
rect 19816 83204 19820 83260
rect 19820 83204 19876 83260
rect 19876 83204 19880 83260
rect 19816 83200 19880 83204
rect 50296 83260 50360 83264
rect 50296 83204 50300 83260
rect 50300 83204 50356 83260
rect 50356 83204 50360 83260
rect 50296 83200 50360 83204
rect 50376 83260 50440 83264
rect 50376 83204 50380 83260
rect 50380 83204 50436 83260
rect 50436 83204 50440 83260
rect 50376 83200 50440 83204
rect 50456 83260 50520 83264
rect 50456 83204 50460 83260
rect 50460 83204 50516 83260
rect 50516 83204 50520 83260
rect 50456 83200 50520 83204
rect 50536 83260 50600 83264
rect 50536 83204 50540 83260
rect 50540 83204 50596 83260
rect 50596 83204 50600 83260
rect 50536 83200 50600 83204
rect 81016 83260 81080 83264
rect 81016 83204 81020 83260
rect 81020 83204 81076 83260
rect 81076 83204 81080 83260
rect 81016 83200 81080 83204
rect 81096 83260 81160 83264
rect 81096 83204 81100 83260
rect 81100 83204 81156 83260
rect 81156 83204 81160 83260
rect 81096 83200 81160 83204
rect 81176 83260 81240 83264
rect 81176 83204 81180 83260
rect 81180 83204 81236 83260
rect 81236 83204 81240 83260
rect 81176 83200 81240 83204
rect 81256 83260 81320 83264
rect 81256 83204 81260 83260
rect 81260 83204 81316 83260
rect 81316 83204 81320 83260
rect 81256 83200 81320 83204
rect 4216 82716 4280 82720
rect 4216 82660 4220 82716
rect 4220 82660 4276 82716
rect 4276 82660 4280 82716
rect 4216 82656 4280 82660
rect 4296 82716 4360 82720
rect 4296 82660 4300 82716
rect 4300 82660 4356 82716
rect 4356 82660 4360 82716
rect 4296 82656 4360 82660
rect 4376 82716 4440 82720
rect 4376 82660 4380 82716
rect 4380 82660 4436 82716
rect 4436 82660 4440 82716
rect 4376 82656 4440 82660
rect 4456 82716 4520 82720
rect 4456 82660 4460 82716
rect 4460 82660 4516 82716
rect 4516 82660 4520 82716
rect 4456 82656 4520 82660
rect 34936 82716 35000 82720
rect 34936 82660 34940 82716
rect 34940 82660 34996 82716
rect 34996 82660 35000 82716
rect 34936 82656 35000 82660
rect 35016 82716 35080 82720
rect 35016 82660 35020 82716
rect 35020 82660 35076 82716
rect 35076 82660 35080 82716
rect 35016 82656 35080 82660
rect 35096 82716 35160 82720
rect 35096 82660 35100 82716
rect 35100 82660 35156 82716
rect 35156 82660 35160 82716
rect 35096 82656 35160 82660
rect 35176 82716 35240 82720
rect 35176 82660 35180 82716
rect 35180 82660 35236 82716
rect 35236 82660 35240 82716
rect 35176 82656 35240 82660
rect 65656 82716 65720 82720
rect 65656 82660 65660 82716
rect 65660 82660 65716 82716
rect 65716 82660 65720 82716
rect 65656 82656 65720 82660
rect 65736 82716 65800 82720
rect 65736 82660 65740 82716
rect 65740 82660 65796 82716
rect 65796 82660 65800 82716
rect 65736 82656 65800 82660
rect 65816 82716 65880 82720
rect 65816 82660 65820 82716
rect 65820 82660 65876 82716
rect 65876 82660 65880 82716
rect 65816 82656 65880 82660
rect 65896 82716 65960 82720
rect 65896 82660 65900 82716
rect 65900 82660 65956 82716
rect 65956 82660 65960 82716
rect 65896 82656 65960 82660
rect 96376 82716 96440 82720
rect 96376 82660 96380 82716
rect 96380 82660 96436 82716
rect 96436 82660 96440 82716
rect 96376 82656 96440 82660
rect 96456 82716 96520 82720
rect 96456 82660 96460 82716
rect 96460 82660 96516 82716
rect 96516 82660 96520 82716
rect 96456 82656 96520 82660
rect 96536 82716 96600 82720
rect 96536 82660 96540 82716
rect 96540 82660 96596 82716
rect 96596 82660 96600 82716
rect 96536 82656 96600 82660
rect 96616 82716 96680 82720
rect 96616 82660 96620 82716
rect 96620 82660 96676 82716
rect 96676 82660 96680 82716
rect 96616 82656 96680 82660
rect 19576 82172 19640 82176
rect 19576 82116 19580 82172
rect 19580 82116 19636 82172
rect 19636 82116 19640 82172
rect 19576 82112 19640 82116
rect 19656 82172 19720 82176
rect 19656 82116 19660 82172
rect 19660 82116 19716 82172
rect 19716 82116 19720 82172
rect 19656 82112 19720 82116
rect 19736 82172 19800 82176
rect 19736 82116 19740 82172
rect 19740 82116 19796 82172
rect 19796 82116 19800 82172
rect 19736 82112 19800 82116
rect 19816 82172 19880 82176
rect 19816 82116 19820 82172
rect 19820 82116 19876 82172
rect 19876 82116 19880 82172
rect 19816 82112 19880 82116
rect 50296 82172 50360 82176
rect 50296 82116 50300 82172
rect 50300 82116 50356 82172
rect 50356 82116 50360 82172
rect 50296 82112 50360 82116
rect 50376 82172 50440 82176
rect 50376 82116 50380 82172
rect 50380 82116 50436 82172
rect 50436 82116 50440 82172
rect 50376 82112 50440 82116
rect 50456 82172 50520 82176
rect 50456 82116 50460 82172
rect 50460 82116 50516 82172
rect 50516 82116 50520 82172
rect 50456 82112 50520 82116
rect 50536 82172 50600 82176
rect 50536 82116 50540 82172
rect 50540 82116 50596 82172
rect 50596 82116 50600 82172
rect 50536 82112 50600 82116
rect 81016 82172 81080 82176
rect 81016 82116 81020 82172
rect 81020 82116 81076 82172
rect 81076 82116 81080 82172
rect 81016 82112 81080 82116
rect 81096 82172 81160 82176
rect 81096 82116 81100 82172
rect 81100 82116 81156 82172
rect 81156 82116 81160 82172
rect 81096 82112 81160 82116
rect 81176 82172 81240 82176
rect 81176 82116 81180 82172
rect 81180 82116 81236 82172
rect 81236 82116 81240 82172
rect 81176 82112 81240 82116
rect 81256 82172 81320 82176
rect 81256 82116 81260 82172
rect 81260 82116 81316 82172
rect 81316 82116 81320 82172
rect 81256 82112 81320 82116
rect 4216 81628 4280 81632
rect 4216 81572 4220 81628
rect 4220 81572 4276 81628
rect 4276 81572 4280 81628
rect 4216 81568 4280 81572
rect 4296 81628 4360 81632
rect 4296 81572 4300 81628
rect 4300 81572 4356 81628
rect 4356 81572 4360 81628
rect 4296 81568 4360 81572
rect 4376 81628 4440 81632
rect 4376 81572 4380 81628
rect 4380 81572 4436 81628
rect 4436 81572 4440 81628
rect 4376 81568 4440 81572
rect 4456 81628 4520 81632
rect 4456 81572 4460 81628
rect 4460 81572 4516 81628
rect 4516 81572 4520 81628
rect 4456 81568 4520 81572
rect 34936 81628 35000 81632
rect 34936 81572 34940 81628
rect 34940 81572 34996 81628
rect 34996 81572 35000 81628
rect 34936 81568 35000 81572
rect 35016 81628 35080 81632
rect 35016 81572 35020 81628
rect 35020 81572 35076 81628
rect 35076 81572 35080 81628
rect 35016 81568 35080 81572
rect 35096 81628 35160 81632
rect 35096 81572 35100 81628
rect 35100 81572 35156 81628
rect 35156 81572 35160 81628
rect 35096 81568 35160 81572
rect 35176 81628 35240 81632
rect 35176 81572 35180 81628
rect 35180 81572 35236 81628
rect 35236 81572 35240 81628
rect 35176 81568 35240 81572
rect 65656 81628 65720 81632
rect 65656 81572 65660 81628
rect 65660 81572 65716 81628
rect 65716 81572 65720 81628
rect 65656 81568 65720 81572
rect 65736 81628 65800 81632
rect 65736 81572 65740 81628
rect 65740 81572 65796 81628
rect 65796 81572 65800 81628
rect 65736 81568 65800 81572
rect 65816 81628 65880 81632
rect 65816 81572 65820 81628
rect 65820 81572 65876 81628
rect 65876 81572 65880 81628
rect 65816 81568 65880 81572
rect 65896 81628 65960 81632
rect 65896 81572 65900 81628
rect 65900 81572 65956 81628
rect 65956 81572 65960 81628
rect 65896 81568 65960 81572
rect 96376 81628 96440 81632
rect 96376 81572 96380 81628
rect 96380 81572 96436 81628
rect 96436 81572 96440 81628
rect 96376 81568 96440 81572
rect 96456 81628 96520 81632
rect 96456 81572 96460 81628
rect 96460 81572 96516 81628
rect 96516 81572 96520 81628
rect 96456 81568 96520 81572
rect 96536 81628 96600 81632
rect 96536 81572 96540 81628
rect 96540 81572 96596 81628
rect 96596 81572 96600 81628
rect 96536 81568 96600 81572
rect 96616 81628 96680 81632
rect 96616 81572 96620 81628
rect 96620 81572 96676 81628
rect 96676 81572 96680 81628
rect 96616 81568 96680 81572
rect 19576 81084 19640 81088
rect 19576 81028 19580 81084
rect 19580 81028 19636 81084
rect 19636 81028 19640 81084
rect 19576 81024 19640 81028
rect 19656 81084 19720 81088
rect 19656 81028 19660 81084
rect 19660 81028 19716 81084
rect 19716 81028 19720 81084
rect 19656 81024 19720 81028
rect 19736 81084 19800 81088
rect 19736 81028 19740 81084
rect 19740 81028 19796 81084
rect 19796 81028 19800 81084
rect 19736 81024 19800 81028
rect 19816 81084 19880 81088
rect 19816 81028 19820 81084
rect 19820 81028 19876 81084
rect 19876 81028 19880 81084
rect 19816 81024 19880 81028
rect 50296 81084 50360 81088
rect 50296 81028 50300 81084
rect 50300 81028 50356 81084
rect 50356 81028 50360 81084
rect 50296 81024 50360 81028
rect 50376 81084 50440 81088
rect 50376 81028 50380 81084
rect 50380 81028 50436 81084
rect 50436 81028 50440 81084
rect 50376 81024 50440 81028
rect 50456 81084 50520 81088
rect 50456 81028 50460 81084
rect 50460 81028 50516 81084
rect 50516 81028 50520 81084
rect 50456 81024 50520 81028
rect 50536 81084 50600 81088
rect 50536 81028 50540 81084
rect 50540 81028 50596 81084
rect 50596 81028 50600 81084
rect 50536 81024 50600 81028
rect 81016 81084 81080 81088
rect 81016 81028 81020 81084
rect 81020 81028 81076 81084
rect 81076 81028 81080 81084
rect 81016 81024 81080 81028
rect 81096 81084 81160 81088
rect 81096 81028 81100 81084
rect 81100 81028 81156 81084
rect 81156 81028 81160 81084
rect 81096 81024 81160 81028
rect 81176 81084 81240 81088
rect 81176 81028 81180 81084
rect 81180 81028 81236 81084
rect 81236 81028 81240 81084
rect 81176 81024 81240 81028
rect 81256 81084 81320 81088
rect 81256 81028 81260 81084
rect 81260 81028 81316 81084
rect 81316 81028 81320 81084
rect 81256 81024 81320 81028
rect 4216 80540 4280 80544
rect 4216 80484 4220 80540
rect 4220 80484 4276 80540
rect 4276 80484 4280 80540
rect 4216 80480 4280 80484
rect 4296 80540 4360 80544
rect 4296 80484 4300 80540
rect 4300 80484 4356 80540
rect 4356 80484 4360 80540
rect 4296 80480 4360 80484
rect 4376 80540 4440 80544
rect 4376 80484 4380 80540
rect 4380 80484 4436 80540
rect 4436 80484 4440 80540
rect 4376 80480 4440 80484
rect 4456 80540 4520 80544
rect 4456 80484 4460 80540
rect 4460 80484 4516 80540
rect 4516 80484 4520 80540
rect 4456 80480 4520 80484
rect 34936 80540 35000 80544
rect 34936 80484 34940 80540
rect 34940 80484 34996 80540
rect 34996 80484 35000 80540
rect 34936 80480 35000 80484
rect 35016 80540 35080 80544
rect 35016 80484 35020 80540
rect 35020 80484 35076 80540
rect 35076 80484 35080 80540
rect 35016 80480 35080 80484
rect 35096 80540 35160 80544
rect 35096 80484 35100 80540
rect 35100 80484 35156 80540
rect 35156 80484 35160 80540
rect 35096 80480 35160 80484
rect 35176 80540 35240 80544
rect 35176 80484 35180 80540
rect 35180 80484 35236 80540
rect 35236 80484 35240 80540
rect 35176 80480 35240 80484
rect 65656 80540 65720 80544
rect 65656 80484 65660 80540
rect 65660 80484 65716 80540
rect 65716 80484 65720 80540
rect 65656 80480 65720 80484
rect 65736 80540 65800 80544
rect 65736 80484 65740 80540
rect 65740 80484 65796 80540
rect 65796 80484 65800 80540
rect 65736 80480 65800 80484
rect 65816 80540 65880 80544
rect 65816 80484 65820 80540
rect 65820 80484 65876 80540
rect 65876 80484 65880 80540
rect 65816 80480 65880 80484
rect 65896 80540 65960 80544
rect 65896 80484 65900 80540
rect 65900 80484 65956 80540
rect 65956 80484 65960 80540
rect 65896 80480 65960 80484
rect 96376 80540 96440 80544
rect 96376 80484 96380 80540
rect 96380 80484 96436 80540
rect 96436 80484 96440 80540
rect 96376 80480 96440 80484
rect 96456 80540 96520 80544
rect 96456 80484 96460 80540
rect 96460 80484 96516 80540
rect 96516 80484 96520 80540
rect 96456 80480 96520 80484
rect 96536 80540 96600 80544
rect 96536 80484 96540 80540
rect 96540 80484 96596 80540
rect 96596 80484 96600 80540
rect 96536 80480 96600 80484
rect 96616 80540 96680 80544
rect 96616 80484 96620 80540
rect 96620 80484 96676 80540
rect 96676 80484 96680 80540
rect 96616 80480 96680 80484
rect 19576 79996 19640 80000
rect 19576 79940 19580 79996
rect 19580 79940 19636 79996
rect 19636 79940 19640 79996
rect 19576 79936 19640 79940
rect 19656 79996 19720 80000
rect 19656 79940 19660 79996
rect 19660 79940 19716 79996
rect 19716 79940 19720 79996
rect 19656 79936 19720 79940
rect 19736 79996 19800 80000
rect 19736 79940 19740 79996
rect 19740 79940 19796 79996
rect 19796 79940 19800 79996
rect 19736 79936 19800 79940
rect 19816 79996 19880 80000
rect 19816 79940 19820 79996
rect 19820 79940 19876 79996
rect 19876 79940 19880 79996
rect 19816 79936 19880 79940
rect 50296 79996 50360 80000
rect 50296 79940 50300 79996
rect 50300 79940 50356 79996
rect 50356 79940 50360 79996
rect 50296 79936 50360 79940
rect 50376 79996 50440 80000
rect 50376 79940 50380 79996
rect 50380 79940 50436 79996
rect 50436 79940 50440 79996
rect 50376 79936 50440 79940
rect 50456 79996 50520 80000
rect 50456 79940 50460 79996
rect 50460 79940 50516 79996
rect 50516 79940 50520 79996
rect 50456 79936 50520 79940
rect 50536 79996 50600 80000
rect 50536 79940 50540 79996
rect 50540 79940 50596 79996
rect 50596 79940 50600 79996
rect 50536 79936 50600 79940
rect 81016 79996 81080 80000
rect 81016 79940 81020 79996
rect 81020 79940 81076 79996
rect 81076 79940 81080 79996
rect 81016 79936 81080 79940
rect 81096 79996 81160 80000
rect 81096 79940 81100 79996
rect 81100 79940 81156 79996
rect 81156 79940 81160 79996
rect 81096 79936 81160 79940
rect 81176 79996 81240 80000
rect 81176 79940 81180 79996
rect 81180 79940 81236 79996
rect 81236 79940 81240 79996
rect 81176 79936 81240 79940
rect 81256 79996 81320 80000
rect 81256 79940 81260 79996
rect 81260 79940 81316 79996
rect 81316 79940 81320 79996
rect 81256 79936 81320 79940
rect 4216 79452 4280 79456
rect 4216 79396 4220 79452
rect 4220 79396 4276 79452
rect 4276 79396 4280 79452
rect 4216 79392 4280 79396
rect 4296 79452 4360 79456
rect 4296 79396 4300 79452
rect 4300 79396 4356 79452
rect 4356 79396 4360 79452
rect 4296 79392 4360 79396
rect 4376 79452 4440 79456
rect 4376 79396 4380 79452
rect 4380 79396 4436 79452
rect 4436 79396 4440 79452
rect 4376 79392 4440 79396
rect 4456 79452 4520 79456
rect 4456 79396 4460 79452
rect 4460 79396 4516 79452
rect 4516 79396 4520 79452
rect 4456 79392 4520 79396
rect 34936 79452 35000 79456
rect 34936 79396 34940 79452
rect 34940 79396 34996 79452
rect 34996 79396 35000 79452
rect 34936 79392 35000 79396
rect 35016 79452 35080 79456
rect 35016 79396 35020 79452
rect 35020 79396 35076 79452
rect 35076 79396 35080 79452
rect 35016 79392 35080 79396
rect 35096 79452 35160 79456
rect 35096 79396 35100 79452
rect 35100 79396 35156 79452
rect 35156 79396 35160 79452
rect 35096 79392 35160 79396
rect 35176 79452 35240 79456
rect 35176 79396 35180 79452
rect 35180 79396 35236 79452
rect 35236 79396 35240 79452
rect 35176 79392 35240 79396
rect 65656 79452 65720 79456
rect 65656 79396 65660 79452
rect 65660 79396 65716 79452
rect 65716 79396 65720 79452
rect 65656 79392 65720 79396
rect 65736 79452 65800 79456
rect 65736 79396 65740 79452
rect 65740 79396 65796 79452
rect 65796 79396 65800 79452
rect 65736 79392 65800 79396
rect 65816 79452 65880 79456
rect 65816 79396 65820 79452
rect 65820 79396 65876 79452
rect 65876 79396 65880 79452
rect 65816 79392 65880 79396
rect 65896 79452 65960 79456
rect 65896 79396 65900 79452
rect 65900 79396 65956 79452
rect 65956 79396 65960 79452
rect 65896 79392 65960 79396
rect 96376 79452 96440 79456
rect 96376 79396 96380 79452
rect 96380 79396 96436 79452
rect 96436 79396 96440 79452
rect 96376 79392 96440 79396
rect 96456 79452 96520 79456
rect 96456 79396 96460 79452
rect 96460 79396 96516 79452
rect 96516 79396 96520 79452
rect 96456 79392 96520 79396
rect 96536 79452 96600 79456
rect 96536 79396 96540 79452
rect 96540 79396 96596 79452
rect 96596 79396 96600 79452
rect 96536 79392 96600 79396
rect 96616 79452 96680 79456
rect 96616 79396 96620 79452
rect 96620 79396 96676 79452
rect 96676 79396 96680 79452
rect 96616 79392 96680 79396
rect 19576 78908 19640 78912
rect 19576 78852 19580 78908
rect 19580 78852 19636 78908
rect 19636 78852 19640 78908
rect 19576 78848 19640 78852
rect 19656 78908 19720 78912
rect 19656 78852 19660 78908
rect 19660 78852 19716 78908
rect 19716 78852 19720 78908
rect 19656 78848 19720 78852
rect 19736 78908 19800 78912
rect 19736 78852 19740 78908
rect 19740 78852 19796 78908
rect 19796 78852 19800 78908
rect 19736 78848 19800 78852
rect 19816 78908 19880 78912
rect 19816 78852 19820 78908
rect 19820 78852 19876 78908
rect 19876 78852 19880 78908
rect 19816 78848 19880 78852
rect 50296 78908 50360 78912
rect 50296 78852 50300 78908
rect 50300 78852 50356 78908
rect 50356 78852 50360 78908
rect 50296 78848 50360 78852
rect 50376 78908 50440 78912
rect 50376 78852 50380 78908
rect 50380 78852 50436 78908
rect 50436 78852 50440 78908
rect 50376 78848 50440 78852
rect 50456 78908 50520 78912
rect 50456 78852 50460 78908
rect 50460 78852 50516 78908
rect 50516 78852 50520 78908
rect 50456 78848 50520 78852
rect 50536 78908 50600 78912
rect 50536 78852 50540 78908
rect 50540 78852 50596 78908
rect 50596 78852 50600 78908
rect 50536 78848 50600 78852
rect 81016 78908 81080 78912
rect 81016 78852 81020 78908
rect 81020 78852 81076 78908
rect 81076 78852 81080 78908
rect 81016 78848 81080 78852
rect 81096 78908 81160 78912
rect 81096 78852 81100 78908
rect 81100 78852 81156 78908
rect 81156 78852 81160 78908
rect 81096 78848 81160 78852
rect 81176 78908 81240 78912
rect 81176 78852 81180 78908
rect 81180 78852 81236 78908
rect 81236 78852 81240 78908
rect 81176 78848 81240 78852
rect 81256 78908 81320 78912
rect 81256 78852 81260 78908
rect 81260 78852 81316 78908
rect 81316 78852 81320 78908
rect 81256 78848 81320 78852
rect 4216 78364 4280 78368
rect 4216 78308 4220 78364
rect 4220 78308 4276 78364
rect 4276 78308 4280 78364
rect 4216 78304 4280 78308
rect 4296 78364 4360 78368
rect 4296 78308 4300 78364
rect 4300 78308 4356 78364
rect 4356 78308 4360 78364
rect 4296 78304 4360 78308
rect 4376 78364 4440 78368
rect 4376 78308 4380 78364
rect 4380 78308 4436 78364
rect 4436 78308 4440 78364
rect 4376 78304 4440 78308
rect 4456 78364 4520 78368
rect 4456 78308 4460 78364
rect 4460 78308 4516 78364
rect 4516 78308 4520 78364
rect 4456 78304 4520 78308
rect 34936 78364 35000 78368
rect 34936 78308 34940 78364
rect 34940 78308 34996 78364
rect 34996 78308 35000 78364
rect 34936 78304 35000 78308
rect 35016 78364 35080 78368
rect 35016 78308 35020 78364
rect 35020 78308 35076 78364
rect 35076 78308 35080 78364
rect 35016 78304 35080 78308
rect 35096 78364 35160 78368
rect 35096 78308 35100 78364
rect 35100 78308 35156 78364
rect 35156 78308 35160 78364
rect 35096 78304 35160 78308
rect 35176 78364 35240 78368
rect 35176 78308 35180 78364
rect 35180 78308 35236 78364
rect 35236 78308 35240 78364
rect 35176 78304 35240 78308
rect 65656 78364 65720 78368
rect 65656 78308 65660 78364
rect 65660 78308 65716 78364
rect 65716 78308 65720 78364
rect 65656 78304 65720 78308
rect 65736 78364 65800 78368
rect 65736 78308 65740 78364
rect 65740 78308 65796 78364
rect 65796 78308 65800 78364
rect 65736 78304 65800 78308
rect 65816 78364 65880 78368
rect 65816 78308 65820 78364
rect 65820 78308 65876 78364
rect 65876 78308 65880 78364
rect 65816 78304 65880 78308
rect 65896 78364 65960 78368
rect 65896 78308 65900 78364
rect 65900 78308 65956 78364
rect 65956 78308 65960 78364
rect 65896 78304 65960 78308
rect 96376 78364 96440 78368
rect 96376 78308 96380 78364
rect 96380 78308 96436 78364
rect 96436 78308 96440 78364
rect 96376 78304 96440 78308
rect 96456 78364 96520 78368
rect 96456 78308 96460 78364
rect 96460 78308 96516 78364
rect 96516 78308 96520 78364
rect 96456 78304 96520 78308
rect 96536 78364 96600 78368
rect 96536 78308 96540 78364
rect 96540 78308 96596 78364
rect 96596 78308 96600 78364
rect 96536 78304 96600 78308
rect 96616 78364 96680 78368
rect 96616 78308 96620 78364
rect 96620 78308 96676 78364
rect 96676 78308 96680 78364
rect 96616 78304 96680 78308
rect 19576 77820 19640 77824
rect 19576 77764 19580 77820
rect 19580 77764 19636 77820
rect 19636 77764 19640 77820
rect 19576 77760 19640 77764
rect 19656 77820 19720 77824
rect 19656 77764 19660 77820
rect 19660 77764 19716 77820
rect 19716 77764 19720 77820
rect 19656 77760 19720 77764
rect 19736 77820 19800 77824
rect 19736 77764 19740 77820
rect 19740 77764 19796 77820
rect 19796 77764 19800 77820
rect 19736 77760 19800 77764
rect 19816 77820 19880 77824
rect 19816 77764 19820 77820
rect 19820 77764 19876 77820
rect 19876 77764 19880 77820
rect 19816 77760 19880 77764
rect 50296 77820 50360 77824
rect 50296 77764 50300 77820
rect 50300 77764 50356 77820
rect 50356 77764 50360 77820
rect 50296 77760 50360 77764
rect 50376 77820 50440 77824
rect 50376 77764 50380 77820
rect 50380 77764 50436 77820
rect 50436 77764 50440 77820
rect 50376 77760 50440 77764
rect 50456 77820 50520 77824
rect 50456 77764 50460 77820
rect 50460 77764 50516 77820
rect 50516 77764 50520 77820
rect 50456 77760 50520 77764
rect 50536 77820 50600 77824
rect 50536 77764 50540 77820
rect 50540 77764 50596 77820
rect 50596 77764 50600 77820
rect 50536 77760 50600 77764
rect 81016 77820 81080 77824
rect 81016 77764 81020 77820
rect 81020 77764 81076 77820
rect 81076 77764 81080 77820
rect 81016 77760 81080 77764
rect 81096 77820 81160 77824
rect 81096 77764 81100 77820
rect 81100 77764 81156 77820
rect 81156 77764 81160 77820
rect 81096 77760 81160 77764
rect 81176 77820 81240 77824
rect 81176 77764 81180 77820
rect 81180 77764 81236 77820
rect 81236 77764 81240 77820
rect 81176 77760 81240 77764
rect 81256 77820 81320 77824
rect 81256 77764 81260 77820
rect 81260 77764 81316 77820
rect 81316 77764 81320 77820
rect 81256 77760 81320 77764
rect 4216 77276 4280 77280
rect 4216 77220 4220 77276
rect 4220 77220 4276 77276
rect 4276 77220 4280 77276
rect 4216 77216 4280 77220
rect 4296 77276 4360 77280
rect 4296 77220 4300 77276
rect 4300 77220 4356 77276
rect 4356 77220 4360 77276
rect 4296 77216 4360 77220
rect 4376 77276 4440 77280
rect 4376 77220 4380 77276
rect 4380 77220 4436 77276
rect 4436 77220 4440 77276
rect 4376 77216 4440 77220
rect 4456 77276 4520 77280
rect 4456 77220 4460 77276
rect 4460 77220 4516 77276
rect 4516 77220 4520 77276
rect 4456 77216 4520 77220
rect 34936 77276 35000 77280
rect 34936 77220 34940 77276
rect 34940 77220 34996 77276
rect 34996 77220 35000 77276
rect 34936 77216 35000 77220
rect 35016 77276 35080 77280
rect 35016 77220 35020 77276
rect 35020 77220 35076 77276
rect 35076 77220 35080 77276
rect 35016 77216 35080 77220
rect 35096 77276 35160 77280
rect 35096 77220 35100 77276
rect 35100 77220 35156 77276
rect 35156 77220 35160 77276
rect 35096 77216 35160 77220
rect 35176 77276 35240 77280
rect 35176 77220 35180 77276
rect 35180 77220 35236 77276
rect 35236 77220 35240 77276
rect 35176 77216 35240 77220
rect 65656 77276 65720 77280
rect 65656 77220 65660 77276
rect 65660 77220 65716 77276
rect 65716 77220 65720 77276
rect 65656 77216 65720 77220
rect 65736 77276 65800 77280
rect 65736 77220 65740 77276
rect 65740 77220 65796 77276
rect 65796 77220 65800 77276
rect 65736 77216 65800 77220
rect 65816 77276 65880 77280
rect 65816 77220 65820 77276
rect 65820 77220 65876 77276
rect 65876 77220 65880 77276
rect 65816 77216 65880 77220
rect 65896 77276 65960 77280
rect 65896 77220 65900 77276
rect 65900 77220 65956 77276
rect 65956 77220 65960 77276
rect 65896 77216 65960 77220
rect 96376 77276 96440 77280
rect 96376 77220 96380 77276
rect 96380 77220 96436 77276
rect 96436 77220 96440 77276
rect 96376 77216 96440 77220
rect 96456 77276 96520 77280
rect 96456 77220 96460 77276
rect 96460 77220 96516 77276
rect 96516 77220 96520 77276
rect 96456 77216 96520 77220
rect 96536 77276 96600 77280
rect 96536 77220 96540 77276
rect 96540 77220 96596 77276
rect 96596 77220 96600 77276
rect 96536 77216 96600 77220
rect 96616 77276 96680 77280
rect 96616 77220 96620 77276
rect 96620 77220 96676 77276
rect 96676 77220 96680 77276
rect 96616 77216 96680 77220
rect 19576 76732 19640 76736
rect 19576 76676 19580 76732
rect 19580 76676 19636 76732
rect 19636 76676 19640 76732
rect 19576 76672 19640 76676
rect 19656 76732 19720 76736
rect 19656 76676 19660 76732
rect 19660 76676 19716 76732
rect 19716 76676 19720 76732
rect 19656 76672 19720 76676
rect 19736 76732 19800 76736
rect 19736 76676 19740 76732
rect 19740 76676 19796 76732
rect 19796 76676 19800 76732
rect 19736 76672 19800 76676
rect 19816 76732 19880 76736
rect 19816 76676 19820 76732
rect 19820 76676 19876 76732
rect 19876 76676 19880 76732
rect 19816 76672 19880 76676
rect 50296 76732 50360 76736
rect 50296 76676 50300 76732
rect 50300 76676 50356 76732
rect 50356 76676 50360 76732
rect 50296 76672 50360 76676
rect 50376 76732 50440 76736
rect 50376 76676 50380 76732
rect 50380 76676 50436 76732
rect 50436 76676 50440 76732
rect 50376 76672 50440 76676
rect 50456 76732 50520 76736
rect 50456 76676 50460 76732
rect 50460 76676 50516 76732
rect 50516 76676 50520 76732
rect 50456 76672 50520 76676
rect 50536 76732 50600 76736
rect 50536 76676 50540 76732
rect 50540 76676 50596 76732
rect 50596 76676 50600 76732
rect 50536 76672 50600 76676
rect 81016 76732 81080 76736
rect 81016 76676 81020 76732
rect 81020 76676 81076 76732
rect 81076 76676 81080 76732
rect 81016 76672 81080 76676
rect 81096 76732 81160 76736
rect 81096 76676 81100 76732
rect 81100 76676 81156 76732
rect 81156 76676 81160 76732
rect 81096 76672 81160 76676
rect 81176 76732 81240 76736
rect 81176 76676 81180 76732
rect 81180 76676 81236 76732
rect 81236 76676 81240 76732
rect 81176 76672 81240 76676
rect 81256 76732 81320 76736
rect 81256 76676 81260 76732
rect 81260 76676 81316 76732
rect 81316 76676 81320 76732
rect 81256 76672 81320 76676
rect 4216 76188 4280 76192
rect 4216 76132 4220 76188
rect 4220 76132 4276 76188
rect 4276 76132 4280 76188
rect 4216 76128 4280 76132
rect 4296 76188 4360 76192
rect 4296 76132 4300 76188
rect 4300 76132 4356 76188
rect 4356 76132 4360 76188
rect 4296 76128 4360 76132
rect 4376 76188 4440 76192
rect 4376 76132 4380 76188
rect 4380 76132 4436 76188
rect 4436 76132 4440 76188
rect 4376 76128 4440 76132
rect 4456 76188 4520 76192
rect 4456 76132 4460 76188
rect 4460 76132 4516 76188
rect 4516 76132 4520 76188
rect 4456 76128 4520 76132
rect 34936 76188 35000 76192
rect 34936 76132 34940 76188
rect 34940 76132 34996 76188
rect 34996 76132 35000 76188
rect 34936 76128 35000 76132
rect 35016 76188 35080 76192
rect 35016 76132 35020 76188
rect 35020 76132 35076 76188
rect 35076 76132 35080 76188
rect 35016 76128 35080 76132
rect 35096 76188 35160 76192
rect 35096 76132 35100 76188
rect 35100 76132 35156 76188
rect 35156 76132 35160 76188
rect 35096 76128 35160 76132
rect 35176 76188 35240 76192
rect 35176 76132 35180 76188
rect 35180 76132 35236 76188
rect 35236 76132 35240 76188
rect 35176 76128 35240 76132
rect 65656 76188 65720 76192
rect 65656 76132 65660 76188
rect 65660 76132 65716 76188
rect 65716 76132 65720 76188
rect 65656 76128 65720 76132
rect 65736 76188 65800 76192
rect 65736 76132 65740 76188
rect 65740 76132 65796 76188
rect 65796 76132 65800 76188
rect 65736 76128 65800 76132
rect 65816 76188 65880 76192
rect 65816 76132 65820 76188
rect 65820 76132 65876 76188
rect 65876 76132 65880 76188
rect 65816 76128 65880 76132
rect 65896 76188 65960 76192
rect 65896 76132 65900 76188
rect 65900 76132 65956 76188
rect 65956 76132 65960 76188
rect 65896 76128 65960 76132
rect 96376 76188 96440 76192
rect 96376 76132 96380 76188
rect 96380 76132 96436 76188
rect 96436 76132 96440 76188
rect 96376 76128 96440 76132
rect 96456 76188 96520 76192
rect 96456 76132 96460 76188
rect 96460 76132 96516 76188
rect 96516 76132 96520 76188
rect 96456 76128 96520 76132
rect 96536 76188 96600 76192
rect 96536 76132 96540 76188
rect 96540 76132 96596 76188
rect 96596 76132 96600 76188
rect 96536 76128 96600 76132
rect 96616 76188 96680 76192
rect 96616 76132 96620 76188
rect 96620 76132 96676 76188
rect 96676 76132 96680 76188
rect 96616 76128 96680 76132
rect 19576 75644 19640 75648
rect 19576 75588 19580 75644
rect 19580 75588 19636 75644
rect 19636 75588 19640 75644
rect 19576 75584 19640 75588
rect 19656 75644 19720 75648
rect 19656 75588 19660 75644
rect 19660 75588 19716 75644
rect 19716 75588 19720 75644
rect 19656 75584 19720 75588
rect 19736 75644 19800 75648
rect 19736 75588 19740 75644
rect 19740 75588 19796 75644
rect 19796 75588 19800 75644
rect 19736 75584 19800 75588
rect 19816 75644 19880 75648
rect 19816 75588 19820 75644
rect 19820 75588 19876 75644
rect 19876 75588 19880 75644
rect 19816 75584 19880 75588
rect 50296 75644 50360 75648
rect 50296 75588 50300 75644
rect 50300 75588 50356 75644
rect 50356 75588 50360 75644
rect 50296 75584 50360 75588
rect 50376 75644 50440 75648
rect 50376 75588 50380 75644
rect 50380 75588 50436 75644
rect 50436 75588 50440 75644
rect 50376 75584 50440 75588
rect 50456 75644 50520 75648
rect 50456 75588 50460 75644
rect 50460 75588 50516 75644
rect 50516 75588 50520 75644
rect 50456 75584 50520 75588
rect 50536 75644 50600 75648
rect 50536 75588 50540 75644
rect 50540 75588 50596 75644
rect 50596 75588 50600 75644
rect 50536 75584 50600 75588
rect 81016 75644 81080 75648
rect 81016 75588 81020 75644
rect 81020 75588 81076 75644
rect 81076 75588 81080 75644
rect 81016 75584 81080 75588
rect 81096 75644 81160 75648
rect 81096 75588 81100 75644
rect 81100 75588 81156 75644
rect 81156 75588 81160 75644
rect 81096 75584 81160 75588
rect 81176 75644 81240 75648
rect 81176 75588 81180 75644
rect 81180 75588 81236 75644
rect 81236 75588 81240 75644
rect 81176 75584 81240 75588
rect 81256 75644 81320 75648
rect 81256 75588 81260 75644
rect 81260 75588 81316 75644
rect 81316 75588 81320 75644
rect 81256 75584 81320 75588
rect 4216 75100 4280 75104
rect 4216 75044 4220 75100
rect 4220 75044 4276 75100
rect 4276 75044 4280 75100
rect 4216 75040 4280 75044
rect 4296 75100 4360 75104
rect 4296 75044 4300 75100
rect 4300 75044 4356 75100
rect 4356 75044 4360 75100
rect 4296 75040 4360 75044
rect 4376 75100 4440 75104
rect 4376 75044 4380 75100
rect 4380 75044 4436 75100
rect 4436 75044 4440 75100
rect 4376 75040 4440 75044
rect 4456 75100 4520 75104
rect 4456 75044 4460 75100
rect 4460 75044 4516 75100
rect 4516 75044 4520 75100
rect 4456 75040 4520 75044
rect 34936 75100 35000 75104
rect 34936 75044 34940 75100
rect 34940 75044 34996 75100
rect 34996 75044 35000 75100
rect 34936 75040 35000 75044
rect 35016 75100 35080 75104
rect 35016 75044 35020 75100
rect 35020 75044 35076 75100
rect 35076 75044 35080 75100
rect 35016 75040 35080 75044
rect 35096 75100 35160 75104
rect 35096 75044 35100 75100
rect 35100 75044 35156 75100
rect 35156 75044 35160 75100
rect 35096 75040 35160 75044
rect 35176 75100 35240 75104
rect 35176 75044 35180 75100
rect 35180 75044 35236 75100
rect 35236 75044 35240 75100
rect 35176 75040 35240 75044
rect 65656 75100 65720 75104
rect 65656 75044 65660 75100
rect 65660 75044 65716 75100
rect 65716 75044 65720 75100
rect 65656 75040 65720 75044
rect 65736 75100 65800 75104
rect 65736 75044 65740 75100
rect 65740 75044 65796 75100
rect 65796 75044 65800 75100
rect 65736 75040 65800 75044
rect 65816 75100 65880 75104
rect 65816 75044 65820 75100
rect 65820 75044 65876 75100
rect 65876 75044 65880 75100
rect 65816 75040 65880 75044
rect 65896 75100 65960 75104
rect 65896 75044 65900 75100
rect 65900 75044 65956 75100
rect 65956 75044 65960 75100
rect 65896 75040 65960 75044
rect 96376 75100 96440 75104
rect 96376 75044 96380 75100
rect 96380 75044 96436 75100
rect 96436 75044 96440 75100
rect 96376 75040 96440 75044
rect 96456 75100 96520 75104
rect 96456 75044 96460 75100
rect 96460 75044 96516 75100
rect 96516 75044 96520 75100
rect 96456 75040 96520 75044
rect 96536 75100 96600 75104
rect 96536 75044 96540 75100
rect 96540 75044 96596 75100
rect 96596 75044 96600 75100
rect 96536 75040 96600 75044
rect 96616 75100 96680 75104
rect 96616 75044 96620 75100
rect 96620 75044 96676 75100
rect 96676 75044 96680 75100
rect 96616 75040 96680 75044
rect 19576 74556 19640 74560
rect 19576 74500 19580 74556
rect 19580 74500 19636 74556
rect 19636 74500 19640 74556
rect 19576 74496 19640 74500
rect 19656 74556 19720 74560
rect 19656 74500 19660 74556
rect 19660 74500 19716 74556
rect 19716 74500 19720 74556
rect 19656 74496 19720 74500
rect 19736 74556 19800 74560
rect 19736 74500 19740 74556
rect 19740 74500 19796 74556
rect 19796 74500 19800 74556
rect 19736 74496 19800 74500
rect 19816 74556 19880 74560
rect 19816 74500 19820 74556
rect 19820 74500 19876 74556
rect 19876 74500 19880 74556
rect 19816 74496 19880 74500
rect 50296 74556 50360 74560
rect 50296 74500 50300 74556
rect 50300 74500 50356 74556
rect 50356 74500 50360 74556
rect 50296 74496 50360 74500
rect 50376 74556 50440 74560
rect 50376 74500 50380 74556
rect 50380 74500 50436 74556
rect 50436 74500 50440 74556
rect 50376 74496 50440 74500
rect 50456 74556 50520 74560
rect 50456 74500 50460 74556
rect 50460 74500 50516 74556
rect 50516 74500 50520 74556
rect 50456 74496 50520 74500
rect 50536 74556 50600 74560
rect 50536 74500 50540 74556
rect 50540 74500 50596 74556
rect 50596 74500 50600 74556
rect 50536 74496 50600 74500
rect 81016 74556 81080 74560
rect 81016 74500 81020 74556
rect 81020 74500 81076 74556
rect 81076 74500 81080 74556
rect 81016 74496 81080 74500
rect 81096 74556 81160 74560
rect 81096 74500 81100 74556
rect 81100 74500 81156 74556
rect 81156 74500 81160 74556
rect 81096 74496 81160 74500
rect 81176 74556 81240 74560
rect 81176 74500 81180 74556
rect 81180 74500 81236 74556
rect 81236 74500 81240 74556
rect 81176 74496 81240 74500
rect 81256 74556 81320 74560
rect 81256 74500 81260 74556
rect 81260 74500 81316 74556
rect 81316 74500 81320 74556
rect 81256 74496 81320 74500
rect 4216 74012 4280 74016
rect 4216 73956 4220 74012
rect 4220 73956 4276 74012
rect 4276 73956 4280 74012
rect 4216 73952 4280 73956
rect 4296 74012 4360 74016
rect 4296 73956 4300 74012
rect 4300 73956 4356 74012
rect 4356 73956 4360 74012
rect 4296 73952 4360 73956
rect 4376 74012 4440 74016
rect 4376 73956 4380 74012
rect 4380 73956 4436 74012
rect 4436 73956 4440 74012
rect 4376 73952 4440 73956
rect 4456 74012 4520 74016
rect 4456 73956 4460 74012
rect 4460 73956 4516 74012
rect 4516 73956 4520 74012
rect 4456 73952 4520 73956
rect 34936 74012 35000 74016
rect 34936 73956 34940 74012
rect 34940 73956 34996 74012
rect 34996 73956 35000 74012
rect 34936 73952 35000 73956
rect 35016 74012 35080 74016
rect 35016 73956 35020 74012
rect 35020 73956 35076 74012
rect 35076 73956 35080 74012
rect 35016 73952 35080 73956
rect 35096 74012 35160 74016
rect 35096 73956 35100 74012
rect 35100 73956 35156 74012
rect 35156 73956 35160 74012
rect 35096 73952 35160 73956
rect 35176 74012 35240 74016
rect 35176 73956 35180 74012
rect 35180 73956 35236 74012
rect 35236 73956 35240 74012
rect 35176 73952 35240 73956
rect 65656 74012 65720 74016
rect 65656 73956 65660 74012
rect 65660 73956 65716 74012
rect 65716 73956 65720 74012
rect 65656 73952 65720 73956
rect 65736 74012 65800 74016
rect 65736 73956 65740 74012
rect 65740 73956 65796 74012
rect 65796 73956 65800 74012
rect 65736 73952 65800 73956
rect 65816 74012 65880 74016
rect 65816 73956 65820 74012
rect 65820 73956 65876 74012
rect 65876 73956 65880 74012
rect 65816 73952 65880 73956
rect 65896 74012 65960 74016
rect 65896 73956 65900 74012
rect 65900 73956 65956 74012
rect 65956 73956 65960 74012
rect 65896 73952 65960 73956
rect 96376 74012 96440 74016
rect 96376 73956 96380 74012
rect 96380 73956 96436 74012
rect 96436 73956 96440 74012
rect 96376 73952 96440 73956
rect 96456 74012 96520 74016
rect 96456 73956 96460 74012
rect 96460 73956 96516 74012
rect 96516 73956 96520 74012
rect 96456 73952 96520 73956
rect 96536 74012 96600 74016
rect 96536 73956 96540 74012
rect 96540 73956 96596 74012
rect 96596 73956 96600 74012
rect 96536 73952 96600 73956
rect 96616 74012 96680 74016
rect 96616 73956 96620 74012
rect 96620 73956 96676 74012
rect 96676 73956 96680 74012
rect 96616 73952 96680 73956
rect 19576 73468 19640 73472
rect 19576 73412 19580 73468
rect 19580 73412 19636 73468
rect 19636 73412 19640 73468
rect 19576 73408 19640 73412
rect 19656 73468 19720 73472
rect 19656 73412 19660 73468
rect 19660 73412 19716 73468
rect 19716 73412 19720 73468
rect 19656 73408 19720 73412
rect 19736 73468 19800 73472
rect 19736 73412 19740 73468
rect 19740 73412 19796 73468
rect 19796 73412 19800 73468
rect 19736 73408 19800 73412
rect 19816 73468 19880 73472
rect 19816 73412 19820 73468
rect 19820 73412 19876 73468
rect 19876 73412 19880 73468
rect 19816 73408 19880 73412
rect 50296 73468 50360 73472
rect 50296 73412 50300 73468
rect 50300 73412 50356 73468
rect 50356 73412 50360 73468
rect 50296 73408 50360 73412
rect 50376 73468 50440 73472
rect 50376 73412 50380 73468
rect 50380 73412 50436 73468
rect 50436 73412 50440 73468
rect 50376 73408 50440 73412
rect 50456 73468 50520 73472
rect 50456 73412 50460 73468
rect 50460 73412 50516 73468
rect 50516 73412 50520 73468
rect 50456 73408 50520 73412
rect 50536 73468 50600 73472
rect 50536 73412 50540 73468
rect 50540 73412 50596 73468
rect 50596 73412 50600 73468
rect 50536 73408 50600 73412
rect 81016 73468 81080 73472
rect 81016 73412 81020 73468
rect 81020 73412 81076 73468
rect 81076 73412 81080 73468
rect 81016 73408 81080 73412
rect 81096 73468 81160 73472
rect 81096 73412 81100 73468
rect 81100 73412 81156 73468
rect 81156 73412 81160 73468
rect 81096 73408 81160 73412
rect 81176 73468 81240 73472
rect 81176 73412 81180 73468
rect 81180 73412 81236 73468
rect 81236 73412 81240 73468
rect 81176 73408 81240 73412
rect 81256 73468 81320 73472
rect 81256 73412 81260 73468
rect 81260 73412 81316 73468
rect 81316 73412 81320 73468
rect 81256 73408 81320 73412
rect 4216 72924 4280 72928
rect 4216 72868 4220 72924
rect 4220 72868 4276 72924
rect 4276 72868 4280 72924
rect 4216 72864 4280 72868
rect 4296 72924 4360 72928
rect 4296 72868 4300 72924
rect 4300 72868 4356 72924
rect 4356 72868 4360 72924
rect 4296 72864 4360 72868
rect 4376 72924 4440 72928
rect 4376 72868 4380 72924
rect 4380 72868 4436 72924
rect 4436 72868 4440 72924
rect 4376 72864 4440 72868
rect 4456 72924 4520 72928
rect 4456 72868 4460 72924
rect 4460 72868 4516 72924
rect 4516 72868 4520 72924
rect 4456 72864 4520 72868
rect 34936 72924 35000 72928
rect 34936 72868 34940 72924
rect 34940 72868 34996 72924
rect 34996 72868 35000 72924
rect 34936 72864 35000 72868
rect 35016 72924 35080 72928
rect 35016 72868 35020 72924
rect 35020 72868 35076 72924
rect 35076 72868 35080 72924
rect 35016 72864 35080 72868
rect 35096 72924 35160 72928
rect 35096 72868 35100 72924
rect 35100 72868 35156 72924
rect 35156 72868 35160 72924
rect 35096 72864 35160 72868
rect 35176 72924 35240 72928
rect 35176 72868 35180 72924
rect 35180 72868 35236 72924
rect 35236 72868 35240 72924
rect 35176 72864 35240 72868
rect 65656 72924 65720 72928
rect 65656 72868 65660 72924
rect 65660 72868 65716 72924
rect 65716 72868 65720 72924
rect 65656 72864 65720 72868
rect 65736 72924 65800 72928
rect 65736 72868 65740 72924
rect 65740 72868 65796 72924
rect 65796 72868 65800 72924
rect 65736 72864 65800 72868
rect 65816 72924 65880 72928
rect 65816 72868 65820 72924
rect 65820 72868 65876 72924
rect 65876 72868 65880 72924
rect 65816 72864 65880 72868
rect 65896 72924 65960 72928
rect 65896 72868 65900 72924
rect 65900 72868 65956 72924
rect 65956 72868 65960 72924
rect 65896 72864 65960 72868
rect 96376 72924 96440 72928
rect 96376 72868 96380 72924
rect 96380 72868 96436 72924
rect 96436 72868 96440 72924
rect 96376 72864 96440 72868
rect 96456 72924 96520 72928
rect 96456 72868 96460 72924
rect 96460 72868 96516 72924
rect 96516 72868 96520 72924
rect 96456 72864 96520 72868
rect 96536 72924 96600 72928
rect 96536 72868 96540 72924
rect 96540 72868 96596 72924
rect 96596 72868 96600 72924
rect 96536 72864 96600 72868
rect 96616 72924 96680 72928
rect 96616 72868 96620 72924
rect 96620 72868 96676 72924
rect 96676 72868 96680 72924
rect 96616 72864 96680 72868
rect 19576 72380 19640 72384
rect 19576 72324 19580 72380
rect 19580 72324 19636 72380
rect 19636 72324 19640 72380
rect 19576 72320 19640 72324
rect 19656 72380 19720 72384
rect 19656 72324 19660 72380
rect 19660 72324 19716 72380
rect 19716 72324 19720 72380
rect 19656 72320 19720 72324
rect 19736 72380 19800 72384
rect 19736 72324 19740 72380
rect 19740 72324 19796 72380
rect 19796 72324 19800 72380
rect 19736 72320 19800 72324
rect 19816 72380 19880 72384
rect 19816 72324 19820 72380
rect 19820 72324 19876 72380
rect 19876 72324 19880 72380
rect 19816 72320 19880 72324
rect 50296 72380 50360 72384
rect 50296 72324 50300 72380
rect 50300 72324 50356 72380
rect 50356 72324 50360 72380
rect 50296 72320 50360 72324
rect 50376 72380 50440 72384
rect 50376 72324 50380 72380
rect 50380 72324 50436 72380
rect 50436 72324 50440 72380
rect 50376 72320 50440 72324
rect 50456 72380 50520 72384
rect 50456 72324 50460 72380
rect 50460 72324 50516 72380
rect 50516 72324 50520 72380
rect 50456 72320 50520 72324
rect 50536 72380 50600 72384
rect 50536 72324 50540 72380
rect 50540 72324 50596 72380
rect 50596 72324 50600 72380
rect 50536 72320 50600 72324
rect 81016 72380 81080 72384
rect 81016 72324 81020 72380
rect 81020 72324 81076 72380
rect 81076 72324 81080 72380
rect 81016 72320 81080 72324
rect 81096 72380 81160 72384
rect 81096 72324 81100 72380
rect 81100 72324 81156 72380
rect 81156 72324 81160 72380
rect 81096 72320 81160 72324
rect 81176 72380 81240 72384
rect 81176 72324 81180 72380
rect 81180 72324 81236 72380
rect 81236 72324 81240 72380
rect 81176 72320 81240 72324
rect 81256 72380 81320 72384
rect 81256 72324 81260 72380
rect 81260 72324 81316 72380
rect 81316 72324 81320 72380
rect 81256 72320 81320 72324
rect 4216 71836 4280 71840
rect 4216 71780 4220 71836
rect 4220 71780 4276 71836
rect 4276 71780 4280 71836
rect 4216 71776 4280 71780
rect 4296 71836 4360 71840
rect 4296 71780 4300 71836
rect 4300 71780 4356 71836
rect 4356 71780 4360 71836
rect 4296 71776 4360 71780
rect 4376 71836 4440 71840
rect 4376 71780 4380 71836
rect 4380 71780 4436 71836
rect 4436 71780 4440 71836
rect 4376 71776 4440 71780
rect 4456 71836 4520 71840
rect 4456 71780 4460 71836
rect 4460 71780 4516 71836
rect 4516 71780 4520 71836
rect 4456 71776 4520 71780
rect 34936 71836 35000 71840
rect 34936 71780 34940 71836
rect 34940 71780 34996 71836
rect 34996 71780 35000 71836
rect 34936 71776 35000 71780
rect 35016 71836 35080 71840
rect 35016 71780 35020 71836
rect 35020 71780 35076 71836
rect 35076 71780 35080 71836
rect 35016 71776 35080 71780
rect 35096 71836 35160 71840
rect 35096 71780 35100 71836
rect 35100 71780 35156 71836
rect 35156 71780 35160 71836
rect 35096 71776 35160 71780
rect 35176 71836 35240 71840
rect 35176 71780 35180 71836
rect 35180 71780 35236 71836
rect 35236 71780 35240 71836
rect 35176 71776 35240 71780
rect 65656 71836 65720 71840
rect 65656 71780 65660 71836
rect 65660 71780 65716 71836
rect 65716 71780 65720 71836
rect 65656 71776 65720 71780
rect 65736 71836 65800 71840
rect 65736 71780 65740 71836
rect 65740 71780 65796 71836
rect 65796 71780 65800 71836
rect 65736 71776 65800 71780
rect 65816 71836 65880 71840
rect 65816 71780 65820 71836
rect 65820 71780 65876 71836
rect 65876 71780 65880 71836
rect 65816 71776 65880 71780
rect 65896 71836 65960 71840
rect 65896 71780 65900 71836
rect 65900 71780 65956 71836
rect 65956 71780 65960 71836
rect 65896 71776 65960 71780
rect 96376 71836 96440 71840
rect 96376 71780 96380 71836
rect 96380 71780 96436 71836
rect 96436 71780 96440 71836
rect 96376 71776 96440 71780
rect 96456 71836 96520 71840
rect 96456 71780 96460 71836
rect 96460 71780 96516 71836
rect 96516 71780 96520 71836
rect 96456 71776 96520 71780
rect 96536 71836 96600 71840
rect 96536 71780 96540 71836
rect 96540 71780 96596 71836
rect 96596 71780 96600 71836
rect 96536 71776 96600 71780
rect 96616 71836 96680 71840
rect 96616 71780 96620 71836
rect 96620 71780 96676 71836
rect 96676 71780 96680 71836
rect 96616 71776 96680 71780
rect 19576 71292 19640 71296
rect 19576 71236 19580 71292
rect 19580 71236 19636 71292
rect 19636 71236 19640 71292
rect 19576 71232 19640 71236
rect 19656 71292 19720 71296
rect 19656 71236 19660 71292
rect 19660 71236 19716 71292
rect 19716 71236 19720 71292
rect 19656 71232 19720 71236
rect 19736 71292 19800 71296
rect 19736 71236 19740 71292
rect 19740 71236 19796 71292
rect 19796 71236 19800 71292
rect 19736 71232 19800 71236
rect 19816 71292 19880 71296
rect 19816 71236 19820 71292
rect 19820 71236 19876 71292
rect 19876 71236 19880 71292
rect 19816 71232 19880 71236
rect 50296 71292 50360 71296
rect 50296 71236 50300 71292
rect 50300 71236 50356 71292
rect 50356 71236 50360 71292
rect 50296 71232 50360 71236
rect 50376 71292 50440 71296
rect 50376 71236 50380 71292
rect 50380 71236 50436 71292
rect 50436 71236 50440 71292
rect 50376 71232 50440 71236
rect 50456 71292 50520 71296
rect 50456 71236 50460 71292
rect 50460 71236 50516 71292
rect 50516 71236 50520 71292
rect 50456 71232 50520 71236
rect 50536 71292 50600 71296
rect 50536 71236 50540 71292
rect 50540 71236 50596 71292
rect 50596 71236 50600 71292
rect 50536 71232 50600 71236
rect 81016 71292 81080 71296
rect 81016 71236 81020 71292
rect 81020 71236 81076 71292
rect 81076 71236 81080 71292
rect 81016 71232 81080 71236
rect 81096 71292 81160 71296
rect 81096 71236 81100 71292
rect 81100 71236 81156 71292
rect 81156 71236 81160 71292
rect 81096 71232 81160 71236
rect 81176 71292 81240 71296
rect 81176 71236 81180 71292
rect 81180 71236 81236 71292
rect 81236 71236 81240 71292
rect 81176 71232 81240 71236
rect 81256 71292 81320 71296
rect 81256 71236 81260 71292
rect 81260 71236 81316 71292
rect 81316 71236 81320 71292
rect 81256 71232 81320 71236
rect 4216 70748 4280 70752
rect 4216 70692 4220 70748
rect 4220 70692 4276 70748
rect 4276 70692 4280 70748
rect 4216 70688 4280 70692
rect 4296 70748 4360 70752
rect 4296 70692 4300 70748
rect 4300 70692 4356 70748
rect 4356 70692 4360 70748
rect 4296 70688 4360 70692
rect 4376 70748 4440 70752
rect 4376 70692 4380 70748
rect 4380 70692 4436 70748
rect 4436 70692 4440 70748
rect 4376 70688 4440 70692
rect 4456 70748 4520 70752
rect 4456 70692 4460 70748
rect 4460 70692 4516 70748
rect 4516 70692 4520 70748
rect 4456 70688 4520 70692
rect 34936 70748 35000 70752
rect 34936 70692 34940 70748
rect 34940 70692 34996 70748
rect 34996 70692 35000 70748
rect 34936 70688 35000 70692
rect 35016 70748 35080 70752
rect 35016 70692 35020 70748
rect 35020 70692 35076 70748
rect 35076 70692 35080 70748
rect 35016 70688 35080 70692
rect 35096 70748 35160 70752
rect 35096 70692 35100 70748
rect 35100 70692 35156 70748
rect 35156 70692 35160 70748
rect 35096 70688 35160 70692
rect 35176 70748 35240 70752
rect 35176 70692 35180 70748
rect 35180 70692 35236 70748
rect 35236 70692 35240 70748
rect 35176 70688 35240 70692
rect 65656 70748 65720 70752
rect 65656 70692 65660 70748
rect 65660 70692 65716 70748
rect 65716 70692 65720 70748
rect 65656 70688 65720 70692
rect 65736 70748 65800 70752
rect 65736 70692 65740 70748
rect 65740 70692 65796 70748
rect 65796 70692 65800 70748
rect 65736 70688 65800 70692
rect 65816 70748 65880 70752
rect 65816 70692 65820 70748
rect 65820 70692 65876 70748
rect 65876 70692 65880 70748
rect 65816 70688 65880 70692
rect 65896 70748 65960 70752
rect 65896 70692 65900 70748
rect 65900 70692 65956 70748
rect 65956 70692 65960 70748
rect 65896 70688 65960 70692
rect 96376 70748 96440 70752
rect 96376 70692 96380 70748
rect 96380 70692 96436 70748
rect 96436 70692 96440 70748
rect 96376 70688 96440 70692
rect 96456 70748 96520 70752
rect 96456 70692 96460 70748
rect 96460 70692 96516 70748
rect 96516 70692 96520 70748
rect 96456 70688 96520 70692
rect 96536 70748 96600 70752
rect 96536 70692 96540 70748
rect 96540 70692 96596 70748
rect 96596 70692 96600 70748
rect 96536 70688 96600 70692
rect 96616 70748 96680 70752
rect 96616 70692 96620 70748
rect 96620 70692 96676 70748
rect 96676 70692 96680 70748
rect 96616 70688 96680 70692
rect 19576 70204 19640 70208
rect 19576 70148 19580 70204
rect 19580 70148 19636 70204
rect 19636 70148 19640 70204
rect 19576 70144 19640 70148
rect 19656 70204 19720 70208
rect 19656 70148 19660 70204
rect 19660 70148 19716 70204
rect 19716 70148 19720 70204
rect 19656 70144 19720 70148
rect 19736 70204 19800 70208
rect 19736 70148 19740 70204
rect 19740 70148 19796 70204
rect 19796 70148 19800 70204
rect 19736 70144 19800 70148
rect 19816 70204 19880 70208
rect 19816 70148 19820 70204
rect 19820 70148 19876 70204
rect 19876 70148 19880 70204
rect 19816 70144 19880 70148
rect 50296 70204 50360 70208
rect 50296 70148 50300 70204
rect 50300 70148 50356 70204
rect 50356 70148 50360 70204
rect 50296 70144 50360 70148
rect 50376 70204 50440 70208
rect 50376 70148 50380 70204
rect 50380 70148 50436 70204
rect 50436 70148 50440 70204
rect 50376 70144 50440 70148
rect 50456 70204 50520 70208
rect 50456 70148 50460 70204
rect 50460 70148 50516 70204
rect 50516 70148 50520 70204
rect 50456 70144 50520 70148
rect 50536 70204 50600 70208
rect 50536 70148 50540 70204
rect 50540 70148 50596 70204
rect 50596 70148 50600 70204
rect 50536 70144 50600 70148
rect 81016 70204 81080 70208
rect 81016 70148 81020 70204
rect 81020 70148 81076 70204
rect 81076 70148 81080 70204
rect 81016 70144 81080 70148
rect 81096 70204 81160 70208
rect 81096 70148 81100 70204
rect 81100 70148 81156 70204
rect 81156 70148 81160 70204
rect 81096 70144 81160 70148
rect 81176 70204 81240 70208
rect 81176 70148 81180 70204
rect 81180 70148 81236 70204
rect 81236 70148 81240 70204
rect 81176 70144 81240 70148
rect 81256 70204 81320 70208
rect 81256 70148 81260 70204
rect 81260 70148 81316 70204
rect 81316 70148 81320 70204
rect 81256 70144 81320 70148
rect 4216 69660 4280 69664
rect 4216 69604 4220 69660
rect 4220 69604 4276 69660
rect 4276 69604 4280 69660
rect 4216 69600 4280 69604
rect 4296 69660 4360 69664
rect 4296 69604 4300 69660
rect 4300 69604 4356 69660
rect 4356 69604 4360 69660
rect 4296 69600 4360 69604
rect 4376 69660 4440 69664
rect 4376 69604 4380 69660
rect 4380 69604 4436 69660
rect 4436 69604 4440 69660
rect 4376 69600 4440 69604
rect 4456 69660 4520 69664
rect 4456 69604 4460 69660
rect 4460 69604 4516 69660
rect 4516 69604 4520 69660
rect 4456 69600 4520 69604
rect 34936 69660 35000 69664
rect 34936 69604 34940 69660
rect 34940 69604 34996 69660
rect 34996 69604 35000 69660
rect 34936 69600 35000 69604
rect 35016 69660 35080 69664
rect 35016 69604 35020 69660
rect 35020 69604 35076 69660
rect 35076 69604 35080 69660
rect 35016 69600 35080 69604
rect 35096 69660 35160 69664
rect 35096 69604 35100 69660
rect 35100 69604 35156 69660
rect 35156 69604 35160 69660
rect 35096 69600 35160 69604
rect 35176 69660 35240 69664
rect 35176 69604 35180 69660
rect 35180 69604 35236 69660
rect 35236 69604 35240 69660
rect 35176 69600 35240 69604
rect 65656 69660 65720 69664
rect 65656 69604 65660 69660
rect 65660 69604 65716 69660
rect 65716 69604 65720 69660
rect 65656 69600 65720 69604
rect 65736 69660 65800 69664
rect 65736 69604 65740 69660
rect 65740 69604 65796 69660
rect 65796 69604 65800 69660
rect 65736 69600 65800 69604
rect 65816 69660 65880 69664
rect 65816 69604 65820 69660
rect 65820 69604 65876 69660
rect 65876 69604 65880 69660
rect 65816 69600 65880 69604
rect 65896 69660 65960 69664
rect 65896 69604 65900 69660
rect 65900 69604 65956 69660
rect 65956 69604 65960 69660
rect 65896 69600 65960 69604
rect 96376 69660 96440 69664
rect 96376 69604 96380 69660
rect 96380 69604 96436 69660
rect 96436 69604 96440 69660
rect 96376 69600 96440 69604
rect 96456 69660 96520 69664
rect 96456 69604 96460 69660
rect 96460 69604 96516 69660
rect 96516 69604 96520 69660
rect 96456 69600 96520 69604
rect 96536 69660 96600 69664
rect 96536 69604 96540 69660
rect 96540 69604 96596 69660
rect 96596 69604 96600 69660
rect 96536 69600 96600 69604
rect 96616 69660 96680 69664
rect 96616 69604 96620 69660
rect 96620 69604 96676 69660
rect 96676 69604 96680 69660
rect 96616 69600 96680 69604
rect 19576 69116 19640 69120
rect 19576 69060 19580 69116
rect 19580 69060 19636 69116
rect 19636 69060 19640 69116
rect 19576 69056 19640 69060
rect 19656 69116 19720 69120
rect 19656 69060 19660 69116
rect 19660 69060 19716 69116
rect 19716 69060 19720 69116
rect 19656 69056 19720 69060
rect 19736 69116 19800 69120
rect 19736 69060 19740 69116
rect 19740 69060 19796 69116
rect 19796 69060 19800 69116
rect 19736 69056 19800 69060
rect 19816 69116 19880 69120
rect 19816 69060 19820 69116
rect 19820 69060 19876 69116
rect 19876 69060 19880 69116
rect 19816 69056 19880 69060
rect 50296 69116 50360 69120
rect 50296 69060 50300 69116
rect 50300 69060 50356 69116
rect 50356 69060 50360 69116
rect 50296 69056 50360 69060
rect 50376 69116 50440 69120
rect 50376 69060 50380 69116
rect 50380 69060 50436 69116
rect 50436 69060 50440 69116
rect 50376 69056 50440 69060
rect 50456 69116 50520 69120
rect 50456 69060 50460 69116
rect 50460 69060 50516 69116
rect 50516 69060 50520 69116
rect 50456 69056 50520 69060
rect 50536 69116 50600 69120
rect 50536 69060 50540 69116
rect 50540 69060 50596 69116
rect 50596 69060 50600 69116
rect 50536 69056 50600 69060
rect 81016 69116 81080 69120
rect 81016 69060 81020 69116
rect 81020 69060 81076 69116
rect 81076 69060 81080 69116
rect 81016 69056 81080 69060
rect 81096 69116 81160 69120
rect 81096 69060 81100 69116
rect 81100 69060 81156 69116
rect 81156 69060 81160 69116
rect 81096 69056 81160 69060
rect 81176 69116 81240 69120
rect 81176 69060 81180 69116
rect 81180 69060 81236 69116
rect 81236 69060 81240 69116
rect 81176 69056 81240 69060
rect 81256 69116 81320 69120
rect 81256 69060 81260 69116
rect 81260 69060 81316 69116
rect 81316 69060 81320 69116
rect 81256 69056 81320 69060
rect 4216 68572 4280 68576
rect 4216 68516 4220 68572
rect 4220 68516 4276 68572
rect 4276 68516 4280 68572
rect 4216 68512 4280 68516
rect 4296 68572 4360 68576
rect 4296 68516 4300 68572
rect 4300 68516 4356 68572
rect 4356 68516 4360 68572
rect 4296 68512 4360 68516
rect 4376 68572 4440 68576
rect 4376 68516 4380 68572
rect 4380 68516 4436 68572
rect 4436 68516 4440 68572
rect 4376 68512 4440 68516
rect 4456 68572 4520 68576
rect 4456 68516 4460 68572
rect 4460 68516 4516 68572
rect 4516 68516 4520 68572
rect 4456 68512 4520 68516
rect 34936 68572 35000 68576
rect 34936 68516 34940 68572
rect 34940 68516 34996 68572
rect 34996 68516 35000 68572
rect 34936 68512 35000 68516
rect 35016 68572 35080 68576
rect 35016 68516 35020 68572
rect 35020 68516 35076 68572
rect 35076 68516 35080 68572
rect 35016 68512 35080 68516
rect 35096 68572 35160 68576
rect 35096 68516 35100 68572
rect 35100 68516 35156 68572
rect 35156 68516 35160 68572
rect 35096 68512 35160 68516
rect 35176 68572 35240 68576
rect 35176 68516 35180 68572
rect 35180 68516 35236 68572
rect 35236 68516 35240 68572
rect 35176 68512 35240 68516
rect 65656 68572 65720 68576
rect 65656 68516 65660 68572
rect 65660 68516 65716 68572
rect 65716 68516 65720 68572
rect 65656 68512 65720 68516
rect 65736 68572 65800 68576
rect 65736 68516 65740 68572
rect 65740 68516 65796 68572
rect 65796 68516 65800 68572
rect 65736 68512 65800 68516
rect 65816 68572 65880 68576
rect 65816 68516 65820 68572
rect 65820 68516 65876 68572
rect 65876 68516 65880 68572
rect 65816 68512 65880 68516
rect 65896 68572 65960 68576
rect 65896 68516 65900 68572
rect 65900 68516 65956 68572
rect 65956 68516 65960 68572
rect 65896 68512 65960 68516
rect 96376 68572 96440 68576
rect 96376 68516 96380 68572
rect 96380 68516 96436 68572
rect 96436 68516 96440 68572
rect 96376 68512 96440 68516
rect 96456 68572 96520 68576
rect 96456 68516 96460 68572
rect 96460 68516 96516 68572
rect 96516 68516 96520 68572
rect 96456 68512 96520 68516
rect 96536 68572 96600 68576
rect 96536 68516 96540 68572
rect 96540 68516 96596 68572
rect 96596 68516 96600 68572
rect 96536 68512 96600 68516
rect 96616 68572 96680 68576
rect 96616 68516 96620 68572
rect 96620 68516 96676 68572
rect 96676 68516 96680 68572
rect 96616 68512 96680 68516
rect 19576 68028 19640 68032
rect 19576 67972 19580 68028
rect 19580 67972 19636 68028
rect 19636 67972 19640 68028
rect 19576 67968 19640 67972
rect 19656 68028 19720 68032
rect 19656 67972 19660 68028
rect 19660 67972 19716 68028
rect 19716 67972 19720 68028
rect 19656 67968 19720 67972
rect 19736 68028 19800 68032
rect 19736 67972 19740 68028
rect 19740 67972 19796 68028
rect 19796 67972 19800 68028
rect 19736 67968 19800 67972
rect 19816 68028 19880 68032
rect 19816 67972 19820 68028
rect 19820 67972 19876 68028
rect 19876 67972 19880 68028
rect 19816 67968 19880 67972
rect 50296 68028 50360 68032
rect 50296 67972 50300 68028
rect 50300 67972 50356 68028
rect 50356 67972 50360 68028
rect 50296 67968 50360 67972
rect 50376 68028 50440 68032
rect 50376 67972 50380 68028
rect 50380 67972 50436 68028
rect 50436 67972 50440 68028
rect 50376 67968 50440 67972
rect 50456 68028 50520 68032
rect 50456 67972 50460 68028
rect 50460 67972 50516 68028
rect 50516 67972 50520 68028
rect 50456 67968 50520 67972
rect 50536 68028 50600 68032
rect 50536 67972 50540 68028
rect 50540 67972 50596 68028
rect 50596 67972 50600 68028
rect 50536 67968 50600 67972
rect 81016 68028 81080 68032
rect 81016 67972 81020 68028
rect 81020 67972 81076 68028
rect 81076 67972 81080 68028
rect 81016 67968 81080 67972
rect 81096 68028 81160 68032
rect 81096 67972 81100 68028
rect 81100 67972 81156 68028
rect 81156 67972 81160 68028
rect 81096 67968 81160 67972
rect 81176 68028 81240 68032
rect 81176 67972 81180 68028
rect 81180 67972 81236 68028
rect 81236 67972 81240 68028
rect 81176 67968 81240 67972
rect 81256 68028 81320 68032
rect 81256 67972 81260 68028
rect 81260 67972 81316 68028
rect 81316 67972 81320 68028
rect 81256 67968 81320 67972
rect 4216 67484 4280 67488
rect 4216 67428 4220 67484
rect 4220 67428 4276 67484
rect 4276 67428 4280 67484
rect 4216 67424 4280 67428
rect 4296 67484 4360 67488
rect 4296 67428 4300 67484
rect 4300 67428 4356 67484
rect 4356 67428 4360 67484
rect 4296 67424 4360 67428
rect 4376 67484 4440 67488
rect 4376 67428 4380 67484
rect 4380 67428 4436 67484
rect 4436 67428 4440 67484
rect 4376 67424 4440 67428
rect 4456 67484 4520 67488
rect 4456 67428 4460 67484
rect 4460 67428 4516 67484
rect 4516 67428 4520 67484
rect 4456 67424 4520 67428
rect 34936 67484 35000 67488
rect 34936 67428 34940 67484
rect 34940 67428 34996 67484
rect 34996 67428 35000 67484
rect 34936 67424 35000 67428
rect 35016 67484 35080 67488
rect 35016 67428 35020 67484
rect 35020 67428 35076 67484
rect 35076 67428 35080 67484
rect 35016 67424 35080 67428
rect 35096 67484 35160 67488
rect 35096 67428 35100 67484
rect 35100 67428 35156 67484
rect 35156 67428 35160 67484
rect 35096 67424 35160 67428
rect 35176 67484 35240 67488
rect 35176 67428 35180 67484
rect 35180 67428 35236 67484
rect 35236 67428 35240 67484
rect 35176 67424 35240 67428
rect 65656 67484 65720 67488
rect 65656 67428 65660 67484
rect 65660 67428 65716 67484
rect 65716 67428 65720 67484
rect 65656 67424 65720 67428
rect 65736 67484 65800 67488
rect 65736 67428 65740 67484
rect 65740 67428 65796 67484
rect 65796 67428 65800 67484
rect 65736 67424 65800 67428
rect 65816 67484 65880 67488
rect 65816 67428 65820 67484
rect 65820 67428 65876 67484
rect 65876 67428 65880 67484
rect 65816 67424 65880 67428
rect 65896 67484 65960 67488
rect 65896 67428 65900 67484
rect 65900 67428 65956 67484
rect 65956 67428 65960 67484
rect 65896 67424 65960 67428
rect 96376 67484 96440 67488
rect 96376 67428 96380 67484
rect 96380 67428 96436 67484
rect 96436 67428 96440 67484
rect 96376 67424 96440 67428
rect 96456 67484 96520 67488
rect 96456 67428 96460 67484
rect 96460 67428 96516 67484
rect 96516 67428 96520 67484
rect 96456 67424 96520 67428
rect 96536 67484 96600 67488
rect 96536 67428 96540 67484
rect 96540 67428 96596 67484
rect 96596 67428 96600 67484
rect 96536 67424 96600 67428
rect 96616 67484 96680 67488
rect 96616 67428 96620 67484
rect 96620 67428 96676 67484
rect 96676 67428 96680 67484
rect 96616 67424 96680 67428
rect 19576 66940 19640 66944
rect 19576 66884 19580 66940
rect 19580 66884 19636 66940
rect 19636 66884 19640 66940
rect 19576 66880 19640 66884
rect 19656 66940 19720 66944
rect 19656 66884 19660 66940
rect 19660 66884 19716 66940
rect 19716 66884 19720 66940
rect 19656 66880 19720 66884
rect 19736 66940 19800 66944
rect 19736 66884 19740 66940
rect 19740 66884 19796 66940
rect 19796 66884 19800 66940
rect 19736 66880 19800 66884
rect 19816 66940 19880 66944
rect 19816 66884 19820 66940
rect 19820 66884 19876 66940
rect 19876 66884 19880 66940
rect 19816 66880 19880 66884
rect 50296 66940 50360 66944
rect 50296 66884 50300 66940
rect 50300 66884 50356 66940
rect 50356 66884 50360 66940
rect 50296 66880 50360 66884
rect 50376 66940 50440 66944
rect 50376 66884 50380 66940
rect 50380 66884 50436 66940
rect 50436 66884 50440 66940
rect 50376 66880 50440 66884
rect 50456 66940 50520 66944
rect 50456 66884 50460 66940
rect 50460 66884 50516 66940
rect 50516 66884 50520 66940
rect 50456 66880 50520 66884
rect 50536 66940 50600 66944
rect 50536 66884 50540 66940
rect 50540 66884 50596 66940
rect 50596 66884 50600 66940
rect 50536 66880 50600 66884
rect 81016 66940 81080 66944
rect 81016 66884 81020 66940
rect 81020 66884 81076 66940
rect 81076 66884 81080 66940
rect 81016 66880 81080 66884
rect 81096 66940 81160 66944
rect 81096 66884 81100 66940
rect 81100 66884 81156 66940
rect 81156 66884 81160 66940
rect 81096 66880 81160 66884
rect 81176 66940 81240 66944
rect 81176 66884 81180 66940
rect 81180 66884 81236 66940
rect 81236 66884 81240 66940
rect 81176 66880 81240 66884
rect 81256 66940 81320 66944
rect 81256 66884 81260 66940
rect 81260 66884 81316 66940
rect 81316 66884 81320 66940
rect 81256 66880 81320 66884
rect 4216 66396 4280 66400
rect 4216 66340 4220 66396
rect 4220 66340 4276 66396
rect 4276 66340 4280 66396
rect 4216 66336 4280 66340
rect 4296 66396 4360 66400
rect 4296 66340 4300 66396
rect 4300 66340 4356 66396
rect 4356 66340 4360 66396
rect 4296 66336 4360 66340
rect 4376 66396 4440 66400
rect 4376 66340 4380 66396
rect 4380 66340 4436 66396
rect 4436 66340 4440 66396
rect 4376 66336 4440 66340
rect 4456 66396 4520 66400
rect 4456 66340 4460 66396
rect 4460 66340 4516 66396
rect 4516 66340 4520 66396
rect 4456 66336 4520 66340
rect 34936 66396 35000 66400
rect 34936 66340 34940 66396
rect 34940 66340 34996 66396
rect 34996 66340 35000 66396
rect 34936 66336 35000 66340
rect 35016 66396 35080 66400
rect 35016 66340 35020 66396
rect 35020 66340 35076 66396
rect 35076 66340 35080 66396
rect 35016 66336 35080 66340
rect 35096 66396 35160 66400
rect 35096 66340 35100 66396
rect 35100 66340 35156 66396
rect 35156 66340 35160 66396
rect 35096 66336 35160 66340
rect 35176 66396 35240 66400
rect 35176 66340 35180 66396
rect 35180 66340 35236 66396
rect 35236 66340 35240 66396
rect 35176 66336 35240 66340
rect 65656 66396 65720 66400
rect 65656 66340 65660 66396
rect 65660 66340 65716 66396
rect 65716 66340 65720 66396
rect 65656 66336 65720 66340
rect 65736 66396 65800 66400
rect 65736 66340 65740 66396
rect 65740 66340 65796 66396
rect 65796 66340 65800 66396
rect 65736 66336 65800 66340
rect 65816 66396 65880 66400
rect 65816 66340 65820 66396
rect 65820 66340 65876 66396
rect 65876 66340 65880 66396
rect 65816 66336 65880 66340
rect 65896 66396 65960 66400
rect 65896 66340 65900 66396
rect 65900 66340 65956 66396
rect 65956 66340 65960 66396
rect 65896 66336 65960 66340
rect 96376 66396 96440 66400
rect 96376 66340 96380 66396
rect 96380 66340 96436 66396
rect 96436 66340 96440 66396
rect 96376 66336 96440 66340
rect 96456 66396 96520 66400
rect 96456 66340 96460 66396
rect 96460 66340 96516 66396
rect 96516 66340 96520 66396
rect 96456 66336 96520 66340
rect 96536 66396 96600 66400
rect 96536 66340 96540 66396
rect 96540 66340 96596 66396
rect 96596 66340 96600 66396
rect 96536 66336 96600 66340
rect 96616 66396 96680 66400
rect 96616 66340 96620 66396
rect 96620 66340 96676 66396
rect 96676 66340 96680 66396
rect 96616 66336 96680 66340
rect 19576 65852 19640 65856
rect 19576 65796 19580 65852
rect 19580 65796 19636 65852
rect 19636 65796 19640 65852
rect 19576 65792 19640 65796
rect 19656 65852 19720 65856
rect 19656 65796 19660 65852
rect 19660 65796 19716 65852
rect 19716 65796 19720 65852
rect 19656 65792 19720 65796
rect 19736 65852 19800 65856
rect 19736 65796 19740 65852
rect 19740 65796 19796 65852
rect 19796 65796 19800 65852
rect 19736 65792 19800 65796
rect 19816 65852 19880 65856
rect 19816 65796 19820 65852
rect 19820 65796 19876 65852
rect 19876 65796 19880 65852
rect 19816 65792 19880 65796
rect 50296 65852 50360 65856
rect 50296 65796 50300 65852
rect 50300 65796 50356 65852
rect 50356 65796 50360 65852
rect 50296 65792 50360 65796
rect 50376 65852 50440 65856
rect 50376 65796 50380 65852
rect 50380 65796 50436 65852
rect 50436 65796 50440 65852
rect 50376 65792 50440 65796
rect 50456 65852 50520 65856
rect 50456 65796 50460 65852
rect 50460 65796 50516 65852
rect 50516 65796 50520 65852
rect 50456 65792 50520 65796
rect 50536 65852 50600 65856
rect 50536 65796 50540 65852
rect 50540 65796 50596 65852
rect 50596 65796 50600 65852
rect 50536 65792 50600 65796
rect 81016 65852 81080 65856
rect 81016 65796 81020 65852
rect 81020 65796 81076 65852
rect 81076 65796 81080 65852
rect 81016 65792 81080 65796
rect 81096 65852 81160 65856
rect 81096 65796 81100 65852
rect 81100 65796 81156 65852
rect 81156 65796 81160 65852
rect 81096 65792 81160 65796
rect 81176 65852 81240 65856
rect 81176 65796 81180 65852
rect 81180 65796 81236 65852
rect 81236 65796 81240 65852
rect 81176 65792 81240 65796
rect 81256 65852 81320 65856
rect 81256 65796 81260 65852
rect 81260 65796 81316 65852
rect 81316 65796 81320 65852
rect 81256 65792 81320 65796
rect 4216 65308 4280 65312
rect 4216 65252 4220 65308
rect 4220 65252 4276 65308
rect 4276 65252 4280 65308
rect 4216 65248 4280 65252
rect 4296 65308 4360 65312
rect 4296 65252 4300 65308
rect 4300 65252 4356 65308
rect 4356 65252 4360 65308
rect 4296 65248 4360 65252
rect 4376 65308 4440 65312
rect 4376 65252 4380 65308
rect 4380 65252 4436 65308
rect 4436 65252 4440 65308
rect 4376 65248 4440 65252
rect 4456 65308 4520 65312
rect 4456 65252 4460 65308
rect 4460 65252 4516 65308
rect 4516 65252 4520 65308
rect 4456 65248 4520 65252
rect 34936 65308 35000 65312
rect 34936 65252 34940 65308
rect 34940 65252 34996 65308
rect 34996 65252 35000 65308
rect 34936 65248 35000 65252
rect 35016 65308 35080 65312
rect 35016 65252 35020 65308
rect 35020 65252 35076 65308
rect 35076 65252 35080 65308
rect 35016 65248 35080 65252
rect 35096 65308 35160 65312
rect 35096 65252 35100 65308
rect 35100 65252 35156 65308
rect 35156 65252 35160 65308
rect 35096 65248 35160 65252
rect 35176 65308 35240 65312
rect 35176 65252 35180 65308
rect 35180 65252 35236 65308
rect 35236 65252 35240 65308
rect 35176 65248 35240 65252
rect 65656 65308 65720 65312
rect 65656 65252 65660 65308
rect 65660 65252 65716 65308
rect 65716 65252 65720 65308
rect 65656 65248 65720 65252
rect 65736 65308 65800 65312
rect 65736 65252 65740 65308
rect 65740 65252 65796 65308
rect 65796 65252 65800 65308
rect 65736 65248 65800 65252
rect 65816 65308 65880 65312
rect 65816 65252 65820 65308
rect 65820 65252 65876 65308
rect 65876 65252 65880 65308
rect 65816 65248 65880 65252
rect 65896 65308 65960 65312
rect 65896 65252 65900 65308
rect 65900 65252 65956 65308
rect 65956 65252 65960 65308
rect 65896 65248 65960 65252
rect 96376 65308 96440 65312
rect 96376 65252 96380 65308
rect 96380 65252 96436 65308
rect 96436 65252 96440 65308
rect 96376 65248 96440 65252
rect 96456 65308 96520 65312
rect 96456 65252 96460 65308
rect 96460 65252 96516 65308
rect 96516 65252 96520 65308
rect 96456 65248 96520 65252
rect 96536 65308 96600 65312
rect 96536 65252 96540 65308
rect 96540 65252 96596 65308
rect 96596 65252 96600 65308
rect 96536 65248 96600 65252
rect 96616 65308 96680 65312
rect 96616 65252 96620 65308
rect 96620 65252 96676 65308
rect 96676 65252 96680 65308
rect 96616 65248 96680 65252
rect 19576 64764 19640 64768
rect 19576 64708 19580 64764
rect 19580 64708 19636 64764
rect 19636 64708 19640 64764
rect 19576 64704 19640 64708
rect 19656 64764 19720 64768
rect 19656 64708 19660 64764
rect 19660 64708 19716 64764
rect 19716 64708 19720 64764
rect 19656 64704 19720 64708
rect 19736 64764 19800 64768
rect 19736 64708 19740 64764
rect 19740 64708 19796 64764
rect 19796 64708 19800 64764
rect 19736 64704 19800 64708
rect 19816 64764 19880 64768
rect 19816 64708 19820 64764
rect 19820 64708 19876 64764
rect 19876 64708 19880 64764
rect 19816 64704 19880 64708
rect 50296 64764 50360 64768
rect 50296 64708 50300 64764
rect 50300 64708 50356 64764
rect 50356 64708 50360 64764
rect 50296 64704 50360 64708
rect 50376 64764 50440 64768
rect 50376 64708 50380 64764
rect 50380 64708 50436 64764
rect 50436 64708 50440 64764
rect 50376 64704 50440 64708
rect 50456 64764 50520 64768
rect 50456 64708 50460 64764
rect 50460 64708 50516 64764
rect 50516 64708 50520 64764
rect 50456 64704 50520 64708
rect 50536 64764 50600 64768
rect 50536 64708 50540 64764
rect 50540 64708 50596 64764
rect 50596 64708 50600 64764
rect 50536 64704 50600 64708
rect 81016 64764 81080 64768
rect 81016 64708 81020 64764
rect 81020 64708 81076 64764
rect 81076 64708 81080 64764
rect 81016 64704 81080 64708
rect 81096 64764 81160 64768
rect 81096 64708 81100 64764
rect 81100 64708 81156 64764
rect 81156 64708 81160 64764
rect 81096 64704 81160 64708
rect 81176 64764 81240 64768
rect 81176 64708 81180 64764
rect 81180 64708 81236 64764
rect 81236 64708 81240 64764
rect 81176 64704 81240 64708
rect 81256 64764 81320 64768
rect 81256 64708 81260 64764
rect 81260 64708 81316 64764
rect 81316 64708 81320 64764
rect 81256 64704 81320 64708
rect 4216 64220 4280 64224
rect 4216 64164 4220 64220
rect 4220 64164 4276 64220
rect 4276 64164 4280 64220
rect 4216 64160 4280 64164
rect 4296 64220 4360 64224
rect 4296 64164 4300 64220
rect 4300 64164 4356 64220
rect 4356 64164 4360 64220
rect 4296 64160 4360 64164
rect 4376 64220 4440 64224
rect 4376 64164 4380 64220
rect 4380 64164 4436 64220
rect 4436 64164 4440 64220
rect 4376 64160 4440 64164
rect 4456 64220 4520 64224
rect 4456 64164 4460 64220
rect 4460 64164 4516 64220
rect 4516 64164 4520 64220
rect 4456 64160 4520 64164
rect 34936 64220 35000 64224
rect 34936 64164 34940 64220
rect 34940 64164 34996 64220
rect 34996 64164 35000 64220
rect 34936 64160 35000 64164
rect 35016 64220 35080 64224
rect 35016 64164 35020 64220
rect 35020 64164 35076 64220
rect 35076 64164 35080 64220
rect 35016 64160 35080 64164
rect 35096 64220 35160 64224
rect 35096 64164 35100 64220
rect 35100 64164 35156 64220
rect 35156 64164 35160 64220
rect 35096 64160 35160 64164
rect 35176 64220 35240 64224
rect 35176 64164 35180 64220
rect 35180 64164 35236 64220
rect 35236 64164 35240 64220
rect 35176 64160 35240 64164
rect 65656 64220 65720 64224
rect 65656 64164 65660 64220
rect 65660 64164 65716 64220
rect 65716 64164 65720 64220
rect 65656 64160 65720 64164
rect 65736 64220 65800 64224
rect 65736 64164 65740 64220
rect 65740 64164 65796 64220
rect 65796 64164 65800 64220
rect 65736 64160 65800 64164
rect 65816 64220 65880 64224
rect 65816 64164 65820 64220
rect 65820 64164 65876 64220
rect 65876 64164 65880 64220
rect 65816 64160 65880 64164
rect 65896 64220 65960 64224
rect 65896 64164 65900 64220
rect 65900 64164 65956 64220
rect 65956 64164 65960 64220
rect 65896 64160 65960 64164
rect 96376 64220 96440 64224
rect 96376 64164 96380 64220
rect 96380 64164 96436 64220
rect 96436 64164 96440 64220
rect 96376 64160 96440 64164
rect 96456 64220 96520 64224
rect 96456 64164 96460 64220
rect 96460 64164 96516 64220
rect 96516 64164 96520 64220
rect 96456 64160 96520 64164
rect 96536 64220 96600 64224
rect 96536 64164 96540 64220
rect 96540 64164 96596 64220
rect 96596 64164 96600 64220
rect 96536 64160 96600 64164
rect 96616 64220 96680 64224
rect 96616 64164 96620 64220
rect 96620 64164 96676 64220
rect 96676 64164 96680 64220
rect 96616 64160 96680 64164
rect 19576 63676 19640 63680
rect 19576 63620 19580 63676
rect 19580 63620 19636 63676
rect 19636 63620 19640 63676
rect 19576 63616 19640 63620
rect 19656 63676 19720 63680
rect 19656 63620 19660 63676
rect 19660 63620 19716 63676
rect 19716 63620 19720 63676
rect 19656 63616 19720 63620
rect 19736 63676 19800 63680
rect 19736 63620 19740 63676
rect 19740 63620 19796 63676
rect 19796 63620 19800 63676
rect 19736 63616 19800 63620
rect 19816 63676 19880 63680
rect 19816 63620 19820 63676
rect 19820 63620 19876 63676
rect 19876 63620 19880 63676
rect 19816 63616 19880 63620
rect 50296 63676 50360 63680
rect 50296 63620 50300 63676
rect 50300 63620 50356 63676
rect 50356 63620 50360 63676
rect 50296 63616 50360 63620
rect 50376 63676 50440 63680
rect 50376 63620 50380 63676
rect 50380 63620 50436 63676
rect 50436 63620 50440 63676
rect 50376 63616 50440 63620
rect 50456 63676 50520 63680
rect 50456 63620 50460 63676
rect 50460 63620 50516 63676
rect 50516 63620 50520 63676
rect 50456 63616 50520 63620
rect 50536 63676 50600 63680
rect 50536 63620 50540 63676
rect 50540 63620 50596 63676
rect 50596 63620 50600 63676
rect 50536 63616 50600 63620
rect 81016 63676 81080 63680
rect 81016 63620 81020 63676
rect 81020 63620 81076 63676
rect 81076 63620 81080 63676
rect 81016 63616 81080 63620
rect 81096 63676 81160 63680
rect 81096 63620 81100 63676
rect 81100 63620 81156 63676
rect 81156 63620 81160 63676
rect 81096 63616 81160 63620
rect 81176 63676 81240 63680
rect 81176 63620 81180 63676
rect 81180 63620 81236 63676
rect 81236 63620 81240 63676
rect 81176 63616 81240 63620
rect 81256 63676 81320 63680
rect 81256 63620 81260 63676
rect 81260 63620 81316 63676
rect 81316 63620 81320 63676
rect 81256 63616 81320 63620
rect 4216 63132 4280 63136
rect 4216 63076 4220 63132
rect 4220 63076 4276 63132
rect 4276 63076 4280 63132
rect 4216 63072 4280 63076
rect 4296 63132 4360 63136
rect 4296 63076 4300 63132
rect 4300 63076 4356 63132
rect 4356 63076 4360 63132
rect 4296 63072 4360 63076
rect 4376 63132 4440 63136
rect 4376 63076 4380 63132
rect 4380 63076 4436 63132
rect 4436 63076 4440 63132
rect 4376 63072 4440 63076
rect 4456 63132 4520 63136
rect 4456 63076 4460 63132
rect 4460 63076 4516 63132
rect 4516 63076 4520 63132
rect 4456 63072 4520 63076
rect 34936 63132 35000 63136
rect 34936 63076 34940 63132
rect 34940 63076 34996 63132
rect 34996 63076 35000 63132
rect 34936 63072 35000 63076
rect 35016 63132 35080 63136
rect 35016 63076 35020 63132
rect 35020 63076 35076 63132
rect 35076 63076 35080 63132
rect 35016 63072 35080 63076
rect 35096 63132 35160 63136
rect 35096 63076 35100 63132
rect 35100 63076 35156 63132
rect 35156 63076 35160 63132
rect 35096 63072 35160 63076
rect 35176 63132 35240 63136
rect 35176 63076 35180 63132
rect 35180 63076 35236 63132
rect 35236 63076 35240 63132
rect 35176 63072 35240 63076
rect 65656 63132 65720 63136
rect 65656 63076 65660 63132
rect 65660 63076 65716 63132
rect 65716 63076 65720 63132
rect 65656 63072 65720 63076
rect 65736 63132 65800 63136
rect 65736 63076 65740 63132
rect 65740 63076 65796 63132
rect 65796 63076 65800 63132
rect 65736 63072 65800 63076
rect 65816 63132 65880 63136
rect 65816 63076 65820 63132
rect 65820 63076 65876 63132
rect 65876 63076 65880 63132
rect 65816 63072 65880 63076
rect 65896 63132 65960 63136
rect 65896 63076 65900 63132
rect 65900 63076 65956 63132
rect 65956 63076 65960 63132
rect 65896 63072 65960 63076
rect 96376 63132 96440 63136
rect 96376 63076 96380 63132
rect 96380 63076 96436 63132
rect 96436 63076 96440 63132
rect 96376 63072 96440 63076
rect 96456 63132 96520 63136
rect 96456 63076 96460 63132
rect 96460 63076 96516 63132
rect 96516 63076 96520 63132
rect 96456 63072 96520 63076
rect 96536 63132 96600 63136
rect 96536 63076 96540 63132
rect 96540 63076 96596 63132
rect 96596 63076 96600 63132
rect 96536 63072 96600 63076
rect 96616 63132 96680 63136
rect 96616 63076 96620 63132
rect 96620 63076 96676 63132
rect 96676 63076 96680 63132
rect 96616 63072 96680 63076
rect 19576 62588 19640 62592
rect 19576 62532 19580 62588
rect 19580 62532 19636 62588
rect 19636 62532 19640 62588
rect 19576 62528 19640 62532
rect 19656 62588 19720 62592
rect 19656 62532 19660 62588
rect 19660 62532 19716 62588
rect 19716 62532 19720 62588
rect 19656 62528 19720 62532
rect 19736 62588 19800 62592
rect 19736 62532 19740 62588
rect 19740 62532 19796 62588
rect 19796 62532 19800 62588
rect 19736 62528 19800 62532
rect 19816 62588 19880 62592
rect 19816 62532 19820 62588
rect 19820 62532 19876 62588
rect 19876 62532 19880 62588
rect 19816 62528 19880 62532
rect 50296 62588 50360 62592
rect 50296 62532 50300 62588
rect 50300 62532 50356 62588
rect 50356 62532 50360 62588
rect 50296 62528 50360 62532
rect 50376 62588 50440 62592
rect 50376 62532 50380 62588
rect 50380 62532 50436 62588
rect 50436 62532 50440 62588
rect 50376 62528 50440 62532
rect 50456 62588 50520 62592
rect 50456 62532 50460 62588
rect 50460 62532 50516 62588
rect 50516 62532 50520 62588
rect 50456 62528 50520 62532
rect 50536 62588 50600 62592
rect 50536 62532 50540 62588
rect 50540 62532 50596 62588
rect 50596 62532 50600 62588
rect 50536 62528 50600 62532
rect 81016 62588 81080 62592
rect 81016 62532 81020 62588
rect 81020 62532 81076 62588
rect 81076 62532 81080 62588
rect 81016 62528 81080 62532
rect 81096 62588 81160 62592
rect 81096 62532 81100 62588
rect 81100 62532 81156 62588
rect 81156 62532 81160 62588
rect 81096 62528 81160 62532
rect 81176 62588 81240 62592
rect 81176 62532 81180 62588
rect 81180 62532 81236 62588
rect 81236 62532 81240 62588
rect 81176 62528 81240 62532
rect 81256 62588 81320 62592
rect 81256 62532 81260 62588
rect 81260 62532 81316 62588
rect 81316 62532 81320 62588
rect 81256 62528 81320 62532
rect 4216 62044 4280 62048
rect 4216 61988 4220 62044
rect 4220 61988 4276 62044
rect 4276 61988 4280 62044
rect 4216 61984 4280 61988
rect 4296 62044 4360 62048
rect 4296 61988 4300 62044
rect 4300 61988 4356 62044
rect 4356 61988 4360 62044
rect 4296 61984 4360 61988
rect 4376 62044 4440 62048
rect 4376 61988 4380 62044
rect 4380 61988 4436 62044
rect 4436 61988 4440 62044
rect 4376 61984 4440 61988
rect 4456 62044 4520 62048
rect 4456 61988 4460 62044
rect 4460 61988 4516 62044
rect 4516 61988 4520 62044
rect 4456 61984 4520 61988
rect 34936 62044 35000 62048
rect 34936 61988 34940 62044
rect 34940 61988 34996 62044
rect 34996 61988 35000 62044
rect 34936 61984 35000 61988
rect 35016 62044 35080 62048
rect 35016 61988 35020 62044
rect 35020 61988 35076 62044
rect 35076 61988 35080 62044
rect 35016 61984 35080 61988
rect 35096 62044 35160 62048
rect 35096 61988 35100 62044
rect 35100 61988 35156 62044
rect 35156 61988 35160 62044
rect 35096 61984 35160 61988
rect 35176 62044 35240 62048
rect 35176 61988 35180 62044
rect 35180 61988 35236 62044
rect 35236 61988 35240 62044
rect 35176 61984 35240 61988
rect 65656 62044 65720 62048
rect 65656 61988 65660 62044
rect 65660 61988 65716 62044
rect 65716 61988 65720 62044
rect 65656 61984 65720 61988
rect 65736 62044 65800 62048
rect 65736 61988 65740 62044
rect 65740 61988 65796 62044
rect 65796 61988 65800 62044
rect 65736 61984 65800 61988
rect 65816 62044 65880 62048
rect 65816 61988 65820 62044
rect 65820 61988 65876 62044
rect 65876 61988 65880 62044
rect 65816 61984 65880 61988
rect 65896 62044 65960 62048
rect 65896 61988 65900 62044
rect 65900 61988 65956 62044
rect 65956 61988 65960 62044
rect 65896 61984 65960 61988
rect 96376 62044 96440 62048
rect 96376 61988 96380 62044
rect 96380 61988 96436 62044
rect 96436 61988 96440 62044
rect 96376 61984 96440 61988
rect 96456 62044 96520 62048
rect 96456 61988 96460 62044
rect 96460 61988 96516 62044
rect 96516 61988 96520 62044
rect 96456 61984 96520 61988
rect 96536 62044 96600 62048
rect 96536 61988 96540 62044
rect 96540 61988 96596 62044
rect 96596 61988 96600 62044
rect 96536 61984 96600 61988
rect 96616 62044 96680 62048
rect 96616 61988 96620 62044
rect 96620 61988 96676 62044
rect 96676 61988 96680 62044
rect 96616 61984 96680 61988
rect 19576 61500 19640 61504
rect 19576 61444 19580 61500
rect 19580 61444 19636 61500
rect 19636 61444 19640 61500
rect 19576 61440 19640 61444
rect 19656 61500 19720 61504
rect 19656 61444 19660 61500
rect 19660 61444 19716 61500
rect 19716 61444 19720 61500
rect 19656 61440 19720 61444
rect 19736 61500 19800 61504
rect 19736 61444 19740 61500
rect 19740 61444 19796 61500
rect 19796 61444 19800 61500
rect 19736 61440 19800 61444
rect 19816 61500 19880 61504
rect 19816 61444 19820 61500
rect 19820 61444 19876 61500
rect 19876 61444 19880 61500
rect 19816 61440 19880 61444
rect 50296 61500 50360 61504
rect 50296 61444 50300 61500
rect 50300 61444 50356 61500
rect 50356 61444 50360 61500
rect 50296 61440 50360 61444
rect 50376 61500 50440 61504
rect 50376 61444 50380 61500
rect 50380 61444 50436 61500
rect 50436 61444 50440 61500
rect 50376 61440 50440 61444
rect 50456 61500 50520 61504
rect 50456 61444 50460 61500
rect 50460 61444 50516 61500
rect 50516 61444 50520 61500
rect 50456 61440 50520 61444
rect 50536 61500 50600 61504
rect 50536 61444 50540 61500
rect 50540 61444 50596 61500
rect 50596 61444 50600 61500
rect 50536 61440 50600 61444
rect 81016 61500 81080 61504
rect 81016 61444 81020 61500
rect 81020 61444 81076 61500
rect 81076 61444 81080 61500
rect 81016 61440 81080 61444
rect 81096 61500 81160 61504
rect 81096 61444 81100 61500
rect 81100 61444 81156 61500
rect 81156 61444 81160 61500
rect 81096 61440 81160 61444
rect 81176 61500 81240 61504
rect 81176 61444 81180 61500
rect 81180 61444 81236 61500
rect 81236 61444 81240 61500
rect 81176 61440 81240 61444
rect 81256 61500 81320 61504
rect 81256 61444 81260 61500
rect 81260 61444 81316 61500
rect 81316 61444 81320 61500
rect 81256 61440 81320 61444
rect 4216 60956 4280 60960
rect 4216 60900 4220 60956
rect 4220 60900 4276 60956
rect 4276 60900 4280 60956
rect 4216 60896 4280 60900
rect 4296 60956 4360 60960
rect 4296 60900 4300 60956
rect 4300 60900 4356 60956
rect 4356 60900 4360 60956
rect 4296 60896 4360 60900
rect 4376 60956 4440 60960
rect 4376 60900 4380 60956
rect 4380 60900 4436 60956
rect 4436 60900 4440 60956
rect 4376 60896 4440 60900
rect 4456 60956 4520 60960
rect 4456 60900 4460 60956
rect 4460 60900 4516 60956
rect 4516 60900 4520 60956
rect 4456 60896 4520 60900
rect 34936 60956 35000 60960
rect 34936 60900 34940 60956
rect 34940 60900 34996 60956
rect 34996 60900 35000 60956
rect 34936 60896 35000 60900
rect 35016 60956 35080 60960
rect 35016 60900 35020 60956
rect 35020 60900 35076 60956
rect 35076 60900 35080 60956
rect 35016 60896 35080 60900
rect 35096 60956 35160 60960
rect 35096 60900 35100 60956
rect 35100 60900 35156 60956
rect 35156 60900 35160 60956
rect 35096 60896 35160 60900
rect 35176 60956 35240 60960
rect 35176 60900 35180 60956
rect 35180 60900 35236 60956
rect 35236 60900 35240 60956
rect 35176 60896 35240 60900
rect 65656 60956 65720 60960
rect 65656 60900 65660 60956
rect 65660 60900 65716 60956
rect 65716 60900 65720 60956
rect 65656 60896 65720 60900
rect 65736 60956 65800 60960
rect 65736 60900 65740 60956
rect 65740 60900 65796 60956
rect 65796 60900 65800 60956
rect 65736 60896 65800 60900
rect 65816 60956 65880 60960
rect 65816 60900 65820 60956
rect 65820 60900 65876 60956
rect 65876 60900 65880 60956
rect 65816 60896 65880 60900
rect 65896 60956 65960 60960
rect 65896 60900 65900 60956
rect 65900 60900 65956 60956
rect 65956 60900 65960 60956
rect 65896 60896 65960 60900
rect 96376 60956 96440 60960
rect 96376 60900 96380 60956
rect 96380 60900 96436 60956
rect 96436 60900 96440 60956
rect 96376 60896 96440 60900
rect 96456 60956 96520 60960
rect 96456 60900 96460 60956
rect 96460 60900 96516 60956
rect 96516 60900 96520 60956
rect 96456 60896 96520 60900
rect 96536 60956 96600 60960
rect 96536 60900 96540 60956
rect 96540 60900 96596 60956
rect 96596 60900 96600 60956
rect 96536 60896 96600 60900
rect 96616 60956 96680 60960
rect 96616 60900 96620 60956
rect 96620 60900 96676 60956
rect 96676 60900 96680 60956
rect 96616 60896 96680 60900
rect 19576 60412 19640 60416
rect 19576 60356 19580 60412
rect 19580 60356 19636 60412
rect 19636 60356 19640 60412
rect 19576 60352 19640 60356
rect 19656 60412 19720 60416
rect 19656 60356 19660 60412
rect 19660 60356 19716 60412
rect 19716 60356 19720 60412
rect 19656 60352 19720 60356
rect 19736 60412 19800 60416
rect 19736 60356 19740 60412
rect 19740 60356 19796 60412
rect 19796 60356 19800 60412
rect 19736 60352 19800 60356
rect 19816 60412 19880 60416
rect 19816 60356 19820 60412
rect 19820 60356 19876 60412
rect 19876 60356 19880 60412
rect 19816 60352 19880 60356
rect 50296 60412 50360 60416
rect 50296 60356 50300 60412
rect 50300 60356 50356 60412
rect 50356 60356 50360 60412
rect 50296 60352 50360 60356
rect 50376 60412 50440 60416
rect 50376 60356 50380 60412
rect 50380 60356 50436 60412
rect 50436 60356 50440 60412
rect 50376 60352 50440 60356
rect 50456 60412 50520 60416
rect 50456 60356 50460 60412
rect 50460 60356 50516 60412
rect 50516 60356 50520 60412
rect 50456 60352 50520 60356
rect 50536 60412 50600 60416
rect 50536 60356 50540 60412
rect 50540 60356 50596 60412
rect 50596 60356 50600 60412
rect 50536 60352 50600 60356
rect 81016 60412 81080 60416
rect 81016 60356 81020 60412
rect 81020 60356 81076 60412
rect 81076 60356 81080 60412
rect 81016 60352 81080 60356
rect 81096 60412 81160 60416
rect 81096 60356 81100 60412
rect 81100 60356 81156 60412
rect 81156 60356 81160 60412
rect 81096 60352 81160 60356
rect 81176 60412 81240 60416
rect 81176 60356 81180 60412
rect 81180 60356 81236 60412
rect 81236 60356 81240 60412
rect 81176 60352 81240 60356
rect 81256 60412 81320 60416
rect 81256 60356 81260 60412
rect 81260 60356 81316 60412
rect 81316 60356 81320 60412
rect 81256 60352 81320 60356
rect 4216 59868 4280 59872
rect 4216 59812 4220 59868
rect 4220 59812 4276 59868
rect 4276 59812 4280 59868
rect 4216 59808 4280 59812
rect 4296 59868 4360 59872
rect 4296 59812 4300 59868
rect 4300 59812 4356 59868
rect 4356 59812 4360 59868
rect 4296 59808 4360 59812
rect 4376 59868 4440 59872
rect 4376 59812 4380 59868
rect 4380 59812 4436 59868
rect 4436 59812 4440 59868
rect 4376 59808 4440 59812
rect 4456 59868 4520 59872
rect 4456 59812 4460 59868
rect 4460 59812 4516 59868
rect 4516 59812 4520 59868
rect 4456 59808 4520 59812
rect 34936 59868 35000 59872
rect 34936 59812 34940 59868
rect 34940 59812 34996 59868
rect 34996 59812 35000 59868
rect 34936 59808 35000 59812
rect 35016 59868 35080 59872
rect 35016 59812 35020 59868
rect 35020 59812 35076 59868
rect 35076 59812 35080 59868
rect 35016 59808 35080 59812
rect 35096 59868 35160 59872
rect 35096 59812 35100 59868
rect 35100 59812 35156 59868
rect 35156 59812 35160 59868
rect 35096 59808 35160 59812
rect 35176 59868 35240 59872
rect 35176 59812 35180 59868
rect 35180 59812 35236 59868
rect 35236 59812 35240 59868
rect 35176 59808 35240 59812
rect 65656 59868 65720 59872
rect 65656 59812 65660 59868
rect 65660 59812 65716 59868
rect 65716 59812 65720 59868
rect 65656 59808 65720 59812
rect 65736 59868 65800 59872
rect 65736 59812 65740 59868
rect 65740 59812 65796 59868
rect 65796 59812 65800 59868
rect 65736 59808 65800 59812
rect 65816 59868 65880 59872
rect 65816 59812 65820 59868
rect 65820 59812 65876 59868
rect 65876 59812 65880 59868
rect 65816 59808 65880 59812
rect 65896 59868 65960 59872
rect 65896 59812 65900 59868
rect 65900 59812 65956 59868
rect 65956 59812 65960 59868
rect 65896 59808 65960 59812
rect 96376 59868 96440 59872
rect 96376 59812 96380 59868
rect 96380 59812 96436 59868
rect 96436 59812 96440 59868
rect 96376 59808 96440 59812
rect 96456 59868 96520 59872
rect 96456 59812 96460 59868
rect 96460 59812 96516 59868
rect 96516 59812 96520 59868
rect 96456 59808 96520 59812
rect 96536 59868 96600 59872
rect 96536 59812 96540 59868
rect 96540 59812 96596 59868
rect 96596 59812 96600 59868
rect 96536 59808 96600 59812
rect 96616 59868 96680 59872
rect 96616 59812 96620 59868
rect 96620 59812 96676 59868
rect 96676 59812 96680 59868
rect 96616 59808 96680 59812
rect 19576 59324 19640 59328
rect 19576 59268 19580 59324
rect 19580 59268 19636 59324
rect 19636 59268 19640 59324
rect 19576 59264 19640 59268
rect 19656 59324 19720 59328
rect 19656 59268 19660 59324
rect 19660 59268 19716 59324
rect 19716 59268 19720 59324
rect 19656 59264 19720 59268
rect 19736 59324 19800 59328
rect 19736 59268 19740 59324
rect 19740 59268 19796 59324
rect 19796 59268 19800 59324
rect 19736 59264 19800 59268
rect 19816 59324 19880 59328
rect 19816 59268 19820 59324
rect 19820 59268 19876 59324
rect 19876 59268 19880 59324
rect 19816 59264 19880 59268
rect 50296 59324 50360 59328
rect 50296 59268 50300 59324
rect 50300 59268 50356 59324
rect 50356 59268 50360 59324
rect 50296 59264 50360 59268
rect 50376 59324 50440 59328
rect 50376 59268 50380 59324
rect 50380 59268 50436 59324
rect 50436 59268 50440 59324
rect 50376 59264 50440 59268
rect 50456 59324 50520 59328
rect 50456 59268 50460 59324
rect 50460 59268 50516 59324
rect 50516 59268 50520 59324
rect 50456 59264 50520 59268
rect 50536 59324 50600 59328
rect 50536 59268 50540 59324
rect 50540 59268 50596 59324
rect 50596 59268 50600 59324
rect 50536 59264 50600 59268
rect 81016 59324 81080 59328
rect 81016 59268 81020 59324
rect 81020 59268 81076 59324
rect 81076 59268 81080 59324
rect 81016 59264 81080 59268
rect 81096 59324 81160 59328
rect 81096 59268 81100 59324
rect 81100 59268 81156 59324
rect 81156 59268 81160 59324
rect 81096 59264 81160 59268
rect 81176 59324 81240 59328
rect 81176 59268 81180 59324
rect 81180 59268 81236 59324
rect 81236 59268 81240 59324
rect 81176 59264 81240 59268
rect 81256 59324 81320 59328
rect 81256 59268 81260 59324
rect 81260 59268 81316 59324
rect 81316 59268 81320 59324
rect 81256 59264 81320 59268
rect 4216 58780 4280 58784
rect 4216 58724 4220 58780
rect 4220 58724 4276 58780
rect 4276 58724 4280 58780
rect 4216 58720 4280 58724
rect 4296 58780 4360 58784
rect 4296 58724 4300 58780
rect 4300 58724 4356 58780
rect 4356 58724 4360 58780
rect 4296 58720 4360 58724
rect 4376 58780 4440 58784
rect 4376 58724 4380 58780
rect 4380 58724 4436 58780
rect 4436 58724 4440 58780
rect 4376 58720 4440 58724
rect 4456 58780 4520 58784
rect 4456 58724 4460 58780
rect 4460 58724 4516 58780
rect 4516 58724 4520 58780
rect 4456 58720 4520 58724
rect 34936 58780 35000 58784
rect 34936 58724 34940 58780
rect 34940 58724 34996 58780
rect 34996 58724 35000 58780
rect 34936 58720 35000 58724
rect 35016 58780 35080 58784
rect 35016 58724 35020 58780
rect 35020 58724 35076 58780
rect 35076 58724 35080 58780
rect 35016 58720 35080 58724
rect 35096 58780 35160 58784
rect 35096 58724 35100 58780
rect 35100 58724 35156 58780
rect 35156 58724 35160 58780
rect 35096 58720 35160 58724
rect 35176 58780 35240 58784
rect 35176 58724 35180 58780
rect 35180 58724 35236 58780
rect 35236 58724 35240 58780
rect 35176 58720 35240 58724
rect 65656 58780 65720 58784
rect 65656 58724 65660 58780
rect 65660 58724 65716 58780
rect 65716 58724 65720 58780
rect 65656 58720 65720 58724
rect 65736 58780 65800 58784
rect 65736 58724 65740 58780
rect 65740 58724 65796 58780
rect 65796 58724 65800 58780
rect 65736 58720 65800 58724
rect 65816 58780 65880 58784
rect 65816 58724 65820 58780
rect 65820 58724 65876 58780
rect 65876 58724 65880 58780
rect 65816 58720 65880 58724
rect 65896 58780 65960 58784
rect 65896 58724 65900 58780
rect 65900 58724 65956 58780
rect 65956 58724 65960 58780
rect 65896 58720 65960 58724
rect 96376 58780 96440 58784
rect 96376 58724 96380 58780
rect 96380 58724 96436 58780
rect 96436 58724 96440 58780
rect 96376 58720 96440 58724
rect 96456 58780 96520 58784
rect 96456 58724 96460 58780
rect 96460 58724 96516 58780
rect 96516 58724 96520 58780
rect 96456 58720 96520 58724
rect 96536 58780 96600 58784
rect 96536 58724 96540 58780
rect 96540 58724 96596 58780
rect 96596 58724 96600 58780
rect 96536 58720 96600 58724
rect 96616 58780 96680 58784
rect 96616 58724 96620 58780
rect 96620 58724 96676 58780
rect 96676 58724 96680 58780
rect 96616 58720 96680 58724
rect 19576 58236 19640 58240
rect 19576 58180 19580 58236
rect 19580 58180 19636 58236
rect 19636 58180 19640 58236
rect 19576 58176 19640 58180
rect 19656 58236 19720 58240
rect 19656 58180 19660 58236
rect 19660 58180 19716 58236
rect 19716 58180 19720 58236
rect 19656 58176 19720 58180
rect 19736 58236 19800 58240
rect 19736 58180 19740 58236
rect 19740 58180 19796 58236
rect 19796 58180 19800 58236
rect 19736 58176 19800 58180
rect 19816 58236 19880 58240
rect 19816 58180 19820 58236
rect 19820 58180 19876 58236
rect 19876 58180 19880 58236
rect 19816 58176 19880 58180
rect 50296 58236 50360 58240
rect 50296 58180 50300 58236
rect 50300 58180 50356 58236
rect 50356 58180 50360 58236
rect 50296 58176 50360 58180
rect 50376 58236 50440 58240
rect 50376 58180 50380 58236
rect 50380 58180 50436 58236
rect 50436 58180 50440 58236
rect 50376 58176 50440 58180
rect 50456 58236 50520 58240
rect 50456 58180 50460 58236
rect 50460 58180 50516 58236
rect 50516 58180 50520 58236
rect 50456 58176 50520 58180
rect 50536 58236 50600 58240
rect 50536 58180 50540 58236
rect 50540 58180 50596 58236
rect 50596 58180 50600 58236
rect 50536 58176 50600 58180
rect 81016 58236 81080 58240
rect 81016 58180 81020 58236
rect 81020 58180 81076 58236
rect 81076 58180 81080 58236
rect 81016 58176 81080 58180
rect 81096 58236 81160 58240
rect 81096 58180 81100 58236
rect 81100 58180 81156 58236
rect 81156 58180 81160 58236
rect 81096 58176 81160 58180
rect 81176 58236 81240 58240
rect 81176 58180 81180 58236
rect 81180 58180 81236 58236
rect 81236 58180 81240 58236
rect 81176 58176 81240 58180
rect 81256 58236 81320 58240
rect 81256 58180 81260 58236
rect 81260 58180 81316 58236
rect 81316 58180 81320 58236
rect 81256 58176 81320 58180
rect 4216 57692 4280 57696
rect 4216 57636 4220 57692
rect 4220 57636 4276 57692
rect 4276 57636 4280 57692
rect 4216 57632 4280 57636
rect 4296 57692 4360 57696
rect 4296 57636 4300 57692
rect 4300 57636 4356 57692
rect 4356 57636 4360 57692
rect 4296 57632 4360 57636
rect 4376 57692 4440 57696
rect 4376 57636 4380 57692
rect 4380 57636 4436 57692
rect 4436 57636 4440 57692
rect 4376 57632 4440 57636
rect 4456 57692 4520 57696
rect 4456 57636 4460 57692
rect 4460 57636 4516 57692
rect 4516 57636 4520 57692
rect 4456 57632 4520 57636
rect 34936 57692 35000 57696
rect 34936 57636 34940 57692
rect 34940 57636 34996 57692
rect 34996 57636 35000 57692
rect 34936 57632 35000 57636
rect 35016 57692 35080 57696
rect 35016 57636 35020 57692
rect 35020 57636 35076 57692
rect 35076 57636 35080 57692
rect 35016 57632 35080 57636
rect 35096 57692 35160 57696
rect 35096 57636 35100 57692
rect 35100 57636 35156 57692
rect 35156 57636 35160 57692
rect 35096 57632 35160 57636
rect 35176 57692 35240 57696
rect 35176 57636 35180 57692
rect 35180 57636 35236 57692
rect 35236 57636 35240 57692
rect 35176 57632 35240 57636
rect 65656 57692 65720 57696
rect 65656 57636 65660 57692
rect 65660 57636 65716 57692
rect 65716 57636 65720 57692
rect 65656 57632 65720 57636
rect 65736 57692 65800 57696
rect 65736 57636 65740 57692
rect 65740 57636 65796 57692
rect 65796 57636 65800 57692
rect 65736 57632 65800 57636
rect 65816 57692 65880 57696
rect 65816 57636 65820 57692
rect 65820 57636 65876 57692
rect 65876 57636 65880 57692
rect 65816 57632 65880 57636
rect 65896 57692 65960 57696
rect 65896 57636 65900 57692
rect 65900 57636 65956 57692
rect 65956 57636 65960 57692
rect 65896 57632 65960 57636
rect 96376 57692 96440 57696
rect 96376 57636 96380 57692
rect 96380 57636 96436 57692
rect 96436 57636 96440 57692
rect 96376 57632 96440 57636
rect 96456 57692 96520 57696
rect 96456 57636 96460 57692
rect 96460 57636 96516 57692
rect 96516 57636 96520 57692
rect 96456 57632 96520 57636
rect 96536 57692 96600 57696
rect 96536 57636 96540 57692
rect 96540 57636 96596 57692
rect 96596 57636 96600 57692
rect 96536 57632 96600 57636
rect 96616 57692 96680 57696
rect 96616 57636 96620 57692
rect 96620 57636 96676 57692
rect 96676 57636 96680 57692
rect 96616 57632 96680 57636
rect 19576 57148 19640 57152
rect 19576 57092 19580 57148
rect 19580 57092 19636 57148
rect 19636 57092 19640 57148
rect 19576 57088 19640 57092
rect 19656 57148 19720 57152
rect 19656 57092 19660 57148
rect 19660 57092 19716 57148
rect 19716 57092 19720 57148
rect 19656 57088 19720 57092
rect 19736 57148 19800 57152
rect 19736 57092 19740 57148
rect 19740 57092 19796 57148
rect 19796 57092 19800 57148
rect 19736 57088 19800 57092
rect 19816 57148 19880 57152
rect 19816 57092 19820 57148
rect 19820 57092 19876 57148
rect 19876 57092 19880 57148
rect 19816 57088 19880 57092
rect 50296 57148 50360 57152
rect 50296 57092 50300 57148
rect 50300 57092 50356 57148
rect 50356 57092 50360 57148
rect 50296 57088 50360 57092
rect 50376 57148 50440 57152
rect 50376 57092 50380 57148
rect 50380 57092 50436 57148
rect 50436 57092 50440 57148
rect 50376 57088 50440 57092
rect 50456 57148 50520 57152
rect 50456 57092 50460 57148
rect 50460 57092 50516 57148
rect 50516 57092 50520 57148
rect 50456 57088 50520 57092
rect 50536 57148 50600 57152
rect 50536 57092 50540 57148
rect 50540 57092 50596 57148
rect 50596 57092 50600 57148
rect 50536 57088 50600 57092
rect 81016 57148 81080 57152
rect 81016 57092 81020 57148
rect 81020 57092 81076 57148
rect 81076 57092 81080 57148
rect 81016 57088 81080 57092
rect 81096 57148 81160 57152
rect 81096 57092 81100 57148
rect 81100 57092 81156 57148
rect 81156 57092 81160 57148
rect 81096 57088 81160 57092
rect 81176 57148 81240 57152
rect 81176 57092 81180 57148
rect 81180 57092 81236 57148
rect 81236 57092 81240 57148
rect 81176 57088 81240 57092
rect 81256 57148 81320 57152
rect 81256 57092 81260 57148
rect 81260 57092 81316 57148
rect 81316 57092 81320 57148
rect 81256 57088 81320 57092
rect 4216 56604 4280 56608
rect 4216 56548 4220 56604
rect 4220 56548 4276 56604
rect 4276 56548 4280 56604
rect 4216 56544 4280 56548
rect 4296 56604 4360 56608
rect 4296 56548 4300 56604
rect 4300 56548 4356 56604
rect 4356 56548 4360 56604
rect 4296 56544 4360 56548
rect 4376 56604 4440 56608
rect 4376 56548 4380 56604
rect 4380 56548 4436 56604
rect 4436 56548 4440 56604
rect 4376 56544 4440 56548
rect 4456 56604 4520 56608
rect 4456 56548 4460 56604
rect 4460 56548 4516 56604
rect 4516 56548 4520 56604
rect 4456 56544 4520 56548
rect 34936 56604 35000 56608
rect 34936 56548 34940 56604
rect 34940 56548 34996 56604
rect 34996 56548 35000 56604
rect 34936 56544 35000 56548
rect 35016 56604 35080 56608
rect 35016 56548 35020 56604
rect 35020 56548 35076 56604
rect 35076 56548 35080 56604
rect 35016 56544 35080 56548
rect 35096 56604 35160 56608
rect 35096 56548 35100 56604
rect 35100 56548 35156 56604
rect 35156 56548 35160 56604
rect 35096 56544 35160 56548
rect 35176 56604 35240 56608
rect 35176 56548 35180 56604
rect 35180 56548 35236 56604
rect 35236 56548 35240 56604
rect 35176 56544 35240 56548
rect 65656 56604 65720 56608
rect 65656 56548 65660 56604
rect 65660 56548 65716 56604
rect 65716 56548 65720 56604
rect 65656 56544 65720 56548
rect 65736 56604 65800 56608
rect 65736 56548 65740 56604
rect 65740 56548 65796 56604
rect 65796 56548 65800 56604
rect 65736 56544 65800 56548
rect 65816 56604 65880 56608
rect 65816 56548 65820 56604
rect 65820 56548 65876 56604
rect 65876 56548 65880 56604
rect 65816 56544 65880 56548
rect 65896 56604 65960 56608
rect 65896 56548 65900 56604
rect 65900 56548 65956 56604
rect 65956 56548 65960 56604
rect 65896 56544 65960 56548
rect 96376 56604 96440 56608
rect 96376 56548 96380 56604
rect 96380 56548 96436 56604
rect 96436 56548 96440 56604
rect 96376 56544 96440 56548
rect 96456 56604 96520 56608
rect 96456 56548 96460 56604
rect 96460 56548 96516 56604
rect 96516 56548 96520 56604
rect 96456 56544 96520 56548
rect 96536 56604 96600 56608
rect 96536 56548 96540 56604
rect 96540 56548 96596 56604
rect 96596 56548 96600 56604
rect 96536 56544 96600 56548
rect 96616 56604 96680 56608
rect 96616 56548 96620 56604
rect 96620 56548 96676 56604
rect 96676 56548 96680 56604
rect 96616 56544 96680 56548
rect 19576 56060 19640 56064
rect 19576 56004 19580 56060
rect 19580 56004 19636 56060
rect 19636 56004 19640 56060
rect 19576 56000 19640 56004
rect 19656 56060 19720 56064
rect 19656 56004 19660 56060
rect 19660 56004 19716 56060
rect 19716 56004 19720 56060
rect 19656 56000 19720 56004
rect 19736 56060 19800 56064
rect 19736 56004 19740 56060
rect 19740 56004 19796 56060
rect 19796 56004 19800 56060
rect 19736 56000 19800 56004
rect 19816 56060 19880 56064
rect 19816 56004 19820 56060
rect 19820 56004 19876 56060
rect 19876 56004 19880 56060
rect 19816 56000 19880 56004
rect 50296 56060 50360 56064
rect 50296 56004 50300 56060
rect 50300 56004 50356 56060
rect 50356 56004 50360 56060
rect 50296 56000 50360 56004
rect 50376 56060 50440 56064
rect 50376 56004 50380 56060
rect 50380 56004 50436 56060
rect 50436 56004 50440 56060
rect 50376 56000 50440 56004
rect 50456 56060 50520 56064
rect 50456 56004 50460 56060
rect 50460 56004 50516 56060
rect 50516 56004 50520 56060
rect 50456 56000 50520 56004
rect 50536 56060 50600 56064
rect 50536 56004 50540 56060
rect 50540 56004 50596 56060
rect 50596 56004 50600 56060
rect 50536 56000 50600 56004
rect 81016 56060 81080 56064
rect 81016 56004 81020 56060
rect 81020 56004 81076 56060
rect 81076 56004 81080 56060
rect 81016 56000 81080 56004
rect 81096 56060 81160 56064
rect 81096 56004 81100 56060
rect 81100 56004 81156 56060
rect 81156 56004 81160 56060
rect 81096 56000 81160 56004
rect 81176 56060 81240 56064
rect 81176 56004 81180 56060
rect 81180 56004 81236 56060
rect 81236 56004 81240 56060
rect 81176 56000 81240 56004
rect 81256 56060 81320 56064
rect 81256 56004 81260 56060
rect 81260 56004 81316 56060
rect 81316 56004 81320 56060
rect 81256 56000 81320 56004
rect 4216 55516 4280 55520
rect 4216 55460 4220 55516
rect 4220 55460 4276 55516
rect 4276 55460 4280 55516
rect 4216 55456 4280 55460
rect 4296 55516 4360 55520
rect 4296 55460 4300 55516
rect 4300 55460 4356 55516
rect 4356 55460 4360 55516
rect 4296 55456 4360 55460
rect 4376 55516 4440 55520
rect 4376 55460 4380 55516
rect 4380 55460 4436 55516
rect 4436 55460 4440 55516
rect 4376 55456 4440 55460
rect 4456 55516 4520 55520
rect 4456 55460 4460 55516
rect 4460 55460 4516 55516
rect 4516 55460 4520 55516
rect 4456 55456 4520 55460
rect 34936 55516 35000 55520
rect 34936 55460 34940 55516
rect 34940 55460 34996 55516
rect 34996 55460 35000 55516
rect 34936 55456 35000 55460
rect 35016 55516 35080 55520
rect 35016 55460 35020 55516
rect 35020 55460 35076 55516
rect 35076 55460 35080 55516
rect 35016 55456 35080 55460
rect 35096 55516 35160 55520
rect 35096 55460 35100 55516
rect 35100 55460 35156 55516
rect 35156 55460 35160 55516
rect 35096 55456 35160 55460
rect 35176 55516 35240 55520
rect 35176 55460 35180 55516
rect 35180 55460 35236 55516
rect 35236 55460 35240 55516
rect 35176 55456 35240 55460
rect 65656 55516 65720 55520
rect 65656 55460 65660 55516
rect 65660 55460 65716 55516
rect 65716 55460 65720 55516
rect 65656 55456 65720 55460
rect 65736 55516 65800 55520
rect 65736 55460 65740 55516
rect 65740 55460 65796 55516
rect 65796 55460 65800 55516
rect 65736 55456 65800 55460
rect 65816 55516 65880 55520
rect 65816 55460 65820 55516
rect 65820 55460 65876 55516
rect 65876 55460 65880 55516
rect 65816 55456 65880 55460
rect 65896 55516 65960 55520
rect 65896 55460 65900 55516
rect 65900 55460 65956 55516
rect 65956 55460 65960 55516
rect 65896 55456 65960 55460
rect 96376 55516 96440 55520
rect 96376 55460 96380 55516
rect 96380 55460 96436 55516
rect 96436 55460 96440 55516
rect 96376 55456 96440 55460
rect 96456 55516 96520 55520
rect 96456 55460 96460 55516
rect 96460 55460 96516 55516
rect 96516 55460 96520 55516
rect 96456 55456 96520 55460
rect 96536 55516 96600 55520
rect 96536 55460 96540 55516
rect 96540 55460 96596 55516
rect 96596 55460 96600 55516
rect 96536 55456 96600 55460
rect 96616 55516 96680 55520
rect 96616 55460 96620 55516
rect 96620 55460 96676 55516
rect 96676 55460 96680 55516
rect 96616 55456 96680 55460
rect 19576 54972 19640 54976
rect 19576 54916 19580 54972
rect 19580 54916 19636 54972
rect 19636 54916 19640 54972
rect 19576 54912 19640 54916
rect 19656 54972 19720 54976
rect 19656 54916 19660 54972
rect 19660 54916 19716 54972
rect 19716 54916 19720 54972
rect 19656 54912 19720 54916
rect 19736 54972 19800 54976
rect 19736 54916 19740 54972
rect 19740 54916 19796 54972
rect 19796 54916 19800 54972
rect 19736 54912 19800 54916
rect 19816 54972 19880 54976
rect 19816 54916 19820 54972
rect 19820 54916 19876 54972
rect 19876 54916 19880 54972
rect 19816 54912 19880 54916
rect 50296 54972 50360 54976
rect 50296 54916 50300 54972
rect 50300 54916 50356 54972
rect 50356 54916 50360 54972
rect 50296 54912 50360 54916
rect 50376 54972 50440 54976
rect 50376 54916 50380 54972
rect 50380 54916 50436 54972
rect 50436 54916 50440 54972
rect 50376 54912 50440 54916
rect 50456 54972 50520 54976
rect 50456 54916 50460 54972
rect 50460 54916 50516 54972
rect 50516 54916 50520 54972
rect 50456 54912 50520 54916
rect 50536 54972 50600 54976
rect 50536 54916 50540 54972
rect 50540 54916 50596 54972
rect 50596 54916 50600 54972
rect 50536 54912 50600 54916
rect 81016 54972 81080 54976
rect 81016 54916 81020 54972
rect 81020 54916 81076 54972
rect 81076 54916 81080 54972
rect 81016 54912 81080 54916
rect 81096 54972 81160 54976
rect 81096 54916 81100 54972
rect 81100 54916 81156 54972
rect 81156 54916 81160 54972
rect 81096 54912 81160 54916
rect 81176 54972 81240 54976
rect 81176 54916 81180 54972
rect 81180 54916 81236 54972
rect 81236 54916 81240 54972
rect 81176 54912 81240 54916
rect 81256 54972 81320 54976
rect 81256 54916 81260 54972
rect 81260 54916 81316 54972
rect 81316 54916 81320 54972
rect 81256 54912 81320 54916
rect 4216 54428 4280 54432
rect 4216 54372 4220 54428
rect 4220 54372 4276 54428
rect 4276 54372 4280 54428
rect 4216 54368 4280 54372
rect 4296 54428 4360 54432
rect 4296 54372 4300 54428
rect 4300 54372 4356 54428
rect 4356 54372 4360 54428
rect 4296 54368 4360 54372
rect 4376 54428 4440 54432
rect 4376 54372 4380 54428
rect 4380 54372 4436 54428
rect 4436 54372 4440 54428
rect 4376 54368 4440 54372
rect 4456 54428 4520 54432
rect 4456 54372 4460 54428
rect 4460 54372 4516 54428
rect 4516 54372 4520 54428
rect 4456 54368 4520 54372
rect 34936 54428 35000 54432
rect 34936 54372 34940 54428
rect 34940 54372 34996 54428
rect 34996 54372 35000 54428
rect 34936 54368 35000 54372
rect 35016 54428 35080 54432
rect 35016 54372 35020 54428
rect 35020 54372 35076 54428
rect 35076 54372 35080 54428
rect 35016 54368 35080 54372
rect 35096 54428 35160 54432
rect 35096 54372 35100 54428
rect 35100 54372 35156 54428
rect 35156 54372 35160 54428
rect 35096 54368 35160 54372
rect 35176 54428 35240 54432
rect 35176 54372 35180 54428
rect 35180 54372 35236 54428
rect 35236 54372 35240 54428
rect 35176 54368 35240 54372
rect 65656 54428 65720 54432
rect 65656 54372 65660 54428
rect 65660 54372 65716 54428
rect 65716 54372 65720 54428
rect 65656 54368 65720 54372
rect 65736 54428 65800 54432
rect 65736 54372 65740 54428
rect 65740 54372 65796 54428
rect 65796 54372 65800 54428
rect 65736 54368 65800 54372
rect 65816 54428 65880 54432
rect 65816 54372 65820 54428
rect 65820 54372 65876 54428
rect 65876 54372 65880 54428
rect 65816 54368 65880 54372
rect 65896 54428 65960 54432
rect 65896 54372 65900 54428
rect 65900 54372 65956 54428
rect 65956 54372 65960 54428
rect 65896 54368 65960 54372
rect 96376 54428 96440 54432
rect 96376 54372 96380 54428
rect 96380 54372 96436 54428
rect 96436 54372 96440 54428
rect 96376 54368 96440 54372
rect 96456 54428 96520 54432
rect 96456 54372 96460 54428
rect 96460 54372 96516 54428
rect 96516 54372 96520 54428
rect 96456 54368 96520 54372
rect 96536 54428 96600 54432
rect 96536 54372 96540 54428
rect 96540 54372 96596 54428
rect 96596 54372 96600 54428
rect 96536 54368 96600 54372
rect 96616 54428 96680 54432
rect 96616 54372 96620 54428
rect 96620 54372 96676 54428
rect 96676 54372 96680 54428
rect 96616 54368 96680 54372
rect 19576 53884 19640 53888
rect 19576 53828 19580 53884
rect 19580 53828 19636 53884
rect 19636 53828 19640 53884
rect 19576 53824 19640 53828
rect 19656 53884 19720 53888
rect 19656 53828 19660 53884
rect 19660 53828 19716 53884
rect 19716 53828 19720 53884
rect 19656 53824 19720 53828
rect 19736 53884 19800 53888
rect 19736 53828 19740 53884
rect 19740 53828 19796 53884
rect 19796 53828 19800 53884
rect 19736 53824 19800 53828
rect 19816 53884 19880 53888
rect 19816 53828 19820 53884
rect 19820 53828 19876 53884
rect 19876 53828 19880 53884
rect 19816 53824 19880 53828
rect 50296 53884 50360 53888
rect 50296 53828 50300 53884
rect 50300 53828 50356 53884
rect 50356 53828 50360 53884
rect 50296 53824 50360 53828
rect 50376 53884 50440 53888
rect 50376 53828 50380 53884
rect 50380 53828 50436 53884
rect 50436 53828 50440 53884
rect 50376 53824 50440 53828
rect 50456 53884 50520 53888
rect 50456 53828 50460 53884
rect 50460 53828 50516 53884
rect 50516 53828 50520 53884
rect 50456 53824 50520 53828
rect 50536 53884 50600 53888
rect 50536 53828 50540 53884
rect 50540 53828 50596 53884
rect 50596 53828 50600 53884
rect 50536 53824 50600 53828
rect 81016 53884 81080 53888
rect 81016 53828 81020 53884
rect 81020 53828 81076 53884
rect 81076 53828 81080 53884
rect 81016 53824 81080 53828
rect 81096 53884 81160 53888
rect 81096 53828 81100 53884
rect 81100 53828 81156 53884
rect 81156 53828 81160 53884
rect 81096 53824 81160 53828
rect 81176 53884 81240 53888
rect 81176 53828 81180 53884
rect 81180 53828 81236 53884
rect 81236 53828 81240 53884
rect 81176 53824 81240 53828
rect 81256 53884 81320 53888
rect 81256 53828 81260 53884
rect 81260 53828 81316 53884
rect 81316 53828 81320 53884
rect 81256 53824 81320 53828
rect 4216 53340 4280 53344
rect 4216 53284 4220 53340
rect 4220 53284 4276 53340
rect 4276 53284 4280 53340
rect 4216 53280 4280 53284
rect 4296 53340 4360 53344
rect 4296 53284 4300 53340
rect 4300 53284 4356 53340
rect 4356 53284 4360 53340
rect 4296 53280 4360 53284
rect 4376 53340 4440 53344
rect 4376 53284 4380 53340
rect 4380 53284 4436 53340
rect 4436 53284 4440 53340
rect 4376 53280 4440 53284
rect 4456 53340 4520 53344
rect 4456 53284 4460 53340
rect 4460 53284 4516 53340
rect 4516 53284 4520 53340
rect 4456 53280 4520 53284
rect 34936 53340 35000 53344
rect 34936 53284 34940 53340
rect 34940 53284 34996 53340
rect 34996 53284 35000 53340
rect 34936 53280 35000 53284
rect 35016 53340 35080 53344
rect 35016 53284 35020 53340
rect 35020 53284 35076 53340
rect 35076 53284 35080 53340
rect 35016 53280 35080 53284
rect 35096 53340 35160 53344
rect 35096 53284 35100 53340
rect 35100 53284 35156 53340
rect 35156 53284 35160 53340
rect 35096 53280 35160 53284
rect 35176 53340 35240 53344
rect 35176 53284 35180 53340
rect 35180 53284 35236 53340
rect 35236 53284 35240 53340
rect 35176 53280 35240 53284
rect 65656 53340 65720 53344
rect 65656 53284 65660 53340
rect 65660 53284 65716 53340
rect 65716 53284 65720 53340
rect 65656 53280 65720 53284
rect 65736 53340 65800 53344
rect 65736 53284 65740 53340
rect 65740 53284 65796 53340
rect 65796 53284 65800 53340
rect 65736 53280 65800 53284
rect 65816 53340 65880 53344
rect 65816 53284 65820 53340
rect 65820 53284 65876 53340
rect 65876 53284 65880 53340
rect 65816 53280 65880 53284
rect 65896 53340 65960 53344
rect 65896 53284 65900 53340
rect 65900 53284 65956 53340
rect 65956 53284 65960 53340
rect 65896 53280 65960 53284
rect 96376 53340 96440 53344
rect 96376 53284 96380 53340
rect 96380 53284 96436 53340
rect 96436 53284 96440 53340
rect 96376 53280 96440 53284
rect 96456 53340 96520 53344
rect 96456 53284 96460 53340
rect 96460 53284 96516 53340
rect 96516 53284 96520 53340
rect 96456 53280 96520 53284
rect 96536 53340 96600 53344
rect 96536 53284 96540 53340
rect 96540 53284 96596 53340
rect 96596 53284 96600 53340
rect 96536 53280 96600 53284
rect 96616 53340 96680 53344
rect 96616 53284 96620 53340
rect 96620 53284 96676 53340
rect 96676 53284 96680 53340
rect 96616 53280 96680 53284
rect 19576 52796 19640 52800
rect 19576 52740 19580 52796
rect 19580 52740 19636 52796
rect 19636 52740 19640 52796
rect 19576 52736 19640 52740
rect 19656 52796 19720 52800
rect 19656 52740 19660 52796
rect 19660 52740 19716 52796
rect 19716 52740 19720 52796
rect 19656 52736 19720 52740
rect 19736 52796 19800 52800
rect 19736 52740 19740 52796
rect 19740 52740 19796 52796
rect 19796 52740 19800 52796
rect 19736 52736 19800 52740
rect 19816 52796 19880 52800
rect 19816 52740 19820 52796
rect 19820 52740 19876 52796
rect 19876 52740 19880 52796
rect 19816 52736 19880 52740
rect 50296 52796 50360 52800
rect 50296 52740 50300 52796
rect 50300 52740 50356 52796
rect 50356 52740 50360 52796
rect 50296 52736 50360 52740
rect 50376 52796 50440 52800
rect 50376 52740 50380 52796
rect 50380 52740 50436 52796
rect 50436 52740 50440 52796
rect 50376 52736 50440 52740
rect 50456 52796 50520 52800
rect 50456 52740 50460 52796
rect 50460 52740 50516 52796
rect 50516 52740 50520 52796
rect 50456 52736 50520 52740
rect 50536 52796 50600 52800
rect 50536 52740 50540 52796
rect 50540 52740 50596 52796
rect 50596 52740 50600 52796
rect 50536 52736 50600 52740
rect 81016 52796 81080 52800
rect 81016 52740 81020 52796
rect 81020 52740 81076 52796
rect 81076 52740 81080 52796
rect 81016 52736 81080 52740
rect 81096 52796 81160 52800
rect 81096 52740 81100 52796
rect 81100 52740 81156 52796
rect 81156 52740 81160 52796
rect 81096 52736 81160 52740
rect 81176 52796 81240 52800
rect 81176 52740 81180 52796
rect 81180 52740 81236 52796
rect 81236 52740 81240 52796
rect 81176 52736 81240 52740
rect 81256 52796 81320 52800
rect 81256 52740 81260 52796
rect 81260 52740 81316 52796
rect 81316 52740 81320 52796
rect 81256 52736 81320 52740
rect 4216 52252 4280 52256
rect 4216 52196 4220 52252
rect 4220 52196 4276 52252
rect 4276 52196 4280 52252
rect 4216 52192 4280 52196
rect 4296 52252 4360 52256
rect 4296 52196 4300 52252
rect 4300 52196 4356 52252
rect 4356 52196 4360 52252
rect 4296 52192 4360 52196
rect 4376 52252 4440 52256
rect 4376 52196 4380 52252
rect 4380 52196 4436 52252
rect 4436 52196 4440 52252
rect 4376 52192 4440 52196
rect 4456 52252 4520 52256
rect 4456 52196 4460 52252
rect 4460 52196 4516 52252
rect 4516 52196 4520 52252
rect 4456 52192 4520 52196
rect 34936 52252 35000 52256
rect 34936 52196 34940 52252
rect 34940 52196 34996 52252
rect 34996 52196 35000 52252
rect 34936 52192 35000 52196
rect 35016 52252 35080 52256
rect 35016 52196 35020 52252
rect 35020 52196 35076 52252
rect 35076 52196 35080 52252
rect 35016 52192 35080 52196
rect 35096 52252 35160 52256
rect 35096 52196 35100 52252
rect 35100 52196 35156 52252
rect 35156 52196 35160 52252
rect 35096 52192 35160 52196
rect 35176 52252 35240 52256
rect 35176 52196 35180 52252
rect 35180 52196 35236 52252
rect 35236 52196 35240 52252
rect 35176 52192 35240 52196
rect 65656 52252 65720 52256
rect 65656 52196 65660 52252
rect 65660 52196 65716 52252
rect 65716 52196 65720 52252
rect 65656 52192 65720 52196
rect 65736 52252 65800 52256
rect 65736 52196 65740 52252
rect 65740 52196 65796 52252
rect 65796 52196 65800 52252
rect 65736 52192 65800 52196
rect 65816 52252 65880 52256
rect 65816 52196 65820 52252
rect 65820 52196 65876 52252
rect 65876 52196 65880 52252
rect 65816 52192 65880 52196
rect 65896 52252 65960 52256
rect 65896 52196 65900 52252
rect 65900 52196 65956 52252
rect 65956 52196 65960 52252
rect 65896 52192 65960 52196
rect 96376 52252 96440 52256
rect 96376 52196 96380 52252
rect 96380 52196 96436 52252
rect 96436 52196 96440 52252
rect 96376 52192 96440 52196
rect 96456 52252 96520 52256
rect 96456 52196 96460 52252
rect 96460 52196 96516 52252
rect 96516 52196 96520 52252
rect 96456 52192 96520 52196
rect 96536 52252 96600 52256
rect 96536 52196 96540 52252
rect 96540 52196 96596 52252
rect 96596 52196 96600 52252
rect 96536 52192 96600 52196
rect 96616 52252 96680 52256
rect 96616 52196 96620 52252
rect 96620 52196 96676 52252
rect 96676 52196 96680 52252
rect 96616 52192 96680 52196
rect 19576 51708 19640 51712
rect 19576 51652 19580 51708
rect 19580 51652 19636 51708
rect 19636 51652 19640 51708
rect 19576 51648 19640 51652
rect 19656 51708 19720 51712
rect 19656 51652 19660 51708
rect 19660 51652 19716 51708
rect 19716 51652 19720 51708
rect 19656 51648 19720 51652
rect 19736 51708 19800 51712
rect 19736 51652 19740 51708
rect 19740 51652 19796 51708
rect 19796 51652 19800 51708
rect 19736 51648 19800 51652
rect 19816 51708 19880 51712
rect 19816 51652 19820 51708
rect 19820 51652 19876 51708
rect 19876 51652 19880 51708
rect 19816 51648 19880 51652
rect 50296 51708 50360 51712
rect 50296 51652 50300 51708
rect 50300 51652 50356 51708
rect 50356 51652 50360 51708
rect 50296 51648 50360 51652
rect 50376 51708 50440 51712
rect 50376 51652 50380 51708
rect 50380 51652 50436 51708
rect 50436 51652 50440 51708
rect 50376 51648 50440 51652
rect 50456 51708 50520 51712
rect 50456 51652 50460 51708
rect 50460 51652 50516 51708
rect 50516 51652 50520 51708
rect 50456 51648 50520 51652
rect 50536 51708 50600 51712
rect 50536 51652 50540 51708
rect 50540 51652 50596 51708
rect 50596 51652 50600 51708
rect 50536 51648 50600 51652
rect 81016 51708 81080 51712
rect 81016 51652 81020 51708
rect 81020 51652 81076 51708
rect 81076 51652 81080 51708
rect 81016 51648 81080 51652
rect 81096 51708 81160 51712
rect 81096 51652 81100 51708
rect 81100 51652 81156 51708
rect 81156 51652 81160 51708
rect 81096 51648 81160 51652
rect 81176 51708 81240 51712
rect 81176 51652 81180 51708
rect 81180 51652 81236 51708
rect 81236 51652 81240 51708
rect 81176 51648 81240 51652
rect 81256 51708 81320 51712
rect 81256 51652 81260 51708
rect 81260 51652 81316 51708
rect 81316 51652 81320 51708
rect 81256 51648 81320 51652
rect 4216 51164 4280 51168
rect 4216 51108 4220 51164
rect 4220 51108 4276 51164
rect 4276 51108 4280 51164
rect 4216 51104 4280 51108
rect 4296 51164 4360 51168
rect 4296 51108 4300 51164
rect 4300 51108 4356 51164
rect 4356 51108 4360 51164
rect 4296 51104 4360 51108
rect 4376 51164 4440 51168
rect 4376 51108 4380 51164
rect 4380 51108 4436 51164
rect 4436 51108 4440 51164
rect 4376 51104 4440 51108
rect 4456 51164 4520 51168
rect 4456 51108 4460 51164
rect 4460 51108 4516 51164
rect 4516 51108 4520 51164
rect 4456 51104 4520 51108
rect 34936 51164 35000 51168
rect 34936 51108 34940 51164
rect 34940 51108 34996 51164
rect 34996 51108 35000 51164
rect 34936 51104 35000 51108
rect 35016 51164 35080 51168
rect 35016 51108 35020 51164
rect 35020 51108 35076 51164
rect 35076 51108 35080 51164
rect 35016 51104 35080 51108
rect 35096 51164 35160 51168
rect 35096 51108 35100 51164
rect 35100 51108 35156 51164
rect 35156 51108 35160 51164
rect 35096 51104 35160 51108
rect 35176 51164 35240 51168
rect 35176 51108 35180 51164
rect 35180 51108 35236 51164
rect 35236 51108 35240 51164
rect 35176 51104 35240 51108
rect 65656 51164 65720 51168
rect 65656 51108 65660 51164
rect 65660 51108 65716 51164
rect 65716 51108 65720 51164
rect 65656 51104 65720 51108
rect 65736 51164 65800 51168
rect 65736 51108 65740 51164
rect 65740 51108 65796 51164
rect 65796 51108 65800 51164
rect 65736 51104 65800 51108
rect 65816 51164 65880 51168
rect 65816 51108 65820 51164
rect 65820 51108 65876 51164
rect 65876 51108 65880 51164
rect 65816 51104 65880 51108
rect 65896 51164 65960 51168
rect 65896 51108 65900 51164
rect 65900 51108 65956 51164
rect 65956 51108 65960 51164
rect 65896 51104 65960 51108
rect 96376 51164 96440 51168
rect 96376 51108 96380 51164
rect 96380 51108 96436 51164
rect 96436 51108 96440 51164
rect 96376 51104 96440 51108
rect 96456 51164 96520 51168
rect 96456 51108 96460 51164
rect 96460 51108 96516 51164
rect 96516 51108 96520 51164
rect 96456 51104 96520 51108
rect 96536 51164 96600 51168
rect 96536 51108 96540 51164
rect 96540 51108 96596 51164
rect 96596 51108 96600 51164
rect 96536 51104 96600 51108
rect 96616 51164 96680 51168
rect 96616 51108 96620 51164
rect 96620 51108 96676 51164
rect 96676 51108 96680 51164
rect 96616 51104 96680 51108
rect 19576 50620 19640 50624
rect 19576 50564 19580 50620
rect 19580 50564 19636 50620
rect 19636 50564 19640 50620
rect 19576 50560 19640 50564
rect 19656 50620 19720 50624
rect 19656 50564 19660 50620
rect 19660 50564 19716 50620
rect 19716 50564 19720 50620
rect 19656 50560 19720 50564
rect 19736 50620 19800 50624
rect 19736 50564 19740 50620
rect 19740 50564 19796 50620
rect 19796 50564 19800 50620
rect 19736 50560 19800 50564
rect 19816 50620 19880 50624
rect 19816 50564 19820 50620
rect 19820 50564 19876 50620
rect 19876 50564 19880 50620
rect 19816 50560 19880 50564
rect 50296 50620 50360 50624
rect 50296 50564 50300 50620
rect 50300 50564 50356 50620
rect 50356 50564 50360 50620
rect 50296 50560 50360 50564
rect 50376 50620 50440 50624
rect 50376 50564 50380 50620
rect 50380 50564 50436 50620
rect 50436 50564 50440 50620
rect 50376 50560 50440 50564
rect 50456 50620 50520 50624
rect 50456 50564 50460 50620
rect 50460 50564 50516 50620
rect 50516 50564 50520 50620
rect 50456 50560 50520 50564
rect 50536 50620 50600 50624
rect 50536 50564 50540 50620
rect 50540 50564 50596 50620
rect 50596 50564 50600 50620
rect 50536 50560 50600 50564
rect 81016 50620 81080 50624
rect 81016 50564 81020 50620
rect 81020 50564 81076 50620
rect 81076 50564 81080 50620
rect 81016 50560 81080 50564
rect 81096 50620 81160 50624
rect 81096 50564 81100 50620
rect 81100 50564 81156 50620
rect 81156 50564 81160 50620
rect 81096 50560 81160 50564
rect 81176 50620 81240 50624
rect 81176 50564 81180 50620
rect 81180 50564 81236 50620
rect 81236 50564 81240 50620
rect 81176 50560 81240 50564
rect 81256 50620 81320 50624
rect 81256 50564 81260 50620
rect 81260 50564 81316 50620
rect 81316 50564 81320 50620
rect 81256 50560 81320 50564
rect 4216 50076 4280 50080
rect 4216 50020 4220 50076
rect 4220 50020 4276 50076
rect 4276 50020 4280 50076
rect 4216 50016 4280 50020
rect 4296 50076 4360 50080
rect 4296 50020 4300 50076
rect 4300 50020 4356 50076
rect 4356 50020 4360 50076
rect 4296 50016 4360 50020
rect 4376 50076 4440 50080
rect 4376 50020 4380 50076
rect 4380 50020 4436 50076
rect 4436 50020 4440 50076
rect 4376 50016 4440 50020
rect 4456 50076 4520 50080
rect 4456 50020 4460 50076
rect 4460 50020 4516 50076
rect 4516 50020 4520 50076
rect 4456 50016 4520 50020
rect 34936 50076 35000 50080
rect 34936 50020 34940 50076
rect 34940 50020 34996 50076
rect 34996 50020 35000 50076
rect 34936 50016 35000 50020
rect 35016 50076 35080 50080
rect 35016 50020 35020 50076
rect 35020 50020 35076 50076
rect 35076 50020 35080 50076
rect 35016 50016 35080 50020
rect 35096 50076 35160 50080
rect 35096 50020 35100 50076
rect 35100 50020 35156 50076
rect 35156 50020 35160 50076
rect 35096 50016 35160 50020
rect 35176 50076 35240 50080
rect 35176 50020 35180 50076
rect 35180 50020 35236 50076
rect 35236 50020 35240 50076
rect 35176 50016 35240 50020
rect 65656 50076 65720 50080
rect 65656 50020 65660 50076
rect 65660 50020 65716 50076
rect 65716 50020 65720 50076
rect 65656 50016 65720 50020
rect 65736 50076 65800 50080
rect 65736 50020 65740 50076
rect 65740 50020 65796 50076
rect 65796 50020 65800 50076
rect 65736 50016 65800 50020
rect 65816 50076 65880 50080
rect 65816 50020 65820 50076
rect 65820 50020 65876 50076
rect 65876 50020 65880 50076
rect 65816 50016 65880 50020
rect 65896 50076 65960 50080
rect 65896 50020 65900 50076
rect 65900 50020 65956 50076
rect 65956 50020 65960 50076
rect 65896 50016 65960 50020
rect 96376 50076 96440 50080
rect 96376 50020 96380 50076
rect 96380 50020 96436 50076
rect 96436 50020 96440 50076
rect 96376 50016 96440 50020
rect 96456 50076 96520 50080
rect 96456 50020 96460 50076
rect 96460 50020 96516 50076
rect 96516 50020 96520 50076
rect 96456 50016 96520 50020
rect 96536 50076 96600 50080
rect 96536 50020 96540 50076
rect 96540 50020 96596 50076
rect 96596 50020 96600 50076
rect 96536 50016 96600 50020
rect 96616 50076 96680 50080
rect 96616 50020 96620 50076
rect 96620 50020 96676 50076
rect 96676 50020 96680 50076
rect 96616 50016 96680 50020
rect 19576 49532 19640 49536
rect 19576 49476 19580 49532
rect 19580 49476 19636 49532
rect 19636 49476 19640 49532
rect 19576 49472 19640 49476
rect 19656 49532 19720 49536
rect 19656 49476 19660 49532
rect 19660 49476 19716 49532
rect 19716 49476 19720 49532
rect 19656 49472 19720 49476
rect 19736 49532 19800 49536
rect 19736 49476 19740 49532
rect 19740 49476 19796 49532
rect 19796 49476 19800 49532
rect 19736 49472 19800 49476
rect 19816 49532 19880 49536
rect 19816 49476 19820 49532
rect 19820 49476 19876 49532
rect 19876 49476 19880 49532
rect 19816 49472 19880 49476
rect 50296 49532 50360 49536
rect 50296 49476 50300 49532
rect 50300 49476 50356 49532
rect 50356 49476 50360 49532
rect 50296 49472 50360 49476
rect 50376 49532 50440 49536
rect 50376 49476 50380 49532
rect 50380 49476 50436 49532
rect 50436 49476 50440 49532
rect 50376 49472 50440 49476
rect 50456 49532 50520 49536
rect 50456 49476 50460 49532
rect 50460 49476 50516 49532
rect 50516 49476 50520 49532
rect 50456 49472 50520 49476
rect 50536 49532 50600 49536
rect 50536 49476 50540 49532
rect 50540 49476 50596 49532
rect 50596 49476 50600 49532
rect 50536 49472 50600 49476
rect 81016 49532 81080 49536
rect 81016 49476 81020 49532
rect 81020 49476 81076 49532
rect 81076 49476 81080 49532
rect 81016 49472 81080 49476
rect 81096 49532 81160 49536
rect 81096 49476 81100 49532
rect 81100 49476 81156 49532
rect 81156 49476 81160 49532
rect 81096 49472 81160 49476
rect 81176 49532 81240 49536
rect 81176 49476 81180 49532
rect 81180 49476 81236 49532
rect 81236 49476 81240 49532
rect 81176 49472 81240 49476
rect 81256 49532 81320 49536
rect 81256 49476 81260 49532
rect 81260 49476 81316 49532
rect 81316 49476 81320 49532
rect 81256 49472 81320 49476
rect 4216 48988 4280 48992
rect 4216 48932 4220 48988
rect 4220 48932 4276 48988
rect 4276 48932 4280 48988
rect 4216 48928 4280 48932
rect 4296 48988 4360 48992
rect 4296 48932 4300 48988
rect 4300 48932 4356 48988
rect 4356 48932 4360 48988
rect 4296 48928 4360 48932
rect 4376 48988 4440 48992
rect 4376 48932 4380 48988
rect 4380 48932 4436 48988
rect 4436 48932 4440 48988
rect 4376 48928 4440 48932
rect 4456 48988 4520 48992
rect 4456 48932 4460 48988
rect 4460 48932 4516 48988
rect 4516 48932 4520 48988
rect 4456 48928 4520 48932
rect 34936 48988 35000 48992
rect 34936 48932 34940 48988
rect 34940 48932 34996 48988
rect 34996 48932 35000 48988
rect 34936 48928 35000 48932
rect 35016 48988 35080 48992
rect 35016 48932 35020 48988
rect 35020 48932 35076 48988
rect 35076 48932 35080 48988
rect 35016 48928 35080 48932
rect 35096 48988 35160 48992
rect 35096 48932 35100 48988
rect 35100 48932 35156 48988
rect 35156 48932 35160 48988
rect 35096 48928 35160 48932
rect 35176 48988 35240 48992
rect 35176 48932 35180 48988
rect 35180 48932 35236 48988
rect 35236 48932 35240 48988
rect 35176 48928 35240 48932
rect 65656 48988 65720 48992
rect 65656 48932 65660 48988
rect 65660 48932 65716 48988
rect 65716 48932 65720 48988
rect 65656 48928 65720 48932
rect 65736 48988 65800 48992
rect 65736 48932 65740 48988
rect 65740 48932 65796 48988
rect 65796 48932 65800 48988
rect 65736 48928 65800 48932
rect 65816 48988 65880 48992
rect 65816 48932 65820 48988
rect 65820 48932 65876 48988
rect 65876 48932 65880 48988
rect 65816 48928 65880 48932
rect 65896 48988 65960 48992
rect 65896 48932 65900 48988
rect 65900 48932 65956 48988
rect 65956 48932 65960 48988
rect 65896 48928 65960 48932
rect 96376 48988 96440 48992
rect 96376 48932 96380 48988
rect 96380 48932 96436 48988
rect 96436 48932 96440 48988
rect 96376 48928 96440 48932
rect 96456 48988 96520 48992
rect 96456 48932 96460 48988
rect 96460 48932 96516 48988
rect 96516 48932 96520 48988
rect 96456 48928 96520 48932
rect 96536 48988 96600 48992
rect 96536 48932 96540 48988
rect 96540 48932 96596 48988
rect 96596 48932 96600 48988
rect 96536 48928 96600 48932
rect 96616 48988 96680 48992
rect 96616 48932 96620 48988
rect 96620 48932 96676 48988
rect 96676 48932 96680 48988
rect 96616 48928 96680 48932
rect 19576 48444 19640 48448
rect 19576 48388 19580 48444
rect 19580 48388 19636 48444
rect 19636 48388 19640 48444
rect 19576 48384 19640 48388
rect 19656 48444 19720 48448
rect 19656 48388 19660 48444
rect 19660 48388 19716 48444
rect 19716 48388 19720 48444
rect 19656 48384 19720 48388
rect 19736 48444 19800 48448
rect 19736 48388 19740 48444
rect 19740 48388 19796 48444
rect 19796 48388 19800 48444
rect 19736 48384 19800 48388
rect 19816 48444 19880 48448
rect 19816 48388 19820 48444
rect 19820 48388 19876 48444
rect 19876 48388 19880 48444
rect 19816 48384 19880 48388
rect 50296 48444 50360 48448
rect 50296 48388 50300 48444
rect 50300 48388 50356 48444
rect 50356 48388 50360 48444
rect 50296 48384 50360 48388
rect 50376 48444 50440 48448
rect 50376 48388 50380 48444
rect 50380 48388 50436 48444
rect 50436 48388 50440 48444
rect 50376 48384 50440 48388
rect 50456 48444 50520 48448
rect 50456 48388 50460 48444
rect 50460 48388 50516 48444
rect 50516 48388 50520 48444
rect 50456 48384 50520 48388
rect 50536 48444 50600 48448
rect 50536 48388 50540 48444
rect 50540 48388 50596 48444
rect 50596 48388 50600 48444
rect 50536 48384 50600 48388
rect 81016 48444 81080 48448
rect 81016 48388 81020 48444
rect 81020 48388 81076 48444
rect 81076 48388 81080 48444
rect 81016 48384 81080 48388
rect 81096 48444 81160 48448
rect 81096 48388 81100 48444
rect 81100 48388 81156 48444
rect 81156 48388 81160 48444
rect 81096 48384 81160 48388
rect 81176 48444 81240 48448
rect 81176 48388 81180 48444
rect 81180 48388 81236 48444
rect 81236 48388 81240 48444
rect 81176 48384 81240 48388
rect 81256 48444 81320 48448
rect 81256 48388 81260 48444
rect 81260 48388 81316 48444
rect 81316 48388 81320 48444
rect 81256 48384 81320 48388
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 34936 47900 35000 47904
rect 34936 47844 34940 47900
rect 34940 47844 34996 47900
rect 34996 47844 35000 47900
rect 34936 47840 35000 47844
rect 35016 47900 35080 47904
rect 35016 47844 35020 47900
rect 35020 47844 35076 47900
rect 35076 47844 35080 47900
rect 35016 47840 35080 47844
rect 35096 47900 35160 47904
rect 35096 47844 35100 47900
rect 35100 47844 35156 47900
rect 35156 47844 35160 47900
rect 35096 47840 35160 47844
rect 35176 47900 35240 47904
rect 35176 47844 35180 47900
rect 35180 47844 35236 47900
rect 35236 47844 35240 47900
rect 35176 47840 35240 47844
rect 65656 47900 65720 47904
rect 65656 47844 65660 47900
rect 65660 47844 65716 47900
rect 65716 47844 65720 47900
rect 65656 47840 65720 47844
rect 65736 47900 65800 47904
rect 65736 47844 65740 47900
rect 65740 47844 65796 47900
rect 65796 47844 65800 47900
rect 65736 47840 65800 47844
rect 65816 47900 65880 47904
rect 65816 47844 65820 47900
rect 65820 47844 65876 47900
rect 65876 47844 65880 47900
rect 65816 47840 65880 47844
rect 65896 47900 65960 47904
rect 65896 47844 65900 47900
rect 65900 47844 65956 47900
rect 65956 47844 65960 47900
rect 65896 47840 65960 47844
rect 96376 47900 96440 47904
rect 96376 47844 96380 47900
rect 96380 47844 96436 47900
rect 96436 47844 96440 47900
rect 96376 47840 96440 47844
rect 96456 47900 96520 47904
rect 96456 47844 96460 47900
rect 96460 47844 96516 47900
rect 96516 47844 96520 47900
rect 96456 47840 96520 47844
rect 96536 47900 96600 47904
rect 96536 47844 96540 47900
rect 96540 47844 96596 47900
rect 96596 47844 96600 47900
rect 96536 47840 96600 47844
rect 96616 47900 96680 47904
rect 96616 47844 96620 47900
rect 96620 47844 96676 47900
rect 96676 47844 96680 47900
rect 96616 47840 96680 47844
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 50296 47356 50360 47360
rect 50296 47300 50300 47356
rect 50300 47300 50356 47356
rect 50356 47300 50360 47356
rect 50296 47296 50360 47300
rect 50376 47356 50440 47360
rect 50376 47300 50380 47356
rect 50380 47300 50436 47356
rect 50436 47300 50440 47356
rect 50376 47296 50440 47300
rect 50456 47356 50520 47360
rect 50456 47300 50460 47356
rect 50460 47300 50516 47356
rect 50516 47300 50520 47356
rect 50456 47296 50520 47300
rect 50536 47356 50600 47360
rect 50536 47300 50540 47356
rect 50540 47300 50596 47356
rect 50596 47300 50600 47356
rect 50536 47296 50600 47300
rect 81016 47356 81080 47360
rect 81016 47300 81020 47356
rect 81020 47300 81076 47356
rect 81076 47300 81080 47356
rect 81016 47296 81080 47300
rect 81096 47356 81160 47360
rect 81096 47300 81100 47356
rect 81100 47300 81156 47356
rect 81156 47300 81160 47356
rect 81096 47296 81160 47300
rect 81176 47356 81240 47360
rect 81176 47300 81180 47356
rect 81180 47300 81236 47356
rect 81236 47300 81240 47356
rect 81176 47296 81240 47300
rect 81256 47356 81320 47360
rect 81256 47300 81260 47356
rect 81260 47300 81316 47356
rect 81316 47300 81320 47356
rect 81256 47296 81320 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 65656 46812 65720 46816
rect 65656 46756 65660 46812
rect 65660 46756 65716 46812
rect 65716 46756 65720 46812
rect 65656 46752 65720 46756
rect 65736 46812 65800 46816
rect 65736 46756 65740 46812
rect 65740 46756 65796 46812
rect 65796 46756 65800 46812
rect 65736 46752 65800 46756
rect 65816 46812 65880 46816
rect 65816 46756 65820 46812
rect 65820 46756 65876 46812
rect 65876 46756 65880 46812
rect 65816 46752 65880 46756
rect 65896 46812 65960 46816
rect 65896 46756 65900 46812
rect 65900 46756 65956 46812
rect 65956 46756 65960 46812
rect 65896 46752 65960 46756
rect 96376 46812 96440 46816
rect 96376 46756 96380 46812
rect 96380 46756 96436 46812
rect 96436 46756 96440 46812
rect 96376 46752 96440 46756
rect 96456 46812 96520 46816
rect 96456 46756 96460 46812
rect 96460 46756 96516 46812
rect 96516 46756 96520 46812
rect 96456 46752 96520 46756
rect 96536 46812 96600 46816
rect 96536 46756 96540 46812
rect 96540 46756 96596 46812
rect 96596 46756 96600 46812
rect 96536 46752 96600 46756
rect 96616 46812 96680 46816
rect 96616 46756 96620 46812
rect 96620 46756 96676 46812
rect 96676 46756 96680 46812
rect 96616 46752 96680 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 50296 46268 50360 46272
rect 50296 46212 50300 46268
rect 50300 46212 50356 46268
rect 50356 46212 50360 46268
rect 50296 46208 50360 46212
rect 50376 46268 50440 46272
rect 50376 46212 50380 46268
rect 50380 46212 50436 46268
rect 50436 46212 50440 46268
rect 50376 46208 50440 46212
rect 50456 46268 50520 46272
rect 50456 46212 50460 46268
rect 50460 46212 50516 46268
rect 50516 46212 50520 46268
rect 50456 46208 50520 46212
rect 50536 46268 50600 46272
rect 50536 46212 50540 46268
rect 50540 46212 50596 46268
rect 50596 46212 50600 46268
rect 50536 46208 50600 46212
rect 81016 46268 81080 46272
rect 81016 46212 81020 46268
rect 81020 46212 81076 46268
rect 81076 46212 81080 46268
rect 81016 46208 81080 46212
rect 81096 46268 81160 46272
rect 81096 46212 81100 46268
rect 81100 46212 81156 46268
rect 81156 46212 81160 46268
rect 81096 46208 81160 46212
rect 81176 46268 81240 46272
rect 81176 46212 81180 46268
rect 81180 46212 81236 46268
rect 81236 46212 81240 46268
rect 81176 46208 81240 46212
rect 81256 46268 81320 46272
rect 81256 46212 81260 46268
rect 81260 46212 81316 46268
rect 81316 46212 81320 46268
rect 81256 46208 81320 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 65656 45724 65720 45728
rect 65656 45668 65660 45724
rect 65660 45668 65716 45724
rect 65716 45668 65720 45724
rect 65656 45664 65720 45668
rect 65736 45724 65800 45728
rect 65736 45668 65740 45724
rect 65740 45668 65796 45724
rect 65796 45668 65800 45724
rect 65736 45664 65800 45668
rect 65816 45724 65880 45728
rect 65816 45668 65820 45724
rect 65820 45668 65876 45724
rect 65876 45668 65880 45724
rect 65816 45664 65880 45668
rect 65896 45724 65960 45728
rect 65896 45668 65900 45724
rect 65900 45668 65956 45724
rect 65956 45668 65960 45724
rect 65896 45664 65960 45668
rect 96376 45724 96440 45728
rect 96376 45668 96380 45724
rect 96380 45668 96436 45724
rect 96436 45668 96440 45724
rect 96376 45664 96440 45668
rect 96456 45724 96520 45728
rect 96456 45668 96460 45724
rect 96460 45668 96516 45724
rect 96516 45668 96520 45724
rect 96456 45664 96520 45668
rect 96536 45724 96600 45728
rect 96536 45668 96540 45724
rect 96540 45668 96596 45724
rect 96596 45668 96600 45724
rect 96536 45664 96600 45668
rect 96616 45724 96680 45728
rect 96616 45668 96620 45724
rect 96620 45668 96676 45724
rect 96676 45668 96680 45724
rect 96616 45664 96680 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 50296 45180 50360 45184
rect 50296 45124 50300 45180
rect 50300 45124 50356 45180
rect 50356 45124 50360 45180
rect 50296 45120 50360 45124
rect 50376 45180 50440 45184
rect 50376 45124 50380 45180
rect 50380 45124 50436 45180
rect 50436 45124 50440 45180
rect 50376 45120 50440 45124
rect 50456 45180 50520 45184
rect 50456 45124 50460 45180
rect 50460 45124 50516 45180
rect 50516 45124 50520 45180
rect 50456 45120 50520 45124
rect 50536 45180 50600 45184
rect 50536 45124 50540 45180
rect 50540 45124 50596 45180
rect 50596 45124 50600 45180
rect 50536 45120 50600 45124
rect 81016 45180 81080 45184
rect 81016 45124 81020 45180
rect 81020 45124 81076 45180
rect 81076 45124 81080 45180
rect 81016 45120 81080 45124
rect 81096 45180 81160 45184
rect 81096 45124 81100 45180
rect 81100 45124 81156 45180
rect 81156 45124 81160 45180
rect 81096 45120 81160 45124
rect 81176 45180 81240 45184
rect 81176 45124 81180 45180
rect 81180 45124 81236 45180
rect 81236 45124 81240 45180
rect 81176 45120 81240 45124
rect 81256 45180 81320 45184
rect 81256 45124 81260 45180
rect 81260 45124 81316 45180
rect 81316 45124 81320 45180
rect 81256 45120 81320 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 65656 44636 65720 44640
rect 65656 44580 65660 44636
rect 65660 44580 65716 44636
rect 65716 44580 65720 44636
rect 65656 44576 65720 44580
rect 65736 44636 65800 44640
rect 65736 44580 65740 44636
rect 65740 44580 65796 44636
rect 65796 44580 65800 44636
rect 65736 44576 65800 44580
rect 65816 44636 65880 44640
rect 65816 44580 65820 44636
rect 65820 44580 65876 44636
rect 65876 44580 65880 44636
rect 65816 44576 65880 44580
rect 65896 44636 65960 44640
rect 65896 44580 65900 44636
rect 65900 44580 65956 44636
rect 65956 44580 65960 44636
rect 65896 44576 65960 44580
rect 96376 44636 96440 44640
rect 96376 44580 96380 44636
rect 96380 44580 96436 44636
rect 96436 44580 96440 44636
rect 96376 44576 96440 44580
rect 96456 44636 96520 44640
rect 96456 44580 96460 44636
rect 96460 44580 96516 44636
rect 96516 44580 96520 44636
rect 96456 44576 96520 44580
rect 96536 44636 96600 44640
rect 96536 44580 96540 44636
rect 96540 44580 96596 44636
rect 96596 44580 96600 44636
rect 96536 44576 96600 44580
rect 96616 44636 96680 44640
rect 96616 44580 96620 44636
rect 96620 44580 96676 44636
rect 96676 44580 96680 44636
rect 96616 44576 96680 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 50296 44092 50360 44096
rect 50296 44036 50300 44092
rect 50300 44036 50356 44092
rect 50356 44036 50360 44092
rect 50296 44032 50360 44036
rect 50376 44092 50440 44096
rect 50376 44036 50380 44092
rect 50380 44036 50436 44092
rect 50436 44036 50440 44092
rect 50376 44032 50440 44036
rect 50456 44092 50520 44096
rect 50456 44036 50460 44092
rect 50460 44036 50516 44092
rect 50516 44036 50520 44092
rect 50456 44032 50520 44036
rect 50536 44092 50600 44096
rect 50536 44036 50540 44092
rect 50540 44036 50596 44092
rect 50596 44036 50600 44092
rect 50536 44032 50600 44036
rect 81016 44092 81080 44096
rect 81016 44036 81020 44092
rect 81020 44036 81076 44092
rect 81076 44036 81080 44092
rect 81016 44032 81080 44036
rect 81096 44092 81160 44096
rect 81096 44036 81100 44092
rect 81100 44036 81156 44092
rect 81156 44036 81160 44092
rect 81096 44032 81160 44036
rect 81176 44092 81240 44096
rect 81176 44036 81180 44092
rect 81180 44036 81236 44092
rect 81236 44036 81240 44092
rect 81176 44032 81240 44036
rect 81256 44092 81320 44096
rect 81256 44036 81260 44092
rect 81260 44036 81316 44092
rect 81316 44036 81320 44092
rect 81256 44032 81320 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 65656 43548 65720 43552
rect 65656 43492 65660 43548
rect 65660 43492 65716 43548
rect 65716 43492 65720 43548
rect 65656 43488 65720 43492
rect 65736 43548 65800 43552
rect 65736 43492 65740 43548
rect 65740 43492 65796 43548
rect 65796 43492 65800 43548
rect 65736 43488 65800 43492
rect 65816 43548 65880 43552
rect 65816 43492 65820 43548
rect 65820 43492 65876 43548
rect 65876 43492 65880 43548
rect 65816 43488 65880 43492
rect 65896 43548 65960 43552
rect 65896 43492 65900 43548
rect 65900 43492 65956 43548
rect 65956 43492 65960 43548
rect 65896 43488 65960 43492
rect 96376 43548 96440 43552
rect 96376 43492 96380 43548
rect 96380 43492 96436 43548
rect 96436 43492 96440 43548
rect 96376 43488 96440 43492
rect 96456 43548 96520 43552
rect 96456 43492 96460 43548
rect 96460 43492 96516 43548
rect 96516 43492 96520 43548
rect 96456 43488 96520 43492
rect 96536 43548 96600 43552
rect 96536 43492 96540 43548
rect 96540 43492 96596 43548
rect 96596 43492 96600 43548
rect 96536 43488 96600 43492
rect 96616 43548 96680 43552
rect 96616 43492 96620 43548
rect 96620 43492 96676 43548
rect 96676 43492 96680 43548
rect 96616 43488 96680 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 50296 43004 50360 43008
rect 50296 42948 50300 43004
rect 50300 42948 50356 43004
rect 50356 42948 50360 43004
rect 50296 42944 50360 42948
rect 50376 43004 50440 43008
rect 50376 42948 50380 43004
rect 50380 42948 50436 43004
rect 50436 42948 50440 43004
rect 50376 42944 50440 42948
rect 50456 43004 50520 43008
rect 50456 42948 50460 43004
rect 50460 42948 50516 43004
rect 50516 42948 50520 43004
rect 50456 42944 50520 42948
rect 50536 43004 50600 43008
rect 50536 42948 50540 43004
rect 50540 42948 50596 43004
rect 50596 42948 50600 43004
rect 50536 42944 50600 42948
rect 81016 43004 81080 43008
rect 81016 42948 81020 43004
rect 81020 42948 81076 43004
rect 81076 42948 81080 43004
rect 81016 42944 81080 42948
rect 81096 43004 81160 43008
rect 81096 42948 81100 43004
rect 81100 42948 81156 43004
rect 81156 42948 81160 43004
rect 81096 42944 81160 42948
rect 81176 43004 81240 43008
rect 81176 42948 81180 43004
rect 81180 42948 81236 43004
rect 81236 42948 81240 43004
rect 81176 42944 81240 42948
rect 81256 43004 81320 43008
rect 81256 42948 81260 43004
rect 81260 42948 81316 43004
rect 81316 42948 81320 43004
rect 81256 42944 81320 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 65656 42460 65720 42464
rect 65656 42404 65660 42460
rect 65660 42404 65716 42460
rect 65716 42404 65720 42460
rect 65656 42400 65720 42404
rect 65736 42460 65800 42464
rect 65736 42404 65740 42460
rect 65740 42404 65796 42460
rect 65796 42404 65800 42460
rect 65736 42400 65800 42404
rect 65816 42460 65880 42464
rect 65816 42404 65820 42460
rect 65820 42404 65876 42460
rect 65876 42404 65880 42460
rect 65816 42400 65880 42404
rect 65896 42460 65960 42464
rect 65896 42404 65900 42460
rect 65900 42404 65956 42460
rect 65956 42404 65960 42460
rect 65896 42400 65960 42404
rect 96376 42460 96440 42464
rect 96376 42404 96380 42460
rect 96380 42404 96436 42460
rect 96436 42404 96440 42460
rect 96376 42400 96440 42404
rect 96456 42460 96520 42464
rect 96456 42404 96460 42460
rect 96460 42404 96516 42460
rect 96516 42404 96520 42460
rect 96456 42400 96520 42404
rect 96536 42460 96600 42464
rect 96536 42404 96540 42460
rect 96540 42404 96596 42460
rect 96596 42404 96600 42460
rect 96536 42400 96600 42404
rect 96616 42460 96680 42464
rect 96616 42404 96620 42460
rect 96620 42404 96676 42460
rect 96676 42404 96680 42460
rect 96616 42400 96680 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 50296 41916 50360 41920
rect 50296 41860 50300 41916
rect 50300 41860 50356 41916
rect 50356 41860 50360 41916
rect 50296 41856 50360 41860
rect 50376 41916 50440 41920
rect 50376 41860 50380 41916
rect 50380 41860 50436 41916
rect 50436 41860 50440 41916
rect 50376 41856 50440 41860
rect 50456 41916 50520 41920
rect 50456 41860 50460 41916
rect 50460 41860 50516 41916
rect 50516 41860 50520 41916
rect 50456 41856 50520 41860
rect 50536 41916 50600 41920
rect 50536 41860 50540 41916
rect 50540 41860 50596 41916
rect 50596 41860 50600 41916
rect 50536 41856 50600 41860
rect 81016 41916 81080 41920
rect 81016 41860 81020 41916
rect 81020 41860 81076 41916
rect 81076 41860 81080 41916
rect 81016 41856 81080 41860
rect 81096 41916 81160 41920
rect 81096 41860 81100 41916
rect 81100 41860 81156 41916
rect 81156 41860 81160 41916
rect 81096 41856 81160 41860
rect 81176 41916 81240 41920
rect 81176 41860 81180 41916
rect 81180 41860 81236 41916
rect 81236 41860 81240 41916
rect 81176 41856 81240 41860
rect 81256 41916 81320 41920
rect 81256 41860 81260 41916
rect 81260 41860 81316 41916
rect 81316 41860 81320 41916
rect 81256 41856 81320 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 65656 41372 65720 41376
rect 65656 41316 65660 41372
rect 65660 41316 65716 41372
rect 65716 41316 65720 41372
rect 65656 41312 65720 41316
rect 65736 41372 65800 41376
rect 65736 41316 65740 41372
rect 65740 41316 65796 41372
rect 65796 41316 65800 41372
rect 65736 41312 65800 41316
rect 65816 41372 65880 41376
rect 65816 41316 65820 41372
rect 65820 41316 65876 41372
rect 65876 41316 65880 41372
rect 65816 41312 65880 41316
rect 65896 41372 65960 41376
rect 65896 41316 65900 41372
rect 65900 41316 65956 41372
rect 65956 41316 65960 41372
rect 65896 41312 65960 41316
rect 96376 41372 96440 41376
rect 96376 41316 96380 41372
rect 96380 41316 96436 41372
rect 96436 41316 96440 41372
rect 96376 41312 96440 41316
rect 96456 41372 96520 41376
rect 96456 41316 96460 41372
rect 96460 41316 96516 41372
rect 96516 41316 96520 41372
rect 96456 41312 96520 41316
rect 96536 41372 96600 41376
rect 96536 41316 96540 41372
rect 96540 41316 96596 41372
rect 96596 41316 96600 41372
rect 96536 41312 96600 41316
rect 96616 41372 96680 41376
rect 96616 41316 96620 41372
rect 96620 41316 96676 41372
rect 96676 41316 96680 41372
rect 96616 41312 96680 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 50296 40828 50360 40832
rect 50296 40772 50300 40828
rect 50300 40772 50356 40828
rect 50356 40772 50360 40828
rect 50296 40768 50360 40772
rect 50376 40828 50440 40832
rect 50376 40772 50380 40828
rect 50380 40772 50436 40828
rect 50436 40772 50440 40828
rect 50376 40768 50440 40772
rect 50456 40828 50520 40832
rect 50456 40772 50460 40828
rect 50460 40772 50516 40828
rect 50516 40772 50520 40828
rect 50456 40768 50520 40772
rect 50536 40828 50600 40832
rect 50536 40772 50540 40828
rect 50540 40772 50596 40828
rect 50596 40772 50600 40828
rect 50536 40768 50600 40772
rect 81016 40828 81080 40832
rect 81016 40772 81020 40828
rect 81020 40772 81076 40828
rect 81076 40772 81080 40828
rect 81016 40768 81080 40772
rect 81096 40828 81160 40832
rect 81096 40772 81100 40828
rect 81100 40772 81156 40828
rect 81156 40772 81160 40828
rect 81096 40768 81160 40772
rect 81176 40828 81240 40832
rect 81176 40772 81180 40828
rect 81180 40772 81236 40828
rect 81236 40772 81240 40828
rect 81176 40768 81240 40772
rect 81256 40828 81320 40832
rect 81256 40772 81260 40828
rect 81260 40772 81316 40828
rect 81316 40772 81320 40828
rect 81256 40768 81320 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 65656 40284 65720 40288
rect 65656 40228 65660 40284
rect 65660 40228 65716 40284
rect 65716 40228 65720 40284
rect 65656 40224 65720 40228
rect 65736 40284 65800 40288
rect 65736 40228 65740 40284
rect 65740 40228 65796 40284
rect 65796 40228 65800 40284
rect 65736 40224 65800 40228
rect 65816 40284 65880 40288
rect 65816 40228 65820 40284
rect 65820 40228 65876 40284
rect 65876 40228 65880 40284
rect 65816 40224 65880 40228
rect 65896 40284 65960 40288
rect 65896 40228 65900 40284
rect 65900 40228 65956 40284
rect 65956 40228 65960 40284
rect 65896 40224 65960 40228
rect 96376 40284 96440 40288
rect 96376 40228 96380 40284
rect 96380 40228 96436 40284
rect 96436 40228 96440 40284
rect 96376 40224 96440 40228
rect 96456 40284 96520 40288
rect 96456 40228 96460 40284
rect 96460 40228 96516 40284
rect 96516 40228 96520 40284
rect 96456 40224 96520 40228
rect 96536 40284 96600 40288
rect 96536 40228 96540 40284
rect 96540 40228 96596 40284
rect 96596 40228 96600 40284
rect 96536 40224 96600 40228
rect 96616 40284 96680 40288
rect 96616 40228 96620 40284
rect 96620 40228 96676 40284
rect 96676 40228 96680 40284
rect 96616 40224 96680 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 50296 39740 50360 39744
rect 50296 39684 50300 39740
rect 50300 39684 50356 39740
rect 50356 39684 50360 39740
rect 50296 39680 50360 39684
rect 50376 39740 50440 39744
rect 50376 39684 50380 39740
rect 50380 39684 50436 39740
rect 50436 39684 50440 39740
rect 50376 39680 50440 39684
rect 50456 39740 50520 39744
rect 50456 39684 50460 39740
rect 50460 39684 50516 39740
rect 50516 39684 50520 39740
rect 50456 39680 50520 39684
rect 50536 39740 50600 39744
rect 50536 39684 50540 39740
rect 50540 39684 50596 39740
rect 50596 39684 50600 39740
rect 50536 39680 50600 39684
rect 81016 39740 81080 39744
rect 81016 39684 81020 39740
rect 81020 39684 81076 39740
rect 81076 39684 81080 39740
rect 81016 39680 81080 39684
rect 81096 39740 81160 39744
rect 81096 39684 81100 39740
rect 81100 39684 81156 39740
rect 81156 39684 81160 39740
rect 81096 39680 81160 39684
rect 81176 39740 81240 39744
rect 81176 39684 81180 39740
rect 81180 39684 81236 39740
rect 81236 39684 81240 39740
rect 81176 39680 81240 39684
rect 81256 39740 81320 39744
rect 81256 39684 81260 39740
rect 81260 39684 81316 39740
rect 81316 39684 81320 39740
rect 81256 39680 81320 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 65656 39196 65720 39200
rect 65656 39140 65660 39196
rect 65660 39140 65716 39196
rect 65716 39140 65720 39196
rect 65656 39136 65720 39140
rect 65736 39196 65800 39200
rect 65736 39140 65740 39196
rect 65740 39140 65796 39196
rect 65796 39140 65800 39196
rect 65736 39136 65800 39140
rect 65816 39196 65880 39200
rect 65816 39140 65820 39196
rect 65820 39140 65876 39196
rect 65876 39140 65880 39196
rect 65816 39136 65880 39140
rect 65896 39196 65960 39200
rect 65896 39140 65900 39196
rect 65900 39140 65956 39196
rect 65956 39140 65960 39196
rect 65896 39136 65960 39140
rect 96376 39196 96440 39200
rect 96376 39140 96380 39196
rect 96380 39140 96436 39196
rect 96436 39140 96440 39196
rect 96376 39136 96440 39140
rect 96456 39196 96520 39200
rect 96456 39140 96460 39196
rect 96460 39140 96516 39196
rect 96516 39140 96520 39196
rect 96456 39136 96520 39140
rect 96536 39196 96600 39200
rect 96536 39140 96540 39196
rect 96540 39140 96596 39196
rect 96596 39140 96600 39196
rect 96536 39136 96600 39140
rect 96616 39196 96680 39200
rect 96616 39140 96620 39196
rect 96620 39140 96676 39196
rect 96676 39140 96680 39196
rect 96616 39136 96680 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 50296 38652 50360 38656
rect 50296 38596 50300 38652
rect 50300 38596 50356 38652
rect 50356 38596 50360 38652
rect 50296 38592 50360 38596
rect 50376 38652 50440 38656
rect 50376 38596 50380 38652
rect 50380 38596 50436 38652
rect 50436 38596 50440 38652
rect 50376 38592 50440 38596
rect 50456 38652 50520 38656
rect 50456 38596 50460 38652
rect 50460 38596 50516 38652
rect 50516 38596 50520 38652
rect 50456 38592 50520 38596
rect 50536 38652 50600 38656
rect 50536 38596 50540 38652
rect 50540 38596 50596 38652
rect 50596 38596 50600 38652
rect 50536 38592 50600 38596
rect 81016 38652 81080 38656
rect 81016 38596 81020 38652
rect 81020 38596 81076 38652
rect 81076 38596 81080 38652
rect 81016 38592 81080 38596
rect 81096 38652 81160 38656
rect 81096 38596 81100 38652
rect 81100 38596 81156 38652
rect 81156 38596 81160 38652
rect 81096 38592 81160 38596
rect 81176 38652 81240 38656
rect 81176 38596 81180 38652
rect 81180 38596 81236 38652
rect 81236 38596 81240 38652
rect 81176 38592 81240 38596
rect 81256 38652 81320 38656
rect 81256 38596 81260 38652
rect 81260 38596 81316 38652
rect 81316 38596 81320 38652
rect 81256 38592 81320 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 65656 38108 65720 38112
rect 65656 38052 65660 38108
rect 65660 38052 65716 38108
rect 65716 38052 65720 38108
rect 65656 38048 65720 38052
rect 65736 38108 65800 38112
rect 65736 38052 65740 38108
rect 65740 38052 65796 38108
rect 65796 38052 65800 38108
rect 65736 38048 65800 38052
rect 65816 38108 65880 38112
rect 65816 38052 65820 38108
rect 65820 38052 65876 38108
rect 65876 38052 65880 38108
rect 65816 38048 65880 38052
rect 65896 38108 65960 38112
rect 65896 38052 65900 38108
rect 65900 38052 65956 38108
rect 65956 38052 65960 38108
rect 65896 38048 65960 38052
rect 96376 38108 96440 38112
rect 96376 38052 96380 38108
rect 96380 38052 96436 38108
rect 96436 38052 96440 38108
rect 96376 38048 96440 38052
rect 96456 38108 96520 38112
rect 96456 38052 96460 38108
rect 96460 38052 96516 38108
rect 96516 38052 96520 38108
rect 96456 38048 96520 38052
rect 96536 38108 96600 38112
rect 96536 38052 96540 38108
rect 96540 38052 96596 38108
rect 96596 38052 96600 38108
rect 96536 38048 96600 38052
rect 96616 38108 96680 38112
rect 96616 38052 96620 38108
rect 96620 38052 96676 38108
rect 96676 38052 96680 38108
rect 96616 38048 96680 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 50296 37564 50360 37568
rect 50296 37508 50300 37564
rect 50300 37508 50356 37564
rect 50356 37508 50360 37564
rect 50296 37504 50360 37508
rect 50376 37564 50440 37568
rect 50376 37508 50380 37564
rect 50380 37508 50436 37564
rect 50436 37508 50440 37564
rect 50376 37504 50440 37508
rect 50456 37564 50520 37568
rect 50456 37508 50460 37564
rect 50460 37508 50516 37564
rect 50516 37508 50520 37564
rect 50456 37504 50520 37508
rect 50536 37564 50600 37568
rect 50536 37508 50540 37564
rect 50540 37508 50596 37564
rect 50596 37508 50600 37564
rect 50536 37504 50600 37508
rect 81016 37564 81080 37568
rect 81016 37508 81020 37564
rect 81020 37508 81076 37564
rect 81076 37508 81080 37564
rect 81016 37504 81080 37508
rect 81096 37564 81160 37568
rect 81096 37508 81100 37564
rect 81100 37508 81156 37564
rect 81156 37508 81160 37564
rect 81096 37504 81160 37508
rect 81176 37564 81240 37568
rect 81176 37508 81180 37564
rect 81180 37508 81236 37564
rect 81236 37508 81240 37564
rect 81176 37504 81240 37508
rect 81256 37564 81320 37568
rect 81256 37508 81260 37564
rect 81260 37508 81316 37564
rect 81316 37508 81320 37564
rect 81256 37504 81320 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 65656 37020 65720 37024
rect 65656 36964 65660 37020
rect 65660 36964 65716 37020
rect 65716 36964 65720 37020
rect 65656 36960 65720 36964
rect 65736 37020 65800 37024
rect 65736 36964 65740 37020
rect 65740 36964 65796 37020
rect 65796 36964 65800 37020
rect 65736 36960 65800 36964
rect 65816 37020 65880 37024
rect 65816 36964 65820 37020
rect 65820 36964 65876 37020
rect 65876 36964 65880 37020
rect 65816 36960 65880 36964
rect 65896 37020 65960 37024
rect 65896 36964 65900 37020
rect 65900 36964 65956 37020
rect 65956 36964 65960 37020
rect 65896 36960 65960 36964
rect 96376 37020 96440 37024
rect 96376 36964 96380 37020
rect 96380 36964 96436 37020
rect 96436 36964 96440 37020
rect 96376 36960 96440 36964
rect 96456 37020 96520 37024
rect 96456 36964 96460 37020
rect 96460 36964 96516 37020
rect 96516 36964 96520 37020
rect 96456 36960 96520 36964
rect 96536 37020 96600 37024
rect 96536 36964 96540 37020
rect 96540 36964 96596 37020
rect 96596 36964 96600 37020
rect 96536 36960 96600 36964
rect 96616 37020 96680 37024
rect 96616 36964 96620 37020
rect 96620 36964 96676 37020
rect 96676 36964 96680 37020
rect 96616 36960 96680 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 50296 36476 50360 36480
rect 50296 36420 50300 36476
rect 50300 36420 50356 36476
rect 50356 36420 50360 36476
rect 50296 36416 50360 36420
rect 50376 36476 50440 36480
rect 50376 36420 50380 36476
rect 50380 36420 50436 36476
rect 50436 36420 50440 36476
rect 50376 36416 50440 36420
rect 50456 36476 50520 36480
rect 50456 36420 50460 36476
rect 50460 36420 50516 36476
rect 50516 36420 50520 36476
rect 50456 36416 50520 36420
rect 50536 36476 50600 36480
rect 50536 36420 50540 36476
rect 50540 36420 50596 36476
rect 50596 36420 50600 36476
rect 50536 36416 50600 36420
rect 81016 36476 81080 36480
rect 81016 36420 81020 36476
rect 81020 36420 81076 36476
rect 81076 36420 81080 36476
rect 81016 36416 81080 36420
rect 81096 36476 81160 36480
rect 81096 36420 81100 36476
rect 81100 36420 81156 36476
rect 81156 36420 81160 36476
rect 81096 36416 81160 36420
rect 81176 36476 81240 36480
rect 81176 36420 81180 36476
rect 81180 36420 81236 36476
rect 81236 36420 81240 36476
rect 81176 36416 81240 36420
rect 81256 36476 81320 36480
rect 81256 36420 81260 36476
rect 81260 36420 81316 36476
rect 81316 36420 81320 36476
rect 81256 36416 81320 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 65656 35932 65720 35936
rect 65656 35876 65660 35932
rect 65660 35876 65716 35932
rect 65716 35876 65720 35932
rect 65656 35872 65720 35876
rect 65736 35932 65800 35936
rect 65736 35876 65740 35932
rect 65740 35876 65796 35932
rect 65796 35876 65800 35932
rect 65736 35872 65800 35876
rect 65816 35932 65880 35936
rect 65816 35876 65820 35932
rect 65820 35876 65876 35932
rect 65876 35876 65880 35932
rect 65816 35872 65880 35876
rect 65896 35932 65960 35936
rect 65896 35876 65900 35932
rect 65900 35876 65956 35932
rect 65956 35876 65960 35932
rect 65896 35872 65960 35876
rect 96376 35932 96440 35936
rect 96376 35876 96380 35932
rect 96380 35876 96436 35932
rect 96436 35876 96440 35932
rect 96376 35872 96440 35876
rect 96456 35932 96520 35936
rect 96456 35876 96460 35932
rect 96460 35876 96516 35932
rect 96516 35876 96520 35932
rect 96456 35872 96520 35876
rect 96536 35932 96600 35936
rect 96536 35876 96540 35932
rect 96540 35876 96596 35932
rect 96596 35876 96600 35932
rect 96536 35872 96600 35876
rect 96616 35932 96680 35936
rect 96616 35876 96620 35932
rect 96620 35876 96676 35932
rect 96676 35876 96680 35932
rect 96616 35872 96680 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 50296 35388 50360 35392
rect 50296 35332 50300 35388
rect 50300 35332 50356 35388
rect 50356 35332 50360 35388
rect 50296 35328 50360 35332
rect 50376 35388 50440 35392
rect 50376 35332 50380 35388
rect 50380 35332 50436 35388
rect 50436 35332 50440 35388
rect 50376 35328 50440 35332
rect 50456 35388 50520 35392
rect 50456 35332 50460 35388
rect 50460 35332 50516 35388
rect 50516 35332 50520 35388
rect 50456 35328 50520 35332
rect 50536 35388 50600 35392
rect 50536 35332 50540 35388
rect 50540 35332 50596 35388
rect 50596 35332 50600 35388
rect 50536 35328 50600 35332
rect 81016 35388 81080 35392
rect 81016 35332 81020 35388
rect 81020 35332 81076 35388
rect 81076 35332 81080 35388
rect 81016 35328 81080 35332
rect 81096 35388 81160 35392
rect 81096 35332 81100 35388
rect 81100 35332 81156 35388
rect 81156 35332 81160 35388
rect 81096 35328 81160 35332
rect 81176 35388 81240 35392
rect 81176 35332 81180 35388
rect 81180 35332 81236 35388
rect 81236 35332 81240 35388
rect 81176 35328 81240 35332
rect 81256 35388 81320 35392
rect 81256 35332 81260 35388
rect 81260 35332 81316 35388
rect 81316 35332 81320 35388
rect 81256 35328 81320 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 65656 34844 65720 34848
rect 65656 34788 65660 34844
rect 65660 34788 65716 34844
rect 65716 34788 65720 34844
rect 65656 34784 65720 34788
rect 65736 34844 65800 34848
rect 65736 34788 65740 34844
rect 65740 34788 65796 34844
rect 65796 34788 65800 34844
rect 65736 34784 65800 34788
rect 65816 34844 65880 34848
rect 65816 34788 65820 34844
rect 65820 34788 65876 34844
rect 65876 34788 65880 34844
rect 65816 34784 65880 34788
rect 65896 34844 65960 34848
rect 65896 34788 65900 34844
rect 65900 34788 65956 34844
rect 65956 34788 65960 34844
rect 65896 34784 65960 34788
rect 96376 34844 96440 34848
rect 96376 34788 96380 34844
rect 96380 34788 96436 34844
rect 96436 34788 96440 34844
rect 96376 34784 96440 34788
rect 96456 34844 96520 34848
rect 96456 34788 96460 34844
rect 96460 34788 96516 34844
rect 96516 34788 96520 34844
rect 96456 34784 96520 34788
rect 96536 34844 96600 34848
rect 96536 34788 96540 34844
rect 96540 34788 96596 34844
rect 96596 34788 96600 34844
rect 96536 34784 96600 34788
rect 96616 34844 96680 34848
rect 96616 34788 96620 34844
rect 96620 34788 96676 34844
rect 96676 34788 96680 34844
rect 96616 34784 96680 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 50296 34300 50360 34304
rect 50296 34244 50300 34300
rect 50300 34244 50356 34300
rect 50356 34244 50360 34300
rect 50296 34240 50360 34244
rect 50376 34300 50440 34304
rect 50376 34244 50380 34300
rect 50380 34244 50436 34300
rect 50436 34244 50440 34300
rect 50376 34240 50440 34244
rect 50456 34300 50520 34304
rect 50456 34244 50460 34300
rect 50460 34244 50516 34300
rect 50516 34244 50520 34300
rect 50456 34240 50520 34244
rect 50536 34300 50600 34304
rect 50536 34244 50540 34300
rect 50540 34244 50596 34300
rect 50596 34244 50600 34300
rect 50536 34240 50600 34244
rect 81016 34300 81080 34304
rect 81016 34244 81020 34300
rect 81020 34244 81076 34300
rect 81076 34244 81080 34300
rect 81016 34240 81080 34244
rect 81096 34300 81160 34304
rect 81096 34244 81100 34300
rect 81100 34244 81156 34300
rect 81156 34244 81160 34300
rect 81096 34240 81160 34244
rect 81176 34300 81240 34304
rect 81176 34244 81180 34300
rect 81180 34244 81236 34300
rect 81236 34244 81240 34300
rect 81176 34240 81240 34244
rect 81256 34300 81320 34304
rect 81256 34244 81260 34300
rect 81260 34244 81316 34300
rect 81316 34244 81320 34300
rect 81256 34240 81320 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 65656 33756 65720 33760
rect 65656 33700 65660 33756
rect 65660 33700 65716 33756
rect 65716 33700 65720 33756
rect 65656 33696 65720 33700
rect 65736 33756 65800 33760
rect 65736 33700 65740 33756
rect 65740 33700 65796 33756
rect 65796 33700 65800 33756
rect 65736 33696 65800 33700
rect 65816 33756 65880 33760
rect 65816 33700 65820 33756
rect 65820 33700 65876 33756
rect 65876 33700 65880 33756
rect 65816 33696 65880 33700
rect 65896 33756 65960 33760
rect 65896 33700 65900 33756
rect 65900 33700 65956 33756
rect 65956 33700 65960 33756
rect 65896 33696 65960 33700
rect 96376 33756 96440 33760
rect 96376 33700 96380 33756
rect 96380 33700 96436 33756
rect 96436 33700 96440 33756
rect 96376 33696 96440 33700
rect 96456 33756 96520 33760
rect 96456 33700 96460 33756
rect 96460 33700 96516 33756
rect 96516 33700 96520 33756
rect 96456 33696 96520 33700
rect 96536 33756 96600 33760
rect 96536 33700 96540 33756
rect 96540 33700 96596 33756
rect 96596 33700 96600 33756
rect 96536 33696 96600 33700
rect 96616 33756 96680 33760
rect 96616 33700 96620 33756
rect 96620 33700 96676 33756
rect 96676 33700 96680 33756
rect 96616 33696 96680 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 50296 33212 50360 33216
rect 50296 33156 50300 33212
rect 50300 33156 50356 33212
rect 50356 33156 50360 33212
rect 50296 33152 50360 33156
rect 50376 33212 50440 33216
rect 50376 33156 50380 33212
rect 50380 33156 50436 33212
rect 50436 33156 50440 33212
rect 50376 33152 50440 33156
rect 50456 33212 50520 33216
rect 50456 33156 50460 33212
rect 50460 33156 50516 33212
rect 50516 33156 50520 33212
rect 50456 33152 50520 33156
rect 50536 33212 50600 33216
rect 50536 33156 50540 33212
rect 50540 33156 50596 33212
rect 50596 33156 50600 33212
rect 50536 33152 50600 33156
rect 81016 33212 81080 33216
rect 81016 33156 81020 33212
rect 81020 33156 81076 33212
rect 81076 33156 81080 33212
rect 81016 33152 81080 33156
rect 81096 33212 81160 33216
rect 81096 33156 81100 33212
rect 81100 33156 81156 33212
rect 81156 33156 81160 33212
rect 81096 33152 81160 33156
rect 81176 33212 81240 33216
rect 81176 33156 81180 33212
rect 81180 33156 81236 33212
rect 81236 33156 81240 33212
rect 81176 33152 81240 33156
rect 81256 33212 81320 33216
rect 81256 33156 81260 33212
rect 81260 33156 81316 33212
rect 81316 33156 81320 33212
rect 81256 33152 81320 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 65656 32668 65720 32672
rect 65656 32612 65660 32668
rect 65660 32612 65716 32668
rect 65716 32612 65720 32668
rect 65656 32608 65720 32612
rect 65736 32668 65800 32672
rect 65736 32612 65740 32668
rect 65740 32612 65796 32668
rect 65796 32612 65800 32668
rect 65736 32608 65800 32612
rect 65816 32668 65880 32672
rect 65816 32612 65820 32668
rect 65820 32612 65876 32668
rect 65876 32612 65880 32668
rect 65816 32608 65880 32612
rect 65896 32668 65960 32672
rect 65896 32612 65900 32668
rect 65900 32612 65956 32668
rect 65956 32612 65960 32668
rect 65896 32608 65960 32612
rect 96376 32668 96440 32672
rect 96376 32612 96380 32668
rect 96380 32612 96436 32668
rect 96436 32612 96440 32668
rect 96376 32608 96440 32612
rect 96456 32668 96520 32672
rect 96456 32612 96460 32668
rect 96460 32612 96516 32668
rect 96516 32612 96520 32668
rect 96456 32608 96520 32612
rect 96536 32668 96600 32672
rect 96536 32612 96540 32668
rect 96540 32612 96596 32668
rect 96596 32612 96600 32668
rect 96536 32608 96600 32612
rect 96616 32668 96680 32672
rect 96616 32612 96620 32668
rect 96620 32612 96676 32668
rect 96676 32612 96680 32668
rect 96616 32608 96680 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 50296 32124 50360 32128
rect 50296 32068 50300 32124
rect 50300 32068 50356 32124
rect 50356 32068 50360 32124
rect 50296 32064 50360 32068
rect 50376 32124 50440 32128
rect 50376 32068 50380 32124
rect 50380 32068 50436 32124
rect 50436 32068 50440 32124
rect 50376 32064 50440 32068
rect 50456 32124 50520 32128
rect 50456 32068 50460 32124
rect 50460 32068 50516 32124
rect 50516 32068 50520 32124
rect 50456 32064 50520 32068
rect 50536 32124 50600 32128
rect 50536 32068 50540 32124
rect 50540 32068 50596 32124
rect 50596 32068 50600 32124
rect 50536 32064 50600 32068
rect 81016 32124 81080 32128
rect 81016 32068 81020 32124
rect 81020 32068 81076 32124
rect 81076 32068 81080 32124
rect 81016 32064 81080 32068
rect 81096 32124 81160 32128
rect 81096 32068 81100 32124
rect 81100 32068 81156 32124
rect 81156 32068 81160 32124
rect 81096 32064 81160 32068
rect 81176 32124 81240 32128
rect 81176 32068 81180 32124
rect 81180 32068 81236 32124
rect 81236 32068 81240 32124
rect 81176 32064 81240 32068
rect 81256 32124 81320 32128
rect 81256 32068 81260 32124
rect 81260 32068 81316 32124
rect 81316 32068 81320 32124
rect 81256 32064 81320 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 65656 31580 65720 31584
rect 65656 31524 65660 31580
rect 65660 31524 65716 31580
rect 65716 31524 65720 31580
rect 65656 31520 65720 31524
rect 65736 31580 65800 31584
rect 65736 31524 65740 31580
rect 65740 31524 65796 31580
rect 65796 31524 65800 31580
rect 65736 31520 65800 31524
rect 65816 31580 65880 31584
rect 65816 31524 65820 31580
rect 65820 31524 65876 31580
rect 65876 31524 65880 31580
rect 65816 31520 65880 31524
rect 65896 31580 65960 31584
rect 65896 31524 65900 31580
rect 65900 31524 65956 31580
rect 65956 31524 65960 31580
rect 65896 31520 65960 31524
rect 96376 31580 96440 31584
rect 96376 31524 96380 31580
rect 96380 31524 96436 31580
rect 96436 31524 96440 31580
rect 96376 31520 96440 31524
rect 96456 31580 96520 31584
rect 96456 31524 96460 31580
rect 96460 31524 96516 31580
rect 96516 31524 96520 31580
rect 96456 31520 96520 31524
rect 96536 31580 96600 31584
rect 96536 31524 96540 31580
rect 96540 31524 96596 31580
rect 96596 31524 96600 31580
rect 96536 31520 96600 31524
rect 96616 31580 96680 31584
rect 96616 31524 96620 31580
rect 96620 31524 96676 31580
rect 96676 31524 96680 31580
rect 96616 31520 96680 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 50296 31036 50360 31040
rect 50296 30980 50300 31036
rect 50300 30980 50356 31036
rect 50356 30980 50360 31036
rect 50296 30976 50360 30980
rect 50376 31036 50440 31040
rect 50376 30980 50380 31036
rect 50380 30980 50436 31036
rect 50436 30980 50440 31036
rect 50376 30976 50440 30980
rect 50456 31036 50520 31040
rect 50456 30980 50460 31036
rect 50460 30980 50516 31036
rect 50516 30980 50520 31036
rect 50456 30976 50520 30980
rect 50536 31036 50600 31040
rect 50536 30980 50540 31036
rect 50540 30980 50596 31036
rect 50596 30980 50600 31036
rect 50536 30976 50600 30980
rect 81016 31036 81080 31040
rect 81016 30980 81020 31036
rect 81020 30980 81076 31036
rect 81076 30980 81080 31036
rect 81016 30976 81080 30980
rect 81096 31036 81160 31040
rect 81096 30980 81100 31036
rect 81100 30980 81156 31036
rect 81156 30980 81160 31036
rect 81096 30976 81160 30980
rect 81176 31036 81240 31040
rect 81176 30980 81180 31036
rect 81180 30980 81236 31036
rect 81236 30980 81240 31036
rect 81176 30976 81240 30980
rect 81256 31036 81320 31040
rect 81256 30980 81260 31036
rect 81260 30980 81316 31036
rect 81316 30980 81320 31036
rect 81256 30976 81320 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 65656 30492 65720 30496
rect 65656 30436 65660 30492
rect 65660 30436 65716 30492
rect 65716 30436 65720 30492
rect 65656 30432 65720 30436
rect 65736 30492 65800 30496
rect 65736 30436 65740 30492
rect 65740 30436 65796 30492
rect 65796 30436 65800 30492
rect 65736 30432 65800 30436
rect 65816 30492 65880 30496
rect 65816 30436 65820 30492
rect 65820 30436 65876 30492
rect 65876 30436 65880 30492
rect 65816 30432 65880 30436
rect 65896 30492 65960 30496
rect 65896 30436 65900 30492
rect 65900 30436 65956 30492
rect 65956 30436 65960 30492
rect 65896 30432 65960 30436
rect 96376 30492 96440 30496
rect 96376 30436 96380 30492
rect 96380 30436 96436 30492
rect 96436 30436 96440 30492
rect 96376 30432 96440 30436
rect 96456 30492 96520 30496
rect 96456 30436 96460 30492
rect 96460 30436 96516 30492
rect 96516 30436 96520 30492
rect 96456 30432 96520 30436
rect 96536 30492 96600 30496
rect 96536 30436 96540 30492
rect 96540 30436 96596 30492
rect 96596 30436 96600 30492
rect 96536 30432 96600 30436
rect 96616 30492 96680 30496
rect 96616 30436 96620 30492
rect 96620 30436 96676 30492
rect 96676 30436 96680 30492
rect 96616 30432 96680 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 50296 29948 50360 29952
rect 50296 29892 50300 29948
rect 50300 29892 50356 29948
rect 50356 29892 50360 29948
rect 50296 29888 50360 29892
rect 50376 29948 50440 29952
rect 50376 29892 50380 29948
rect 50380 29892 50436 29948
rect 50436 29892 50440 29948
rect 50376 29888 50440 29892
rect 50456 29948 50520 29952
rect 50456 29892 50460 29948
rect 50460 29892 50516 29948
rect 50516 29892 50520 29948
rect 50456 29888 50520 29892
rect 50536 29948 50600 29952
rect 50536 29892 50540 29948
rect 50540 29892 50596 29948
rect 50596 29892 50600 29948
rect 50536 29888 50600 29892
rect 81016 29948 81080 29952
rect 81016 29892 81020 29948
rect 81020 29892 81076 29948
rect 81076 29892 81080 29948
rect 81016 29888 81080 29892
rect 81096 29948 81160 29952
rect 81096 29892 81100 29948
rect 81100 29892 81156 29948
rect 81156 29892 81160 29948
rect 81096 29888 81160 29892
rect 81176 29948 81240 29952
rect 81176 29892 81180 29948
rect 81180 29892 81236 29948
rect 81236 29892 81240 29948
rect 81176 29888 81240 29892
rect 81256 29948 81320 29952
rect 81256 29892 81260 29948
rect 81260 29892 81316 29948
rect 81316 29892 81320 29948
rect 81256 29888 81320 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 65656 29404 65720 29408
rect 65656 29348 65660 29404
rect 65660 29348 65716 29404
rect 65716 29348 65720 29404
rect 65656 29344 65720 29348
rect 65736 29404 65800 29408
rect 65736 29348 65740 29404
rect 65740 29348 65796 29404
rect 65796 29348 65800 29404
rect 65736 29344 65800 29348
rect 65816 29404 65880 29408
rect 65816 29348 65820 29404
rect 65820 29348 65876 29404
rect 65876 29348 65880 29404
rect 65816 29344 65880 29348
rect 65896 29404 65960 29408
rect 65896 29348 65900 29404
rect 65900 29348 65956 29404
rect 65956 29348 65960 29404
rect 65896 29344 65960 29348
rect 96376 29404 96440 29408
rect 96376 29348 96380 29404
rect 96380 29348 96436 29404
rect 96436 29348 96440 29404
rect 96376 29344 96440 29348
rect 96456 29404 96520 29408
rect 96456 29348 96460 29404
rect 96460 29348 96516 29404
rect 96516 29348 96520 29404
rect 96456 29344 96520 29348
rect 96536 29404 96600 29408
rect 96536 29348 96540 29404
rect 96540 29348 96596 29404
rect 96596 29348 96600 29404
rect 96536 29344 96600 29348
rect 96616 29404 96680 29408
rect 96616 29348 96620 29404
rect 96620 29348 96676 29404
rect 96676 29348 96680 29404
rect 96616 29344 96680 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 50296 28860 50360 28864
rect 50296 28804 50300 28860
rect 50300 28804 50356 28860
rect 50356 28804 50360 28860
rect 50296 28800 50360 28804
rect 50376 28860 50440 28864
rect 50376 28804 50380 28860
rect 50380 28804 50436 28860
rect 50436 28804 50440 28860
rect 50376 28800 50440 28804
rect 50456 28860 50520 28864
rect 50456 28804 50460 28860
rect 50460 28804 50516 28860
rect 50516 28804 50520 28860
rect 50456 28800 50520 28804
rect 50536 28860 50600 28864
rect 50536 28804 50540 28860
rect 50540 28804 50596 28860
rect 50596 28804 50600 28860
rect 50536 28800 50600 28804
rect 81016 28860 81080 28864
rect 81016 28804 81020 28860
rect 81020 28804 81076 28860
rect 81076 28804 81080 28860
rect 81016 28800 81080 28804
rect 81096 28860 81160 28864
rect 81096 28804 81100 28860
rect 81100 28804 81156 28860
rect 81156 28804 81160 28860
rect 81096 28800 81160 28804
rect 81176 28860 81240 28864
rect 81176 28804 81180 28860
rect 81180 28804 81236 28860
rect 81236 28804 81240 28860
rect 81176 28800 81240 28804
rect 81256 28860 81320 28864
rect 81256 28804 81260 28860
rect 81260 28804 81316 28860
rect 81316 28804 81320 28860
rect 81256 28800 81320 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 65656 28316 65720 28320
rect 65656 28260 65660 28316
rect 65660 28260 65716 28316
rect 65716 28260 65720 28316
rect 65656 28256 65720 28260
rect 65736 28316 65800 28320
rect 65736 28260 65740 28316
rect 65740 28260 65796 28316
rect 65796 28260 65800 28316
rect 65736 28256 65800 28260
rect 65816 28316 65880 28320
rect 65816 28260 65820 28316
rect 65820 28260 65876 28316
rect 65876 28260 65880 28316
rect 65816 28256 65880 28260
rect 65896 28316 65960 28320
rect 65896 28260 65900 28316
rect 65900 28260 65956 28316
rect 65956 28260 65960 28316
rect 65896 28256 65960 28260
rect 96376 28316 96440 28320
rect 96376 28260 96380 28316
rect 96380 28260 96436 28316
rect 96436 28260 96440 28316
rect 96376 28256 96440 28260
rect 96456 28316 96520 28320
rect 96456 28260 96460 28316
rect 96460 28260 96516 28316
rect 96516 28260 96520 28316
rect 96456 28256 96520 28260
rect 96536 28316 96600 28320
rect 96536 28260 96540 28316
rect 96540 28260 96596 28316
rect 96596 28260 96600 28316
rect 96536 28256 96600 28260
rect 96616 28316 96680 28320
rect 96616 28260 96620 28316
rect 96620 28260 96676 28316
rect 96676 28260 96680 28316
rect 96616 28256 96680 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 50296 27772 50360 27776
rect 50296 27716 50300 27772
rect 50300 27716 50356 27772
rect 50356 27716 50360 27772
rect 50296 27712 50360 27716
rect 50376 27772 50440 27776
rect 50376 27716 50380 27772
rect 50380 27716 50436 27772
rect 50436 27716 50440 27772
rect 50376 27712 50440 27716
rect 50456 27772 50520 27776
rect 50456 27716 50460 27772
rect 50460 27716 50516 27772
rect 50516 27716 50520 27772
rect 50456 27712 50520 27716
rect 50536 27772 50600 27776
rect 50536 27716 50540 27772
rect 50540 27716 50596 27772
rect 50596 27716 50600 27772
rect 50536 27712 50600 27716
rect 81016 27772 81080 27776
rect 81016 27716 81020 27772
rect 81020 27716 81076 27772
rect 81076 27716 81080 27772
rect 81016 27712 81080 27716
rect 81096 27772 81160 27776
rect 81096 27716 81100 27772
rect 81100 27716 81156 27772
rect 81156 27716 81160 27772
rect 81096 27712 81160 27716
rect 81176 27772 81240 27776
rect 81176 27716 81180 27772
rect 81180 27716 81236 27772
rect 81236 27716 81240 27772
rect 81176 27712 81240 27716
rect 81256 27772 81320 27776
rect 81256 27716 81260 27772
rect 81260 27716 81316 27772
rect 81316 27716 81320 27772
rect 81256 27712 81320 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 65656 27228 65720 27232
rect 65656 27172 65660 27228
rect 65660 27172 65716 27228
rect 65716 27172 65720 27228
rect 65656 27168 65720 27172
rect 65736 27228 65800 27232
rect 65736 27172 65740 27228
rect 65740 27172 65796 27228
rect 65796 27172 65800 27228
rect 65736 27168 65800 27172
rect 65816 27228 65880 27232
rect 65816 27172 65820 27228
rect 65820 27172 65876 27228
rect 65876 27172 65880 27228
rect 65816 27168 65880 27172
rect 65896 27228 65960 27232
rect 65896 27172 65900 27228
rect 65900 27172 65956 27228
rect 65956 27172 65960 27228
rect 65896 27168 65960 27172
rect 96376 27228 96440 27232
rect 96376 27172 96380 27228
rect 96380 27172 96436 27228
rect 96436 27172 96440 27228
rect 96376 27168 96440 27172
rect 96456 27228 96520 27232
rect 96456 27172 96460 27228
rect 96460 27172 96516 27228
rect 96516 27172 96520 27228
rect 96456 27168 96520 27172
rect 96536 27228 96600 27232
rect 96536 27172 96540 27228
rect 96540 27172 96596 27228
rect 96596 27172 96600 27228
rect 96536 27168 96600 27172
rect 96616 27228 96680 27232
rect 96616 27172 96620 27228
rect 96620 27172 96676 27228
rect 96676 27172 96680 27228
rect 96616 27168 96680 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 50296 26684 50360 26688
rect 50296 26628 50300 26684
rect 50300 26628 50356 26684
rect 50356 26628 50360 26684
rect 50296 26624 50360 26628
rect 50376 26684 50440 26688
rect 50376 26628 50380 26684
rect 50380 26628 50436 26684
rect 50436 26628 50440 26684
rect 50376 26624 50440 26628
rect 50456 26684 50520 26688
rect 50456 26628 50460 26684
rect 50460 26628 50516 26684
rect 50516 26628 50520 26684
rect 50456 26624 50520 26628
rect 50536 26684 50600 26688
rect 50536 26628 50540 26684
rect 50540 26628 50596 26684
rect 50596 26628 50600 26684
rect 50536 26624 50600 26628
rect 81016 26684 81080 26688
rect 81016 26628 81020 26684
rect 81020 26628 81076 26684
rect 81076 26628 81080 26684
rect 81016 26624 81080 26628
rect 81096 26684 81160 26688
rect 81096 26628 81100 26684
rect 81100 26628 81156 26684
rect 81156 26628 81160 26684
rect 81096 26624 81160 26628
rect 81176 26684 81240 26688
rect 81176 26628 81180 26684
rect 81180 26628 81236 26684
rect 81236 26628 81240 26684
rect 81176 26624 81240 26628
rect 81256 26684 81320 26688
rect 81256 26628 81260 26684
rect 81260 26628 81316 26684
rect 81316 26628 81320 26684
rect 81256 26624 81320 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 65656 26140 65720 26144
rect 65656 26084 65660 26140
rect 65660 26084 65716 26140
rect 65716 26084 65720 26140
rect 65656 26080 65720 26084
rect 65736 26140 65800 26144
rect 65736 26084 65740 26140
rect 65740 26084 65796 26140
rect 65796 26084 65800 26140
rect 65736 26080 65800 26084
rect 65816 26140 65880 26144
rect 65816 26084 65820 26140
rect 65820 26084 65876 26140
rect 65876 26084 65880 26140
rect 65816 26080 65880 26084
rect 65896 26140 65960 26144
rect 65896 26084 65900 26140
rect 65900 26084 65956 26140
rect 65956 26084 65960 26140
rect 65896 26080 65960 26084
rect 96376 26140 96440 26144
rect 96376 26084 96380 26140
rect 96380 26084 96436 26140
rect 96436 26084 96440 26140
rect 96376 26080 96440 26084
rect 96456 26140 96520 26144
rect 96456 26084 96460 26140
rect 96460 26084 96516 26140
rect 96516 26084 96520 26140
rect 96456 26080 96520 26084
rect 96536 26140 96600 26144
rect 96536 26084 96540 26140
rect 96540 26084 96596 26140
rect 96596 26084 96600 26140
rect 96536 26080 96600 26084
rect 96616 26140 96680 26144
rect 96616 26084 96620 26140
rect 96620 26084 96676 26140
rect 96676 26084 96680 26140
rect 96616 26080 96680 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 50296 25596 50360 25600
rect 50296 25540 50300 25596
rect 50300 25540 50356 25596
rect 50356 25540 50360 25596
rect 50296 25536 50360 25540
rect 50376 25596 50440 25600
rect 50376 25540 50380 25596
rect 50380 25540 50436 25596
rect 50436 25540 50440 25596
rect 50376 25536 50440 25540
rect 50456 25596 50520 25600
rect 50456 25540 50460 25596
rect 50460 25540 50516 25596
rect 50516 25540 50520 25596
rect 50456 25536 50520 25540
rect 50536 25596 50600 25600
rect 50536 25540 50540 25596
rect 50540 25540 50596 25596
rect 50596 25540 50600 25596
rect 50536 25536 50600 25540
rect 81016 25596 81080 25600
rect 81016 25540 81020 25596
rect 81020 25540 81076 25596
rect 81076 25540 81080 25596
rect 81016 25536 81080 25540
rect 81096 25596 81160 25600
rect 81096 25540 81100 25596
rect 81100 25540 81156 25596
rect 81156 25540 81160 25596
rect 81096 25536 81160 25540
rect 81176 25596 81240 25600
rect 81176 25540 81180 25596
rect 81180 25540 81236 25596
rect 81236 25540 81240 25596
rect 81176 25536 81240 25540
rect 81256 25596 81320 25600
rect 81256 25540 81260 25596
rect 81260 25540 81316 25596
rect 81316 25540 81320 25596
rect 81256 25536 81320 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 65656 25052 65720 25056
rect 65656 24996 65660 25052
rect 65660 24996 65716 25052
rect 65716 24996 65720 25052
rect 65656 24992 65720 24996
rect 65736 25052 65800 25056
rect 65736 24996 65740 25052
rect 65740 24996 65796 25052
rect 65796 24996 65800 25052
rect 65736 24992 65800 24996
rect 65816 25052 65880 25056
rect 65816 24996 65820 25052
rect 65820 24996 65876 25052
rect 65876 24996 65880 25052
rect 65816 24992 65880 24996
rect 65896 25052 65960 25056
rect 65896 24996 65900 25052
rect 65900 24996 65956 25052
rect 65956 24996 65960 25052
rect 65896 24992 65960 24996
rect 96376 25052 96440 25056
rect 96376 24996 96380 25052
rect 96380 24996 96436 25052
rect 96436 24996 96440 25052
rect 96376 24992 96440 24996
rect 96456 25052 96520 25056
rect 96456 24996 96460 25052
rect 96460 24996 96516 25052
rect 96516 24996 96520 25052
rect 96456 24992 96520 24996
rect 96536 25052 96600 25056
rect 96536 24996 96540 25052
rect 96540 24996 96596 25052
rect 96596 24996 96600 25052
rect 96536 24992 96600 24996
rect 96616 25052 96680 25056
rect 96616 24996 96620 25052
rect 96620 24996 96676 25052
rect 96676 24996 96680 25052
rect 96616 24992 96680 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 50296 24508 50360 24512
rect 50296 24452 50300 24508
rect 50300 24452 50356 24508
rect 50356 24452 50360 24508
rect 50296 24448 50360 24452
rect 50376 24508 50440 24512
rect 50376 24452 50380 24508
rect 50380 24452 50436 24508
rect 50436 24452 50440 24508
rect 50376 24448 50440 24452
rect 50456 24508 50520 24512
rect 50456 24452 50460 24508
rect 50460 24452 50516 24508
rect 50516 24452 50520 24508
rect 50456 24448 50520 24452
rect 50536 24508 50600 24512
rect 50536 24452 50540 24508
rect 50540 24452 50596 24508
rect 50596 24452 50600 24508
rect 50536 24448 50600 24452
rect 81016 24508 81080 24512
rect 81016 24452 81020 24508
rect 81020 24452 81076 24508
rect 81076 24452 81080 24508
rect 81016 24448 81080 24452
rect 81096 24508 81160 24512
rect 81096 24452 81100 24508
rect 81100 24452 81156 24508
rect 81156 24452 81160 24508
rect 81096 24448 81160 24452
rect 81176 24508 81240 24512
rect 81176 24452 81180 24508
rect 81180 24452 81236 24508
rect 81236 24452 81240 24508
rect 81176 24448 81240 24452
rect 81256 24508 81320 24512
rect 81256 24452 81260 24508
rect 81260 24452 81316 24508
rect 81316 24452 81320 24508
rect 81256 24448 81320 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 65656 23964 65720 23968
rect 65656 23908 65660 23964
rect 65660 23908 65716 23964
rect 65716 23908 65720 23964
rect 65656 23904 65720 23908
rect 65736 23964 65800 23968
rect 65736 23908 65740 23964
rect 65740 23908 65796 23964
rect 65796 23908 65800 23964
rect 65736 23904 65800 23908
rect 65816 23964 65880 23968
rect 65816 23908 65820 23964
rect 65820 23908 65876 23964
rect 65876 23908 65880 23964
rect 65816 23904 65880 23908
rect 65896 23964 65960 23968
rect 65896 23908 65900 23964
rect 65900 23908 65956 23964
rect 65956 23908 65960 23964
rect 65896 23904 65960 23908
rect 96376 23964 96440 23968
rect 96376 23908 96380 23964
rect 96380 23908 96436 23964
rect 96436 23908 96440 23964
rect 96376 23904 96440 23908
rect 96456 23964 96520 23968
rect 96456 23908 96460 23964
rect 96460 23908 96516 23964
rect 96516 23908 96520 23964
rect 96456 23904 96520 23908
rect 96536 23964 96600 23968
rect 96536 23908 96540 23964
rect 96540 23908 96596 23964
rect 96596 23908 96600 23964
rect 96536 23904 96600 23908
rect 96616 23964 96680 23968
rect 96616 23908 96620 23964
rect 96620 23908 96676 23964
rect 96676 23908 96680 23964
rect 96616 23904 96680 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 50296 23420 50360 23424
rect 50296 23364 50300 23420
rect 50300 23364 50356 23420
rect 50356 23364 50360 23420
rect 50296 23360 50360 23364
rect 50376 23420 50440 23424
rect 50376 23364 50380 23420
rect 50380 23364 50436 23420
rect 50436 23364 50440 23420
rect 50376 23360 50440 23364
rect 50456 23420 50520 23424
rect 50456 23364 50460 23420
rect 50460 23364 50516 23420
rect 50516 23364 50520 23420
rect 50456 23360 50520 23364
rect 50536 23420 50600 23424
rect 50536 23364 50540 23420
rect 50540 23364 50596 23420
rect 50596 23364 50600 23420
rect 50536 23360 50600 23364
rect 81016 23420 81080 23424
rect 81016 23364 81020 23420
rect 81020 23364 81076 23420
rect 81076 23364 81080 23420
rect 81016 23360 81080 23364
rect 81096 23420 81160 23424
rect 81096 23364 81100 23420
rect 81100 23364 81156 23420
rect 81156 23364 81160 23420
rect 81096 23360 81160 23364
rect 81176 23420 81240 23424
rect 81176 23364 81180 23420
rect 81180 23364 81236 23420
rect 81236 23364 81240 23420
rect 81176 23360 81240 23364
rect 81256 23420 81320 23424
rect 81256 23364 81260 23420
rect 81260 23364 81316 23420
rect 81316 23364 81320 23420
rect 81256 23360 81320 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 65656 22876 65720 22880
rect 65656 22820 65660 22876
rect 65660 22820 65716 22876
rect 65716 22820 65720 22876
rect 65656 22816 65720 22820
rect 65736 22876 65800 22880
rect 65736 22820 65740 22876
rect 65740 22820 65796 22876
rect 65796 22820 65800 22876
rect 65736 22816 65800 22820
rect 65816 22876 65880 22880
rect 65816 22820 65820 22876
rect 65820 22820 65876 22876
rect 65876 22820 65880 22876
rect 65816 22816 65880 22820
rect 65896 22876 65960 22880
rect 65896 22820 65900 22876
rect 65900 22820 65956 22876
rect 65956 22820 65960 22876
rect 65896 22816 65960 22820
rect 96376 22876 96440 22880
rect 96376 22820 96380 22876
rect 96380 22820 96436 22876
rect 96436 22820 96440 22876
rect 96376 22816 96440 22820
rect 96456 22876 96520 22880
rect 96456 22820 96460 22876
rect 96460 22820 96516 22876
rect 96516 22820 96520 22876
rect 96456 22816 96520 22820
rect 96536 22876 96600 22880
rect 96536 22820 96540 22876
rect 96540 22820 96596 22876
rect 96596 22820 96600 22876
rect 96536 22816 96600 22820
rect 96616 22876 96680 22880
rect 96616 22820 96620 22876
rect 96620 22820 96676 22876
rect 96676 22820 96680 22876
rect 96616 22816 96680 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 50296 22332 50360 22336
rect 50296 22276 50300 22332
rect 50300 22276 50356 22332
rect 50356 22276 50360 22332
rect 50296 22272 50360 22276
rect 50376 22332 50440 22336
rect 50376 22276 50380 22332
rect 50380 22276 50436 22332
rect 50436 22276 50440 22332
rect 50376 22272 50440 22276
rect 50456 22332 50520 22336
rect 50456 22276 50460 22332
rect 50460 22276 50516 22332
rect 50516 22276 50520 22332
rect 50456 22272 50520 22276
rect 50536 22332 50600 22336
rect 50536 22276 50540 22332
rect 50540 22276 50596 22332
rect 50596 22276 50600 22332
rect 50536 22272 50600 22276
rect 81016 22332 81080 22336
rect 81016 22276 81020 22332
rect 81020 22276 81076 22332
rect 81076 22276 81080 22332
rect 81016 22272 81080 22276
rect 81096 22332 81160 22336
rect 81096 22276 81100 22332
rect 81100 22276 81156 22332
rect 81156 22276 81160 22332
rect 81096 22272 81160 22276
rect 81176 22332 81240 22336
rect 81176 22276 81180 22332
rect 81180 22276 81236 22332
rect 81236 22276 81240 22332
rect 81176 22272 81240 22276
rect 81256 22332 81320 22336
rect 81256 22276 81260 22332
rect 81260 22276 81316 22332
rect 81316 22276 81320 22332
rect 81256 22272 81320 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 65656 21788 65720 21792
rect 65656 21732 65660 21788
rect 65660 21732 65716 21788
rect 65716 21732 65720 21788
rect 65656 21728 65720 21732
rect 65736 21788 65800 21792
rect 65736 21732 65740 21788
rect 65740 21732 65796 21788
rect 65796 21732 65800 21788
rect 65736 21728 65800 21732
rect 65816 21788 65880 21792
rect 65816 21732 65820 21788
rect 65820 21732 65876 21788
rect 65876 21732 65880 21788
rect 65816 21728 65880 21732
rect 65896 21788 65960 21792
rect 65896 21732 65900 21788
rect 65900 21732 65956 21788
rect 65956 21732 65960 21788
rect 65896 21728 65960 21732
rect 96376 21788 96440 21792
rect 96376 21732 96380 21788
rect 96380 21732 96436 21788
rect 96436 21732 96440 21788
rect 96376 21728 96440 21732
rect 96456 21788 96520 21792
rect 96456 21732 96460 21788
rect 96460 21732 96516 21788
rect 96516 21732 96520 21788
rect 96456 21728 96520 21732
rect 96536 21788 96600 21792
rect 96536 21732 96540 21788
rect 96540 21732 96596 21788
rect 96596 21732 96600 21788
rect 96536 21728 96600 21732
rect 96616 21788 96680 21792
rect 96616 21732 96620 21788
rect 96620 21732 96676 21788
rect 96676 21732 96680 21788
rect 96616 21728 96680 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 50296 21244 50360 21248
rect 50296 21188 50300 21244
rect 50300 21188 50356 21244
rect 50356 21188 50360 21244
rect 50296 21184 50360 21188
rect 50376 21244 50440 21248
rect 50376 21188 50380 21244
rect 50380 21188 50436 21244
rect 50436 21188 50440 21244
rect 50376 21184 50440 21188
rect 50456 21244 50520 21248
rect 50456 21188 50460 21244
rect 50460 21188 50516 21244
rect 50516 21188 50520 21244
rect 50456 21184 50520 21188
rect 50536 21244 50600 21248
rect 50536 21188 50540 21244
rect 50540 21188 50596 21244
rect 50596 21188 50600 21244
rect 50536 21184 50600 21188
rect 81016 21244 81080 21248
rect 81016 21188 81020 21244
rect 81020 21188 81076 21244
rect 81076 21188 81080 21244
rect 81016 21184 81080 21188
rect 81096 21244 81160 21248
rect 81096 21188 81100 21244
rect 81100 21188 81156 21244
rect 81156 21188 81160 21244
rect 81096 21184 81160 21188
rect 81176 21244 81240 21248
rect 81176 21188 81180 21244
rect 81180 21188 81236 21244
rect 81236 21188 81240 21244
rect 81176 21184 81240 21188
rect 81256 21244 81320 21248
rect 81256 21188 81260 21244
rect 81260 21188 81316 21244
rect 81316 21188 81320 21244
rect 81256 21184 81320 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 65656 20700 65720 20704
rect 65656 20644 65660 20700
rect 65660 20644 65716 20700
rect 65716 20644 65720 20700
rect 65656 20640 65720 20644
rect 65736 20700 65800 20704
rect 65736 20644 65740 20700
rect 65740 20644 65796 20700
rect 65796 20644 65800 20700
rect 65736 20640 65800 20644
rect 65816 20700 65880 20704
rect 65816 20644 65820 20700
rect 65820 20644 65876 20700
rect 65876 20644 65880 20700
rect 65816 20640 65880 20644
rect 65896 20700 65960 20704
rect 65896 20644 65900 20700
rect 65900 20644 65956 20700
rect 65956 20644 65960 20700
rect 65896 20640 65960 20644
rect 96376 20700 96440 20704
rect 96376 20644 96380 20700
rect 96380 20644 96436 20700
rect 96436 20644 96440 20700
rect 96376 20640 96440 20644
rect 96456 20700 96520 20704
rect 96456 20644 96460 20700
rect 96460 20644 96516 20700
rect 96516 20644 96520 20700
rect 96456 20640 96520 20644
rect 96536 20700 96600 20704
rect 96536 20644 96540 20700
rect 96540 20644 96596 20700
rect 96596 20644 96600 20700
rect 96536 20640 96600 20644
rect 96616 20700 96680 20704
rect 96616 20644 96620 20700
rect 96620 20644 96676 20700
rect 96676 20644 96680 20700
rect 96616 20640 96680 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 50296 20156 50360 20160
rect 50296 20100 50300 20156
rect 50300 20100 50356 20156
rect 50356 20100 50360 20156
rect 50296 20096 50360 20100
rect 50376 20156 50440 20160
rect 50376 20100 50380 20156
rect 50380 20100 50436 20156
rect 50436 20100 50440 20156
rect 50376 20096 50440 20100
rect 50456 20156 50520 20160
rect 50456 20100 50460 20156
rect 50460 20100 50516 20156
rect 50516 20100 50520 20156
rect 50456 20096 50520 20100
rect 50536 20156 50600 20160
rect 50536 20100 50540 20156
rect 50540 20100 50596 20156
rect 50596 20100 50600 20156
rect 50536 20096 50600 20100
rect 81016 20156 81080 20160
rect 81016 20100 81020 20156
rect 81020 20100 81076 20156
rect 81076 20100 81080 20156
rect 81016 20096 81080 20100
rect 81096 20156 81160 20160
rect 81096 20100 81100 20156
rect 81100 20100 81156 20156
rect 81156 20100 81160 20156
rect 81096 20096 81160 20100
rect 81176 20156 81240 20160
rect 81176 20100 81180 20156
rect 81180 20100 81236 20156
rect 81236 20100 81240 20156
rect 81176 20096 81240 20100
rect 81256 20156 81320 20160
rect 81256 20100 81260 20156
rect 81260 20100 81316 20156
rect 81316 20100 81320 20156
rect 81256 20096 81320 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 65656 19612 65720 19616
rect 65656 19556 65660 19612
rect 65660 19556 65716 19612
rect 65716 19556 65720 19612
rect 65656 19552 65720 19556
rect 65736 19612 65800 19616
rect 65736 19556 65740 19612
rect 65740 19556 65796 19612
rect 65796 19556 65800 19612
rect 65736 19552 65800 19556
rect 65816 19612 65880 19616
rect 65816 19556 65820 19612
rect 65820 19556 65876 19612
rect 65876 19556 65880 19612
rect 65816 19552 65880 19556
rect 65896 19612 65960 19616
rect 65896 19556 65900 19612
rect 65900 19556 65956 19612
rect 65956 19556 65960 19612
rect 65896 19552 65960 19556
rect 96376 19612 96440 19616
rect 96376 19556 96380 19612
rect 96380 19556 96436 19612
rect 96436 19556 96440 19612
rect 96376 19552 96440 19556
rect 96456 19612 96520 19616
rect 96456 19556 96460 19612
rect 96460 19556 96516 19612
rect 96516 19556 96520 19612
rect 96456 19552 96520 19556
rect 96536 19612 96600 19616
rect 96536 19556 96540 19612
rect 96540 19556 96596 19612
rect 96596 19556 96600 19612
rect 96536 19552 96600 19556
rect 96616 19612 96680 19616
rect 96616 19556 96620 19612
rect 96620 19556 96676 19612
rect 96676 19556 96680 19612
rect 96616 19552 96680 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 50296 19068 50360 19072
rect 50296 19012 50300 19068
rect 50300 19012 50356 19068
rect 50356 19012 50360 19068
rect 50296 19008 50360 19012
rect 50376 19068 50440 19072
rect 50376 19012 50380 19068
rect 50380 19012 50436 19068
rect 50436 19012 50440 19068
rect 50376 19008 50440 19012
rect 50456 19068 50520 19072
rect 50456 19012 50460 19068
rect 50460 19012 50516 19068
rect 50516 19012 50520 19068
rect 50456 19008 50520 19012
rect 50536 19068 50600 19072
rect 50536 19012 50540 19068
rect 50540 19012 50596 19068
rect 50596 19012 50600 19068
rect 50536 19008 50600 19012
rect 81016 19068 81080 19072
rect 81016 19012 81020 19068
rect 81020 19012 81076 19068
rect 81076 19012 81080 19068
rect 81016 19008 81080 19012
rect 81096 19068 81160 19072
rect 81096 19012 81100 19068
rect 81100 19012 81156 19068
rect 81156 19012 81160 19068
rect 81096 19008 81160 19012
rect 81176 19068 81240 19072
rect 81176 19012 81180 19068
rect 81180 19012 81236 19068
rect 81236 19012 81240 19068
rect 81176 19008 81240 19012
rect 81256 19068 81320 19072
rect 81256 19012 81260 19068
rect 81260 19012 81316 19068
rect 81316 19012 81320 19068
rect 81256 19008 81320 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 65656 18524 65720 18528
rect 65656 18468 65660 18524
rect 65660 18468 65716 18524
rect 65716 18468 65720 18524
rect 65656 18464 65720 18468
rect 65736 18524 65800 18528
rect 65736 18468 65740 18524
rect 65740 18468 65796 18524
rect 65796 18468 65800 18524
rect 65736 18464 65800 18468
rect 65816 18524 65880 18528
rect 65816 18468 65820 18524
rect 65820 18468 65876 18524
rect 65876 18468 65880 18524
rect 65816 18464 65880 18468
rect 65896 18524 65960 18528
rect 65896 18468 65900 18524
rect 65900 18468 65956 18524
rect 65956 18468 65960 18524
rect 65896 18464 65960 18468
rect 96376 18524 96440 18528
rect 96376 18468 96380 18524
rect 96380 18468 96436 18524
rect 96436 18468 96440 18524
rect 96376 18464 96440 18468
rect 96456 18524 96520 18528
rect 96456 18468 96460 18524
rect 96460 18468 96516 18524
rect 96516 18468 96520 18524
rect 96456 18464 96520 18468
rect 96536 18524 96600 18528
rect 96536 18468 96540 18524
rect 96540 18468 96596 18524
rect 96596 18468 96600 18524
rect 96536 18464 96600 18468
rect 96616 18524 96680 18528
rect 96616 18468 96620 18524
rect 96620 18468 96676 18524
rect 96676 18468 96680 18524
rect 96616 18464 96680 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 50296 17980 50360 17984
rect 50296 17924 50300 17980
rect 50300 17924 50356 17980
rect 50356 17924 50360 17980
rect 50296 17920 50360 17924
rect 50376 17980 50440 17984
rect 50376 17924 50380 17980
rect 50380 17924 50436 17980
rect 50436 17924 50440 17980
rect 50376 17920 50440 17924
rect 50456 17980 50520 17984
rect 50456 17924 50460 17980
rect 50460 17924 50516 17980
rect 50516 17924 50520 17980
rect 50456 17920 50520 17924
rect 50536 17980 50600 17984
rect 50536 17924 50540 17980
rect 50540 17924 50596 17980
rect 50596 17924 50600 17980
rect 50536 17920 50600 17924
rect 81016 17980 81080 17984
rect 81016 17924 81020 17980
rect 81020 17924 81076 17980
rect 81076 17924 81080 17980
rect 81016 17920 81080 17924
rect 81096 17980 81160 17984
rect 81096 17924 81100 17980
rect 81100 17924 81156 17980
rect 81156 17924 81160 17980
rect 81096 17920 81160 17924
rect 81176 17980 81240 17984
rect 81176 17924 81180 17980
rect 81180 17924 81236 17980
rect 81236 17924 81240 17980
rect 81176 17920 81240 17924
rect 81256 17980 81320 17984
rect 81256 17924 81260 17980
rect 81260 17924 81316 17980
rect 81316 17924 81320 17980
rect 81256 17920 81320 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 65656 17436 65720 17440
rect 65656 17380 65660 17436
rect 65660 17380 65716 17436
rect 65716 17380 65720 17436
rect 65656 17376 65720 17380
rect 65736 17436 65800 17440
rect 65736 17380 65740 17436
rect 65740 17380 65796 17436
rect 65796 17380 65800 17436
rect 65736 17376 65800 17380
rect 65816 17436 65880 17440
rect 65816 17380 65820 17436
rect 65820 17380 65876 17436
rect 65876 17380 65880 17436
rect 65816 17376 65880 17380
rect 65896 17436 65960 17440
rect 65896 17380 65900 17436
rect 65900 17380 65956 17436
rect 65956 17380 65960 17436
rect 65896 17376 65960 17380
rect 96376 17436 96440 17440
rect 96376 17380 96380 17436
rect 96380 17380 96436 17436
rect 96436 17380 96440 17436
rect 96376 17376 96440 17380
rect 96456 17436 96520 17440
rect 96456 17380 96460 17436
rect 96460 17380 96516 17436
rect 96516 17380 96520 17436
rect 96456 17376 96520 17380
rect 96536 17436 96600 17440
rect 96536 17380 96540 17436
rect 96540 17380 96596 17436
rect 96596 17380 96600 17436
rect 96536 17376 96600 17380
rect 96616 17436 96680 17440
rect 96616 17380 96620 17436
rect 96620 17380 96676 17436
rect 96676 17380 96680 17436
rect 96616 17376 96680 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 50296 16892 50360 16896
rect 50296 16836 50300 16892
rect 50300 16836 50356 16892
rect 50356 16836 50360 16892
rect 50296 16832 50360 16836
rect 50376 16892 50440 16896
rect 50376 16836 50380 16892
rect 50380 16836 50436 16892
rect 50436 16836 50440 16892
rect 50376 16832 50440 16836
rect 50456 16892 50520 16896
rect 50456 16836 50460 16892
rect 50460 16836 50516 16892
rect 50516 16836 50520 16892
rect 50456 16832 50520 16836
rect 50536 16892 50600 16896
rect 50536 16836 50540 16892
rect 50540 16836 50596 16892
rect 50596 16836 50600 16892
rect 50536 16832 50600 16836
rect 81016 16892 81080 16896
rect 81016 16836 81020 16892
rect 81020 16836 81076 16892
rect 81076 16836 81080 16892
rect 81016 16832 81080 16836
rect 81096 16892 81160 16896
rect 81096 16836 81100 16892
rect 81100 16836 81156 16892
rect 81156 16836 81160 16892
rect 81096 16832 81160 16836
rect 81176 16892 81240 16896
rect 81176 16836 81180 16892
rect 81180 16836 81236 16892
rect 81236 16836 81240 16892
rect 81176 16832 81240 16836
rect 81256 16892 81320 16896
rect 81256 16836 81260 16892
rect 81260 16836 81316 16892
rect 81316 16836 81320 16892
rect 81256 16832 81320 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 65656 16348 65720 16352
rect 65656 16292 65660 16348
rect 65660 16292 65716 16348
rect 65716 16292 65720 16348
rect 65656 16288 65720 16292
rect 65736 16348 65800 16352
rect 65736 16292 65740 16348
rect 65740 16292 65796 16348
rect 65796 16292 65800 16348
rect 65736 16288 65800 16292
rect 65816 16348 65880 16352
rect 65816 16292 65820 16348
rect 65820 16292 65876 16348
rect 65876 16292 65880 16348
rect 65816 16288 65880 16292
rect 65896 16348 65960 16352
rect 65896 16292 65900 16348
rect 65900 16292 65956 16348
rect 65956 16292 65960 16348
rect 65896 16288 65960 16292
rect 96376 16348 96440 16352
rect 96376 16292 96380 16348
rect 96380 16292 96436 16348
rect 96436 16292 96440 16348
rect 96376 16288 96440 16292
rect 96456 16348 96520 16352
rect 96456 16292 96460 16348
rect 96460 16292 96516 16348
rect 96516 16292 96520 16348
rect 96456 16288 96520 16292
rect 96536 16348 96600 16352
rect 96536 16292 96540 16348
rect 96540 16292 96596 16348
rect 96596 16292 96600 16348
rect 96536 16288 96600 16292
rect 96616 16348 96680 16352
rect 96616 16292 96620 16348
rect 96620 16292 96676 16348
rect 96676 16292 96680 16348
rect 96616 16288 96680 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 50296 15804 50360 15808
rect 50296 15748 50300 15804
rect 50300 15748 50356 15804
rect 50356 15748 50360 15804
rect 50296 15744 50360 15748
rect 50376 15804 50440 15808
rect 50376 15748 50380 15804
rect 50380 15748 50436 15804
rect 50436 15748 50440 15804
rect 50376 15744 50440 15748
rect 50456 15804 50520 15808
rect 50456 15748 50460 15804
rect 50460 15748 50516 15804
rect 50516 15748 50520 15804
rect 50456 15744 50520 15748
rect 50536 15804 50600 15808
rect 50536 15748 50540 15804
rect 50540 15748 50596 15804
rect 50596 15748 50600 15804
rect 50536 15744 50600 15748
rect 81016 15804 81080 15808
rect 81016 15748 81020 15804
rect 81020 15748 81076 15804
rect 81076 15748 81080 15804
rect 81016 15744 81080 15748
rect 81096 15804 81160 15808
rect 81096 15748 81100 15804
rect 81100 15748 81156 15804
rect 81156 15748 81160 15804
rect 81096 15744 81160 15748
rect 81176 15804 81240 15808
rect 81176 15748 81180 15804
rect 81180 15748 81236 15804
rect 81236 15748 81240 15804
rect 81176 15744 81240 15748
rect 81256 15804 81320 15808
rect 81256 15748 81260 15804
rect 81260 15748 81316 15804
rect 81316 15748 81320 15804
rect 81256 15744 81320 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 65656 15260 65720 15264
rect 65656 15204 65660 15260
rect 65660 15204 65716 15260
rect 65716 15204 65720 15260
rect 65656 15200 65720 15204
rect 65736 15260 65800 15264
rect 65736 15204 65740 15260
rect 65740 15204 65796 15260
rect 65796 15204 65800 15260
rect 65736 15200 65800 15204
rect 65816 15260 65880 15264
rect 65816 15204 65820 15260
rect 65820 15204 65876 15260
rect 65876 15204 65880 15260
rect 65816 15200 65880 15204
rect 65896 15260 65960 15264
rect 65896 15204 65900 15260
rect 65900 15204 65956 15260
rect 65956 15204 65960 15260
rect 65896 15200 65960 15204
rect 96376 15260 96440 15264
rect 96376 15204 96380 15260
rect 96380 15204 96436 15260
rect 96436 15204 96440 15260
rect 96376 15200 96440 15204
rect 96456 15260 96520 15264
rect 96456 15204 96460 15260
rect 96460 15204 96516 15260
rect 96516 15204 96520 15260
rect 96456 15200 96520 15204
rect 96536 15260 96600 15264
rect 96536 15204 96540 15260
rect 96540 15204 96596 15260
rect 96596 15204 96600 15260
rect 96536 15200 96600 15204
rect 96616 15260 96680 15264
rect 96616 15204 96620 15260
rect 96620 15204 96676 15260
rect 96676 15204 96680 15260
rect 96616 15200 96680 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 50296 14716 50360 14720
rect 50296 14660 50300 14716
rect 50300 14660 50356 14716
rect 50356 14660 50360 14716
rect 50296 14656 50360 14660
rect 50376 14716 50440 14720
rect 50376 14660 50380 14716
rect 50380 14660 50436 14716
rect 50436 14660 50440 14716
rect 50376 14656 50440 14660
rect 50456 14716 50520 14720
rect 50456 14660 50460 14716
rect 50460 14660 50516 14716
rect 50516 14660 50520 14716
rect 50456 14656 50520 14660
rect 50536 14716 50600 14720
rect 50536 14660 50540 14716
rect 50540 14660 50596 14716
rect 50596 14660 50600 14716
rect 50536 14656 50600 14660
rect 81016 14716 81080 14720
rect 81016 14660 81020 14716
rect 81020 14660 81076 14716
rect 81076 14660 81080 14716
rect 81016 14656 81080 14660
rect 81096 14716 81160 14720
rect 81096 14660 81100 14716
rect 81100 14660 81156 14716
rect 81156 14660 81160 14716
rect 81096 14656 81160 14660
rect 81176 14716 81240 14720
rect 81176 14660 81180 14716
rect 81180 14660 81236 14716
rect 81236 14660 81240 14716
rect 81176 14656 81240 14660
rect 81256 14716 81320 14720
rect 81256 14660 81260 14716
rect 81260 14660 81316 14716
rect 81316 14660 81320 14716
rect 81256 14656 81320 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 65656 14172 65720 14176
rect 65656 14116 65660 14172
rect 65660 14116 65716 14172
rect 65716 14116 65720 14172
rect 65656 14112 65720 14116
rect 65736 14172 65800 14176
rect 65736 14116 65740 14172
rect 65740 14116 65796 14172
rect 65796 14116 65800 14172
rect 65736 14112 65800 14116
rect 65816 14172 65880 14176
rect 65816 14116 65820 14172
rect 65820 14116 65876 14172
rect 65876 14116 65880 14172
rect 65816 14112 65880 14116
rect 65896 14172 65960 14176
rect 65896 14116 65900 14172
rect 65900 14116 65956 14172
rect 65956 14116 65960 14172
rect 65896 14112 65960 14116
rect 96376 14172 96440 14176
rect 96376 14116 96380 14172
rect 96380 14116 96436 14172
rect 96436 14116 96440 14172
rect 96376 14112 96440 14116
rect 96456 14172 96520 14176
rect 96456 14116 96460 14172
rect 96460 14116 96516 14172
rect 96516 14116 96520 14172
rect 96456 14112 96520 14116
rect 96536 14172 96600 14176
rect 96536 14116 96540 14172
rect 96540 14116 96596 14172
rect 96596 14116 96600 14172
rect 96536 14112 96600 14116
rect 96616 14172 96680 14176
rect 96616 14116 96620 14172
rect 96620 14116 96676 14172
rect 96676 14116 96680 14172
rect 96616 14112 96680 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 50296 13628 50360 13632
rect 50296 13572 50300 13628
rect 50300 13572 50356 13628
rect 50356 13572 50360 13628
rect 50296 13568 50360 13572
rect 50376 13628 50440 13632
rect 50376 13572 50380 13628
rect 50380 13572 50436 13628
rect 50436 13572 50440 13628
rect 50376 13568 50440 13572
rect 50456 13628 50520 13632
rect 50456 13572 50460 13628
rect 50460 13572 50516 13628
rect 50516 13572 50520 13628
rect 50456 13568 50520 13572
rect 50536 13628 50600 13632
rect 50536 13572 50540 13628
rect 50540 13572 50596 13628
rect 50596 13572 50600 13628
rect 50536 13568 50600 13572
rect 81016 13628 81080 13632
rect 81016 13572 81020 13628
rect 81020 13572 81076 13628
rect 81076 13572 81080 13628
rect 81016 13568 81080 13572
rect 81096 13628 81160 13632
rect 81096 13572 81100 13628
rect 81100 13572 81156 13628
rect 81156 13572 81160 13628
rect 81096 13568 81160 13572
rect 81176 13628 81240 13632
rect 81176 13572 81180 13628
rect 81180 13572 81236 13628
rect 81236 13572 81240 13628
rect 81176 13568 81240 13572
rect 81256 13628 81320 13632
rect 81256 13572 81260 13628
rect 81260 13572 81316 13628
rect 81316 13572 81320 13628
rect 81256 13568 81320 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 65656 13084 65720 13088
rect 65656 13028 65660 13084
rect 65660 13028 65716 13084
rect 65716 13028 65720 13084
rect 65656 13024 65720 13028
rect 65736 13084 65800 13088
rect 65736 13028 65740 13084
rect 65740 13028 65796 13084
rect 65796 13028 65800 13084
rect 65736 13024 65800 13028
rect 65816 13084 65880 13088
rect 65816 13028 65820 13084
rect 65820 13028 65876 13084
rect 65876 13028 65880 13084
rect 65816 13024 65880 13028
rect 65896 13084 65960 13088
rect 65896 13028 65900 13084
rect 65900 13028 65956 13084
rect 65956 13028 65960 13084
rect 65896 13024 65960 13028
rect 96376 13084 96440 13088
rect 96376 13028 96380 13084
rect 96380 13028 96436 13084
rect 96436 13028 96440 13084
rect 96376 13024 96440 13028
rect 96456 13084 96520 13088
rect 96456 13028 96460 13084
rect 96460 13028 96516 13084
rect 96516 13028 96520 13084
rect 96456 13024 96520 13028
rect 96536 13084 96600 13088
rect 96536 13028 96540 13084
rect 96540 13028 96596 13084
rect 96596 13028 96600 13084
rect 96536 13024 96600 13028
rect 96616 13084 96680 13088
rect 96616 13028 96620 13084
rect 96620 13028 96676 13084
rect 96676 13028 96680 13084
rect 96616 13024 96680 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 50296 12540 50360 12544
rect 50296 12484 50300 12540
rect 50300 12484 50356 12540
rect 50356 12484 50360 12540
rect 50296 12480 50360 12484
rect 50376 12540 50440 12544
rect 50376 12484 50380 12540
rect 50380 12484 50436 12540
rect 50436 12484 50440 12540
rect 50376 12480 50440 12484
rect 50456 12540 50520 12544
rect 50456 12484 50460 12540
rect 50460 12484 50516 12540
rect 50516 12484 50520 12540
rect 50456 12480 50520 12484
rect 50536 12540 50600 12544
rect 50536 12484 50540 12540
rect 50540 12484 50596 12540
rect 50596 12484 50600 12540
rect 50536 12480 50600 12484
rect 81016 12540 81080 12544
rect 81016 12484 81020 12540
rect 81020 12484 81076 12540
rect 81076 12484 81080 12540
rect 81016 12480 81080 12484
rect 81096 12540 81160 12544
rect 81096 12484 81100 12540
rect 81100 12484 81156 12540
rect 81156 12484 81160 12540
rect 81096 12480 81160 12484
rect 81176 12540 81240 12544
rect 81176 12484 81180 12540
rect 81180 12484 81236 12540
rect 81236 12484 81240 12540
rect 81176 12480 81240 12484
rect 81256 12540 81320 12544
rect 81256 12484 81260 12540
rect 81260 12484 81316 12540
rect 81316 12484 81320 12540
rect 81256 12480 81320 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 65656 11996 65720 12000
rect 65656 11940 65660 11996
rect 65660 11940 65716 11996
rect 65716 11940 65720 11996
rect 65656 11936 65720 11940
rect 65736 11996 65800 12000
rect 65736 11940 65740 11996
rect 65740 11940 65796 11996
rect 65796 11940 65800 11996
rect 65736 11936 65800 11940
rect 65816 11996 65880 12000
rect 65816 11940 65820 11996
rect 65820 11940 65876 11996
rect 65876 11940 65880 11996
rect 65816 11936 65880 11940
rect 65896 11996 65960 12000
rect 65896 11940 65900 11996
rect 65900 11940 65956 11996
rect 65956 11940 65960 11996
rect 65896 11936 65960 11940
rect 96376 11996 96440 12000
rect 96376 11940 96380 11996
rect 96380 11940 96436 11996
rect 96436 11940 96440 11996
rect 96376 11936 96440 11940
rect 96456 11996 96520 12000
rect 96456 11940 96460 11996
rect 96460 11940 96516 11996
rect 96516 11940 96520 11996
rect 96456 11936 96520 11940
rect 96536 11996 96600 12000
rect 96536 11940 96540 11996
rect 96540 11940 96596 11996
rect 96596 11940 96600 11996
rect 96536 11936 96600 11940
rect 96616 11996 96680 12000
rect 96616 11940 96620 11996
rect 96620 11940 96676 11996
rect 96676 11940 96680 11996
rect 96616 11936 96680 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 50296 11452 50360 11456
rect 50296 11396 50300 11452
rect 50300 11396 50356 11452
rect 50356 11396 50360 11452
rect 50296 11392 50360 11396
rect 50376 11452 50440 11456
rect 50376 11396 50380 11452
rect 50380 11396 50436 11452
rect 50436 11396 50440 11452
rect 50376 11392 50440 11396
rect 50456 11452 50520 11456
rect 50456 11396 50460 11452
rect 50460 11396 50516 11452
rect 50516 11396 50520 11452
rect 50456 11392 50520 11396
rect 50536 11452 50600 11456
rect 50536 11396 50540 11452
rect 50540 11396 50596 11452
rect 50596 11396 50600 11452
rect 50536 11392 50600 11396
rect 81016 11452 81080 11456
rect 81016 11396 81020 11452
rect 81020 11396 81076 11452
rect 81076 11396 81080 11452
rect 81016 11392 81080 11396
rect 81096 11452 81160 11456
rect 81096 11396 81100 11452
rect 81100 11396 81156 11452
rect 81156 11396 81160 11452
rect 81096 11392 81160 11396
rect 81176 11452 81240 11456
rect 81176 11396 81180 11452
rect 81180 11396 81236 11452
rect 81236 11396 81240 11452
rect 81176 11392 81240 11396
rect 81256 11452 81320 11456
rect 81256 11396 81260 11452
rect 81260 11396 81316 11452
rect 81316 11396 81320 11452
rect 81256 11392 81320 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 65656 10908 65720 10912
rect 65656 10852 65660 10908
rect 65660 10852 65716 10908
rect 65716 10852 65720 10908
rect 65656 10848 65720 10852
rect 65736 10908 65800 10912
rect 65736 10852 65740 10908
rect 65740 10852 65796 10908
rect 65796 10852 65800 10908
rect 65736 10848 65800 10852
rect 65816 10908 65880 10912
rect 65816 10852 65820 10908
rect 65820 10852 65876 10908
rect 65876 10852 65880 10908
rect 65816 10848 65880 10852
rect 65896 10908 65960 10912
rect 65896 10852 65900 10908
rect 65900 10852 65956 10908
rect 65956 10852 65960 10908
rect 65896 10848 65960 10852
rect 96376 10908 96440 10912
rect 96376 10852 96380 10908
rect 96380 10852 96436 10908
rect 96436 10852 96440 10908
rect 96376 10848 96440 10852
rect 96456 10908 96520 10912
rect 96456 10852 96460 10908
rect 96460 10852 96516 10908
rect 96516 10852 96520 10908
rect 96456 10848 96520 10852
rect 96536 10908 96600 10912
rect 96536 10852 96540 10908
rect 96540 10852 96596 10908
rect 96596 10852 96600 10908
rect 96536 10848 96600 10852
rect 96616 10908 96680 10912
rect 96616 10852 96620 10908
rect 96620 10852 96676 10908
rect 96676 10852 96680 10908
rect 96616 10848 96680 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 50296 10364 50360 10368
rect 50296 10308 50300 10364
rect 50300 10308 50356 10364
rect 50356 10308 50360 10364
rect 50296 10304 50360 10308
rect 50376 10364 50440 10368
rect 50376 10308 50380 10364
rect 50380 10308 50436 10364
rect 50436 10308 50440 10364
rect 50376 10304 50440 10308
rect 50456 10364 50520 10368
rect 50456 10308 50460 10364
rect 50460 10308 50516 10364
rect 50516 10308 50520 10364
rect 50456 10304 50520 10308
rect 50536 10364 50600 10368
rect 50536 10308 50540 10364
rect 50540 10308 50596 10364
rect 50596 10308 50600 10364
rect 50536 10304 50600 10308
rect 81016 10364 81080 10368
rect 81016 10308 81020 10364
rect 81020 10308 81076 10364
rect 81076 10308 81080 10364
rect 81016 10304 81080 10308
rect 81096 10364 81160 10368
rect 81096 10308 81100 10364
rect 81100 10308 81156 10364
rect 81156 10308 81160 10364
rect 81096 10304 81160 10308
rect 81176 10364 81240 10368
rect 81176 10308 81180 10364
rect 81180 10308 81236 10364
rect 81236 10308 81240 10364
rect 81176 10304 81240 10308
rect 81256 10364 81320 10368
rect 81256 10308 81260 10364
rect 81260 10308 81316 10364
rect 81316 10308 81320 10364
rect 81256 10304 81320 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 65656 9820 65720 9824
rect 65656 9764 65660 9820
rect 65660 9764 65716 9820
rect 65716 9764 65720 9820
rect 65656 9760 65720 9764
rect 65736 9820 65800 9824
rect 65736 9764 65740 9820
rect 65740 9764 65796 9820
rect 65796 9764 65800 9820
rect 65736 9760 65800 9764
rect 65816 9820 65880 9824
rect 65816 9764 65820 9820
rect 65820 9764 65876 9820
rect 65876 9764 65880 9820
rect 65816 9760 65880 9764
rect 65896 9820 65960 9824
rect 65896 9764 65900 9820
rect 65900 9764 65956 9820
rect 65956 9764 65960 9820
rect 65896 9760 65960 9764
rect 96376 9820 96440 9824
rect 96376 9764 96380 9820
rect 96380 9764 96436 9820
rect 96436 9764 96440 9820
rect 96376 9760 96440 9764
rect 96456 9820 96520 9824
rect 96456 9764 96460 9820
rect 96460 9764 96516 9820
rect 96516 9764 96520 9820
rect 96456 9760 96520 9764
rect 96536 9820 96600 9824
rect 96536 9764 96540 9820
rect 96540 9764 96596 9820
rect 96596 9764 96600 9820
rect 96536 9760 96600 9764
rect 96616 9820 96680 9824
rect 96616 9764 96620 9820
rect 96620 9764 96676 9820
rect 96676 9764 96680 9820
rect 96616 9760 96680 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 50296 9276 50360 9280
rect 50296 9220 50300 9276
rect 50300 9220 50356 9276
rect 50356 9220 50360 9276
rect 50296 9216 50360 9220
rect 50376 9276 50440 9280
rect 50376 9220 50380 9276
rect 50380 9220 50436 9276
rect 50436 9220 50440 9276
rect 50376 9216 50440 9220
rect 50456 9276 50520 9280
rect 50456 9220 50460 9276
rect 50460 9220 50516 9276
rect 50516 9220 50520 9276
rect 50456 9216 50520 9220
rect 50536 9276 50600 9280
rect 50536 9220 50540 9276
rect 50540 9220 50596 9276
rect 50596 9220 50600 9276
rect 50536 9216 50600 9220
rect 81016 9276 81080 9280
rect 81016 9220 81020 9276
rect 81020 9220 81076 9276
rect 81076 9220 81080 9276
rect 81016 9216 81080 9220
rect 81096 9276 81160 9280
rect 81096 9220 81100 9276
rect 81100 9220 81156 9276
rect 81156 9220 81160 9276
rect 81096 9216 81160 9220
rect 81176 9276 81240 9280
rect 81176 9220 81180 9276
rect 81180 9220 81236 9276
rect 81236 9220 81240 9276
rect 81176 9216 81240 9220
rect 81256 9276 81320 9280
rect 81256 9220 81260 9276
rect 81260 9220 81316 9276
rect 81316 9220 81320 9276
rect 81256 9216 81320 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 65656 8732 65720 8736
rect 65656 8676 65660 8732
rect 65660 8676 65716 8732
rect 65716 8676 65720 8732
rect 65656 8672 65720 8676
rect 65736 8732 65800 8736
rect 65736 8676 65740 8732
rect 65740 8676 65796 8732
rect 65796 8676 65800 8732
rect 65736 8672 65800 8676
rect 65816 8732 65880 8736
rect 65816 8676 65820 8732
rect 65820 8676 65876 8732
rect 65876 8676 65880 8732
rect 65816 8672 65880 8676
rect 65896 8732 65960 8736
rect 65896 8676 65900 8732
rect 65900 8676 65956 8732
rect 65956 8676 65960 8732
rect 65896 8672 65960 8676
rect 96376 8732 96440 8736
rect 96376 8676 96380 8732
rect 96380 8676 96436 8732
rect 96436 8676 96440 8732
rect 96376 8672 96440 8676
rect 96456 8732 96520 8736
rect 96456 8676 96460 8732
rect 96460 8676 96516 8732
rect 96516 8676 96520 8732
rect 96456 8672 96520 8676
rect 96536 8732 96600 8736
rect 96536 8676 96540 8732
rect 96540 8676 96596 8732
rect 96596 8676 96600 8732
rect 96536 8672 96600 8676
rect 96616 8732 96680 8736
rect 96616 8676 96620 8732
rect 96620 8676 96676 8732
rect 96676 8676 96680 8732
rect 96616 8672 96680 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 50296 8188 50360 8192
rect 50296 8132 50300 8188
rect 50300 8132 50356 8188
rect 50356 8132 50360 8188
rect 50296 8128 50360 8132
rect 50376 8188 50440 8192
rect 50376 8132 50380 8188
rect 50380 8132 50436 8188
rect 50436 8132 50440 8188
rect 50376 8128 50440 8132
rect 50456 8188 50520 8192
rect 50456 8132 50460 8188
rect 50460 8132 50516 8188
rect 50516 8132 50520 8188
rect 50456 8128 50520 8132
rect 50536 8188 50600 8192
rect 50536 8132 50540 8188
rect 50540 8132 50596 8188
rect 50596 8132 50600 8188
rect 50536 8128 50600 8132
rect 81016 8188 81080 8192
rect 81016 8132 81020 8188
rect 81020 8132 81076 8188
rect 81076 8132 81080 8188
rect 81016 8128 81080 8132
rect 81096 8188 81160 8192
rect 81096 8132 81100 8188
rect 81100 8132 81156 8188
rect 81156 8132 81160 8188
rect 81096 8128 81160 8132
rect 81176 8188 81240 8192
rect 81176 8132 81180 8188
rect 81180 8132 81236 8188
rect 81236 8132 81240 8188
rect 81176 8128 81240 8132
rect 81256 8188 81320 8192
rect 81256 8132 81260 8188
rect 81260 8132 81316 8188
rect 81316 8132 81320 8188
rect 81256 8128 81320 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 65656 7644 65720 7648
rect 65656 7588 65660 7644
rect 65660 7588 65716 7644
rect 65716 7588 65720 7644
rect 65656 7584 65720 7588
rect 65736 7644 65800 7648
rect 65736 7588 65740 7644
rect 65740 7588 65796 7644
rect 65796 7588 65800 7644
rect 65736 7584 65800 7588
rect 65816 7644 65880 7648
rect 65816 7588 65820 7644
rect 65820 7588 65876 7644
rect 65876 7588 65880 7644
rect 65816 7584 65880 7588
rect 65896 7644 65960 7648
rect 65896 7588 65900 7644
rect 65900 7588 65956 7644
rect 65956 7588 65960 7644
rect 65896 7584 65960 7588
rect 96376 7644 96440 7648
rect 96376 7588 96380 7644
rect 96380 7588 96436 7644
rect 96436 7588 96440 7644
rect 96376 7584 96440 7588
rect 96456 7644 96520 7648
rect 96456 7588 96460 7644
rect 96460 7588 96516 7644
rect 96516 7588 96520 7644
rect 96456 7584 96520 7588
rect 96536 7644 96600 7648
rect 96536 7588 96540 7644
rect 96540 7588 96596 7644
rect 96596 7588 96600 7644
rect 96536 7584 96600 7588
rect 96616 7644 96680 7648
rect 96616 7588 96620 7644
rect 96620 7588 96676 7644
rect 96676 7588 96680 7644
rect 96616 7584 96680 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 50296 7100 50360 7104
rect 50296 7044 50300 7100
rect 50300 7044 50356 7100
rect 50356 7044 50360 7100
rect 50296 7040 50360 7044
rect 50376 7100 50440 7104
rect 50376 7044 50380 7100
rect 50380 7044 50436 7100
rect 50436 7044 50440 7100
rect 50376 7040 50440 7044
rect 50456 7100 50520 7104
rect 50456 7044 50460 7100
rect 50460 7044 50516 7100
rect 50516 7044 50520 7100
rect 50456 7040 50520 7044
rect 50536 7100 50600 7104
rect 50536 7044 50540 7100
rect 50540 7044 50596 7100
rect 50596 7044 50600 7100
rect 50536 7040 50600 7044
rect 81016 7100 81080 7104
rect 81016 7044 81020 7100
rect 81020 7044 81076 7100
rect 81076 7044 81080 7100
rect 81016 7040 81080 7044
rect 81096 7100 81160 7104
rect 81096 7044 81100 7100
rect 81100 7044 81156 7100
rect 81156 7044 81160 7100
rect 81096 7040 81160 7044
rect 81176 7100 81240 7104
rect 81176 7044 81180 7100
rect 81180 7044 81236 7100
rect 81236 7044 81240 7100
rect 81176 7040 81240 7044
rect 81256 7100 81320 7104
rect 81256 7044 81260 7100
rect 81260 7044 81316 7100
rect 81316 7044 81320 7100
rect 81256 7040 81320 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 65656 6556 65720 6560
rect 65656 6500 65660 6556
rect 65660 6500 65716 6556
rect 65716 6500 65720 6556
rect 65656 6496 65720 6500
rect 65736 6556 65800 6560
rect 65736 6500 65740 6556
rect 65740 6500 65796 6556
rect 65796 6500 65800 6556
rect 65736 6496 65800 6500
rect 65816 6556 65880 6560
rect 65816 6500 65820 6556
rect 65820 6500 65876 6556
rect 65876 6500 65880 6556
rect 65816 6496 65880 6500
rect 65896 6556 65960 6560
rect 65896 6500 65900 6556
rect 65900 6500 65956 6556
rect 65956 6500 65960 6556
rect 65896 6496 65960 6500
rect 96376 6556 96440 6560
rect 96376 6500 96380 6556
rect 96380 6500 96436 6556
rect 96436 6500 96440 6556
rect 96376 6496 96440 6500
rect 96456 6556 96520 6560
rect 96456 6500 96460 6556
rect 96460 6500 96516 6556
rect 96516 6500 96520 6556
rect 96456 6496 96520 6500
rect 96536 6556 96600 6560
rect 96536 6500 96540 6556
rect 96540 6500 96596 6556
rect 96596 6500 96600 6556
rect 96536 6496 96600 6500
rect 96616 6556 96680 6560
rect 96616 6500 96620 6556
rect 96620 6500 96676 6556
rect 96676 6500 96680 6556
rect 96616 6496 96680 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 50296 6012 50360 6016
rect 50296 5956 50300 6012
rect 50300 5956 50356 6012
rect 50356 5956 50360 6012
rect 50296 5952 50360 5956
rect 50376 6012 50440 6016
rect 50376 5956 50380 6012
rect 50380 5956 50436 6012
rect 50436 5956 50440 6012
rect 50376 5952 50440 5956
rect 50456 6012 50520 6016
rect 50456 5956 50460 6012
rect 50460 5956 50516 6012
rect 50516 5956 50520 6012
rect 50456 5952 50520 5956
rect 50536 6012 50600 6016
rect 50536 5956 50540 6012
rect 50540 5956 50596 6012
rect 50596 5956 50600 6012
rect 50536 5952 50600 5956
rect 81016 6012 81080 6016
rect 81016 5956 81020 6012
rect 81020 5956 81076 6012
rect 81076 5956 81080 6012
rect 81016 5952 81080 5956
rect 81096 6012 81160 6016
rect 81096 5956 81100 6012
rect 81100 5956 81156 6012
rect 81156 5956 81160 6012
rect 81096 5952 81160 5956
rect 81176 6012 81240 6016
rect 81176 5956 81180 6012
rect 81180 5956 81236 6012
rect 81236 5956 81240 6012
rect 81176 5952 81240 5956
rect 81256 6012 81320 6016
rect 81256 5956 81260 6012
rect 81260 5956 81316 6012
rect 81316 5956 81320 6012
rect 81256 5952 81320 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 65656 5468 65720 5472
rect 65656 5412 65660 5468
rect 65660 5412 65716 5468
rect 65716 5412 65720 5468
rect 65656 5408 65720 5412
rect 65736 5468 65800 5472
rect 65736 5412 65740 5468
rect 65740 5412 65796 5468
rect 65796 5412 65800 5468
rect 65736 5408 65800 5412
rect 65816 5468 65880 5472
rect 65816 5412 65820 5468
rect 65820 5412 65876 5468
rect 65876 5412 65880 5468
rect 65816 5408 65880 5412
rect 65896 5468 65960 5472
rect 65896 5412 65900 5468
rect 65900 5412 65956 5468
rect 65956 5412 65960 5468
rect 65896 5408 65960 5412
rect 96376 5468 96440 5472
rect 96376 5412 96380 5468
rect 96380 5412 96436 5468
rect 96436 5412 96440 5468
rect 96376 5408 96440 5412
rect 96456 5468 96520 5472
rect 96456 5412 96460 5468
rect 96460 5412 96516 5468
rect 96516 5412 96520 5468
rect 96456 5408 96520 5412
rect 96536 5468 96600 5472
rect 96536 5412 96540 5468
rect 96540 5412 96596 5468
rect 96596 5412 96600 5468
rect 96536 5408 96600 5412
rect 96616 5468 96680 5472
rect 96616 5412 96620 5468
rect 96620 5412 96676 5468
rect 96676 5412 96680 5468
rect 96616 5408 96680 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 50296 4924 50360 4928
rect 50296 4868 50300 4924
rect 50300 4868 50356 4924
rect 50356 4868 50360 4924
rect 50296 4864 50360 4868
rect 50376 4924 50440 4928
rect 50376 4868 50380 4924
rect 50380 4868 50436 4924
rect 50436 4868 50440 4924
rect 50376 4864 50440 4868
rect 50456 4924 50520 4928
rect 50456 4868 50460 4924
rect 50460 4868 50516 4924
rect 50516 4868 50520 4924
rect 50456 4864 50520 4868
rect 50536 4924 50600 4928
rect 50536 4868 50540 4924
rect 50540 4868 50596 4924
rect 50596 4868 50600 4924
rect 50536 4864 50600 4868
rect 81016 4924 81080 4928
rect 81016 4868 81020 4924
rect 81020 4868 81076 4924
rect 81076 4868 81080 4924
rect 81016 4864 81080 4868
rect 81096 4924 81160 4928
rect 81096 4868 81100 4924
rect 81100 4868 81156 4924
rect 81156 4868 81160 4924
rect 81096 4864 81160 4868
rect 81176 4924 81240 4928
rect 81176 4868 81180 4924
rect 81180 4868 81236 4924
rect 81236 4868 81240 4924
rect 81176 4864 81240 4868
rect 81256 4924 81320 4928
rect 81256 4868 81260 4924
rect 81260 4868 81316 4924
rect 81316 4868 81320 4924
rect 81256 4864 81320 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 65656 4380 65720 4384
rect 65656 4324 65660 4380
rect 65660 4324 65716 4380
rect 65716 4324 65720 4380
rect 65656 4320 65720 4324
rect 65736 4380 65800 4384
rect 65736 4324 65740 4380
rect 65740 4324 65796 4380
rect 65796 4324 65800 4380
rect 65736 4320 65800 4324
rect 65816 4380 65880 4384
rect 65816 4324 65820 4380
rect 65820 4324 65876 4380
rect 65876 4324 65880 4380
rect 65816 4320 65880 4324
rect 65896 4380 65960 4384
rect 65896 4324 65900 4380
rect 65900 4324 65956 4380
rect 65956 4324 65960 4380
rect 65896 4320 65960 4324
rect 96376 4380 96440 4384
rect 96376 4324 96380 4380
rect 96380 4324 96436 4380
rect 96436 4324 96440 4380
rect 96376 4320 96440 4324
rect 96456 4380 96520 4384
rect 96456 4324 96460 4380
rect 96460 4324 96516 4380
rect 96516 4324 96520 4380
rect 96456 4320 96520 4324
rect 96536 4380 96600 4384
rect 96536 4324 96540 4380
rect 96540 4324 96596 4380
rect 96596 4324 96600 4380
rect 96536 4320 96600 4324
rect 96616 4380 96680 4384
rect 96616 4324 96620 4380
rect 96620 4324 96676 4380
rect 96676 4324 96680 4380
rect 96616 4320 96680 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 50296 3836 50360 3840
rect 50296 3780 50300 3836
rect 50300 3780 50356 3836
rect 50356 3780 50360 3836
rect 50296 3776 50360 3780
rect 50376 3836 50440 3840
rect 50376 3780 50380 3836
rect 50380 3780 50436 3836
rect 50436 3780 50440 3836
rect 50376 3776 50440 3780
rect 50456 3836 50520 3840
rect 50456 3780 50460 3836
rect 50460 3780 50516 3836
rect 50516 3780 50520 3836
rect 50456 3776 50520 3780
rect 50536 3836 50600 3840
rect 50536 3780 50540 3836
rect 50540 3780 50596 3836
rect 50596 3780 50600 3836
rect 50536 3776 50600 3780
rect 81016 3836 81080 3840
rect 81016 3780 81020 3836
rect 81020 3780 81076 3836
rect 81076 3780 81080 3836
rect 81016 3776 81080 3780
rect 81096 3836 81160 3840
rect 81096 3780 81100 3836
rect 81100 3780 81156 3836
rect 81156 3780 81160 3836
rect 81096 3776 81160 3780
rect 81176 3836 81240 3840
rect 81176 3780 81180 3836
rect 81180 3780 81236 3836
rect 81236 3780 81240 3836
rect 81176 3776 81240 3780
rect 81256 3836 81320 3840
rect 81256 3780 81260 3836
rect 81260 3780 81316 3836
rect 81316 3780 81320 3836
rect 81256 3776 81320 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 65656 3292 65720 3296
rect 65656 3236 65660 3292
rect 65660 3236 65716 3292
rect 65716 3236 65720 3292
rect 65656 3232 65720 3236
rect 65736 3292 65800 3296
rect 65736 3236 65740 3292
rect 65740 3236 65796 3292
rect 65796 3236 65800 3292
rect 65736 3232 65800 3236
rect 65816 3292 65880 3296
rect 65816 3236 65820 3292
rect 65820 3236 65876 3292
rect 65876 3236 65880 3292
rect 65816 3232 65880 3236
rect 65896 3292 65960 3296
rect 65896 3236 65900 3292
rect 65900 3236 65956 3292
rect 65956 3236 65960 3292
rect 65896 3232 65960 3236
rect 96376 3292 96440 3296
rect 96376 3236 96380 3292
rect 96380 3236 96436 3292
rect 96436 3236 96440 3292
rect 96376 3232 96440 3236
rect 96456 3292 96520 3296
rect 96456 3236 96460 3292
rect 96460 3236 96516 3292
rect 96516 3236 96520 3292
rect 96456 3232 96520 3236
rect 96536 3292 96600 3296
rect 96536 3236 96540 3292
rect 96540 3236 96596 3292
rect 96596 3236 96600 3292
rect 96536 3232 96600 3236
rect 96616 3292 96680 3296
rect 96616 3236 96620 3292
rect 96620 3236 96676 3292
rect 96676 3236 96680 3292
rect 96616 3232 96680 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 50296 2748 50360 2752
rect 50296 2692 50300 2748
rect 50300 2692 50356 2748
rect 50356 2692 50360 2748
rect 50296 2688 50360 2692
rect 50376 2748 50440 2752
rect 50376 2692 50380 2748
rect 50380 2692 50436 2748
rect 50436 2692 50440 2748
rect 50376 2688 50440 2692
rect 50456 2748 50520 2752
rect 50456 2692 50460 2748
rect 50460 2692 50516 2748
rect 50516 2692 50520 2748
rect 50456 2688 50520 2692
rect 50536 2748 50600 2752
rect 50536 2692 50540 2748
rect 50540 2692 50596 2748
rect 50596 2692 50600 2748
rect 50536 2688 50600 2692
rect 81016 2748 81080 2752
rect 81016 2692 81020 2748
rect 81020 2692 81076 2748
rect 81076 2692 81080 2748
rect 81016 2688 81080 2692
rect 81096 2748 81160 2752
rect 81096 2692 81100 2748
rect 81100 2692 81156 2748
rect 81156 2692 81160 2748
rect 81096 2688 81160 2692
rect 81176 2748 81240 2752
rect 81176 2692 81180 2748
rect 81180 2692 81236 2748
rect 81236 2692 81240 2748
rect 81176 2688 81240 2692
rect 81256 2748 81320 2752
rect 81256 2692 81260 2748
rect 81260 2692 81316 2748
rect 81316 2692 81320 2748
rect 81256 2688 81320 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
rect 65656 2204 65720 2208
rect 65656 2148 65660 2204
rect 65660 2148 65716 2204
rect 65716 2148 65720 2204
rect 65656 2144 65720 2148
rect 65736 2204 65800 2208
rect 65736 2148 65740 2204
rect 65740 2148 65796 2204
rect 65796 2148 65800 2204
rect 65736 2144 65800 2148
rect 65816 2204 65880 2208
rect 65816 2148 65820 2204
rect 65820 2148 65876 2204
rect 65876 2148 65880 2204
rect 65816 2144 65880 2148
rect 65896 2204 65960 2208
rect 65896 2148 65900 2204
rect 65900 2148 65956 2204
rect 65956 2148 65960 2204
rect 65896 2144 65960 2148
rect 96376 2204 96440 2208
rect 96376 2148 96380 2204
rect 96380 2148 96436 2204
rect 96436 2148 96440 2204
rect 96376 2144 96440 2148
rect 96456 2204 96520 2208
rect 96456 2148 96460 2204
rect 96460 2148 96516 2204
rect 96516 2148 96520 2204
rect 96456 2144 96520 2148
rect 96536 2204 96600 2208
rect 96536 2148 96540 2204
rect 96540 2148 96596 2204
rect 96596 2148 96600 2204
rect 96536 2144 96600 2148
rect 96616 2204 96680 2208
rect 96616 2148 96620 2204
rect 96620 2148 96676 2204
rect 96676 2148 96680 2204
rect 96616 2144 96680 2148
<< metal4 >>
rect 4208 96864 4528 97424
rect 19568 97408 19888 97424
rect 4208 96800 4216 96864
rect 4280 96800 4296 96864
rect 4360 96800 4376 96864
rect 4440 96800 4456 96864
rect 4520 96800 4528 96864
rect 4208 95776 4528 96800
rect 4208 95712 4216 95776
rect 4280 95712 4296 95776
rect 4360 95712 4376 95776
rect 4440 95712 4456 95776
rect 4520 95712 4528 95776
rect 4208 94688 4528 95712
rect 4208 94624 4216 94688
rect 4280 94624 4296 94688
rect 4360 94624 4376 94688
rect 4440 94624 4456 94688
rect 4520 94624 4528 94688
rect 4208 93600 4528 94624
rect 4208 93536 4216 93600
rect 4280 93536 4296 93600
rect 4360 93536 4376 93600
rect 4440 93536 4456 93600
rect 4520 93536 4528 93600
rect 4208 92512 4528 93536
rect 4208 92448 4216 92512
rect 4280 92448 4296 92512
rect 4360 92448 4376 92512
rect 4440 92448 4456 92512
rect 4520 92448 4528 92512
rect 4208 91424 4528 92448
rect 4208 91360 4216 91424
rect 4280 91360 4296 91424
rect 4360 91360 4376 91424
rect 4440 91360 4456 91424
rect 4520 91360 4528 91424
rect 4208 90336 4528 91360
rect 4208 90272 4216 90336
rect 4280 90272 4296 90336
rect 4360 90272 4376 90336
rect 4440 90272 4456 90336
rect 4520 90272 4528 90336
rect 4208 89248 4528 90272
rect 4208 89184 4216 89248
rect 4280 89184 4296 89248
rect 4360 89184 4376 89248
rect 4440 89184 4456 89248
rect 4520 89184 4528 89248
rect 4208 88160 4528 89184
rect 4208 88096 4216 88160
rect 4280 88096 4296 88160
rect 4360 88096 4376 88160
rect 4440 88096 4456 88160
rect 4520 88096 4528 88160
rect 4208 87072 4528 88096
rect 4208 87008 4216 87072
rect 4280 87008 4296 87072
rect 4360 87008 4376 87072
rect 4440 87008 4456 87072
rect 4520 87008 4528 87072
rect 4208 85984 4528 87008
rect 4208 85920 4216 85984
rect 4280 85920 4296 85984
rect 4360 85920 4376 85984
rect 4440 85920 4456 85984
rect 4520 85920 4528 85984
rect 4208 84896 4528 85920
rect 4208 84832 4216 84896
rect 4280 84832 4296 84896
rect 4360 84832 4376 84896
rect 4440 84832 4456 84896
rect 4520 84832 4528 84896
rect 4208 83808 4528 84832
rect 4208 83744 4216 83808
rect 4280 83744 4296 83808
rect 4360 83744 4376 83808
rect 4440 83744 4456 83808
rect 4520 83744 4528 83808
rect 4208 82720 4528 83744
rect 4208 82656 4216 82720
rect 4280 82656 4296 82720
rect 4360 82656 4376 82720
rect 4440 82656 4456 82720
rect 4520 82656 4528 82720
rect 4208 81632 4528 82656
rect 4208 81568 4216 81632
rect 4280 81568 4296 81632
rect 4360 81568 4376 81632
rect 4440 81568 4456 81632
rect 4520 81568 4528 81632
rect 4208 80544 4528 81568
rect 4208 80480 4216 80544
rect 4280 80480 4296 80544
rect 4360 80480 4376 80544
rect 4440 80480 4456 80544
rect 4520 80480 4528 80544
rect 4208 79456 4528 80480
rect 4208 79392 4216 79456
rect 4280 79392 4296 79456
rect 4360 79392 4376 79456
rect 4440 79392 4456 79456
rect 4520 79392 4528 79456
rect 4208 78368 4528 79392
rect 4208 78304 4216 78368
rect 4280 78304 4296 78368
rect 4360 78304 4376 78368
rect 4440 78304 4456 78368
rect 4520 78304 4528 78368
rect 4208 77280 4528 78304
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 76192 4528 77216
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 75104 4528 76128
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 74016 4528 75040
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 72928 4528 73952
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 71840 4528 72864
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 70752 4528 71776
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 69664 4528 70688
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 68576 4528 69600
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 67488 4528 68512
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 66400 4528 67424
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 65312 4528 66336
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 64224 4528 65248
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 63136 4528 64160
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 62048 4528 63072
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 60960 4528 61984
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 59872 4528 60896
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 58784 4528 59808
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 57696 4528 58720
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 56608 4528 57632
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 55520 4528 56544
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 54432 4528 55456
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 53344 4528 54368
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 52256 4528 53280
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 51168 4528 52192
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 50080 4528 51104
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 48992 4528 50016
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 47904 4528 48928
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4868 2176 5188 97376
rect 5528 2176 5848 97376
rect 6188 2176 6508 97376
rect 19568 97344 19576 97408
rect 19640 97344 19656 97408
rect 19720 97344 19736 97408
rect 19800 97344 19816 97408
rect 19880 97344 19888 97408
rect 19568 96320 19888 97344
rect 19568 96256 19576 96320
rect 19640 96256 19656 96320
rect 19720 96256 19736 96320
rect 19800 96256 19816 96320
rect 19880 96256 19888 96320
rect 19568 95232 19888 96256
rect 19568 95168 19576 95232
rect 19640 95168 19656 95232
rect 19720 95168 19736 95232
rect 19800 95168 19816 95232
rect 19880 95168 19888 95232
rect 19568 94144 19888 95168
rect 19568 94080 19576 94144
rect 19640 94080 19656 94144
rect 19720 94080 19736 94144
rect 19800 94080 19816 94144
rect 19880 94080 19888 94144
rect 19568 93056 19888 94080
rect 19568 92992 19576 93056
rect 19640 92992 19656 93056
rect 19720 92992 19736 93056
rect 19800 92992 19816 93056
rect 19880 92992 19888 93056
rect 19568 91968 19888 92992
rect 19568 91904 19576 91968
rect 19640 91904 19656 91968
rect 19720 91904 19736 91968
rect 19800 91904 19816 91968
rect 19880 91904 19888 91968
rect 19568 90880 19888 91904
rect 19568 90816 19576 90880
rect 19640 90816 19656 90880
rect 19720 90816 19736 90880
rect 19800 90816 19816 90880
rect 19880 90816 19888 90880
rect 19568 89792 19888 90816
rect 19568 89728 19576 89792
rect 19640 89728 19656 89792
rect 19720 89728 19736 89792
rect 19800 89728 19816 89792
rect 19880 89728 19888 89792
rect 19568 88704 19888 89728
rect 19568 88640 19576 88704
rect 19640 88640 19656 88704
rect 19720 88640 19736 88704
rect 19800 88640 19816 88704
rect 19880 88640 19888 88704
rect 19568 87616 19888 88640
rect 19568 87552 19576 87616
rect 19640 87552 19656 87616
rect 19720 87552 19736 87616
rect 19800 87552 19816 87616
rect 19880 87552 19888 87616
rect 19568 86528 19888 87552
rect 19568 86464 19576 86528
rect 19640 86464 19656 86528
rect 19720 86464 19736 86528
rect 19800 86464 19816 86528
rect 19880 86464 19888 86528
rect 19568 85440 19888 86464
rect 19568 85376 19576 85440
rect 19640 85376 19656 85440
rect 19720 85376 19736 85440
rect 19800 85376 19816 85440
rect 19880 85376 19888 85440
rect 19568 84352 19888 85376
rect 19568 84288 19576 84352
rect 19640 84288 19656 84352
rect 19720 84288 19736 84352
rect 19800 84288 19816 84352
rect 19880 84288 19888 84352
rect 19568 83264 19888 84288
rect 19568 83200 19576 83264
rect 19640 83200 19656 83264
rect 19720 83200 19736 83264
rect 19800 83200 19816 83264
rect 19880 83200 19888 83264
rect 19568 82176 19888 83200
rect 19568 82112 19576 82176
rect 19640 82112 19656 82176
rect 19720 82112 19736 82176
rect 19800 82112 19816 82176
rect 19880 82112 19888 82176
rect 19568 81088 19888 82112
rect 19568 81024 19576 81088
rect 19640 81024 19656 81088
rect 19720 81024 19736 81088
rect 19800 81024 19816 81088
rect 19880 81024 19888 81088
rect 19568 80000 19888 81024
rect 19568 79936 19576 80000
rect 19640 79936 19656 80000
rect 19720 79936 19736 80000
rect 19800 79936 19816 80000
rect 19880 79936 19888 80000
rect 19568 78912 19888 79936
rect 19568 78848 19576 78912
rect 19640 78848 19656 78912
rect 19720 78848 19736 78912
rect 19800 78848 19816 78912
rect 19880 78848 19888 78912
rect 19568 77824 19888 78848
rect 19568 77760 19576 77824
rect 19640 77760 19656 77824
rect 19720 77760 19736 77824
rect 19800 77760 19816 77824
rect 19880 77760 19888 77824
rect 19568 76736 19888 77760
rect 19568 76672 19576 76736
rect 19640 76672 19656 76736
rect 19720 76672 19736 76736
rect 19800 76672 19816 76736
rect 19880 76672 19888 76736
rect 19568 75648 19888 76672
rect 19568 75584 19576 75648
rect 19640 75584 19656 75648
rect 19720 75584 19736 75648
rect 19800 75584 19816 75648
rect 19880 75584 19888 75648
rect 19568 74560 19888 75584
rect 19568 74496 19576 74560
rect 19640 74496 19656 74560
rect 19720 74496 19736 74560
rect 19800 74496 19816 74560
rect 19880 74496 19888 74560
rect 19568 73472 19888 74496
rect 19568 73408 19576 73472
rect 19640 73408 19656 73472
rect 19720 73408 19736 73472
rect 19800 73408 19816 73472
rect 19880 73408 19888 73472
rect 19568 72384 19888 73408
rect 19568 72320 19576 72384
rect 19640 72320 19656 72384
rect 19720 72320 19736 72384
rect 19800 72320 19816 72384
rect 19880 72320 19888 72384
rect 19568 71296 19888 72320
rect 19568 71232 19576 71296
rect 19640 71232 19656 71296
rect 19720 71232 19736 71296
rect 19800 71232 19816 71296
rect 19880 71232 19888 71296
rect 19568 70208 19888 71232
rect 19568 70144 19576 70208
rect 19640 70144 19656 70208
rect 19720 70144 19736 70208
rect 19800 70144 19816 70208
rect 19880 70144 19888 70208
rect 19568 69120 19888 70144
rect 19568 69056 19576 69120
rect 19640 69056 19656 69120
rect 19720 69056 19736 69120
rect 19800 69056 19816 69120
rect 19880 69056 19888 69120
rect 19568 68032 19888 69056
rect 19568 67968 19576 68032
rect 19640 67968 19656 68032
rect 19720 67968 19736 68032
rect 19800 67968 19816 68032
rect 19880 67968 19888 68032
rect 19568 66944 19888 67968
rect 19568 66880 19576 66944
rect 19640 66880 19656 66944
rect 19720 66880 19736 66944
rect 19800 66880 19816 66944
rect 19880 66880 19888 66944
rect 19568 65856 19888 66880
rect 19568 65792 19576 65856
rect 19640 65792 19656 65856
rect 19720 65792 19736 65856
rect 19800 65792 19816 65856
rect 19880 65792 19888 65856
rect 19568 64768 19888 65792
rect 19568 64704 19576 64768
rect 19640 64704 19656 64768
rect 19720 64704 19736 64768
rect 19800 64704 19816 64768
rect 19880 64704 19888 64768
rect 19568 63680 19888 64704
rect 19568 63616 19576 63680
rect 19640 63616 19656 63680
rect 19720 63616 19736 63680
rect 19800 63616 19816 63680
rect 19880 63616 19888 63680
rect 19568 62592 19888 63616
rect 19568 62528 19576 62592
rect 19640 62528 19656 62592
rect 19720 62528 19736 62592
rect 19800 62528 19816 62592
rect 19880 62528 19888 62592
rect 19568 61504 19888 62528
rect 19568 61440 19576 61504
rect 19640 61440 19656 61504
rect 19720 61440 19736 61504
rect 19800 61440 19816 61504
rect 19880 61440 19888 61504
rect 19568 60416 19888 61440
rect 19568 60352 19576 60416
rect 19640 60352 19656 60416
rect 19720 60352 19736 60416
rect 19800 60352 19816 60416
rect 19880 60352 19888 60416
rect 19568 59328 19888 60352
rect 19568 59264 19576 59328
rect 19640 59264 19656 59328
rect 19720 59264 19736 59328
rect 19800 59264 19816 59328
rect 19880 59264 19888 59328
rect 19568 58240 19888 59264
rect 19568 58176 19576 58240
rect 19640 58176 19656 58240
rect 19720 58176 19736 58240
rect 19800 58176 19816 58240
rect 19880 58176 19888 58240
rect 19568 57152 19888 58176
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 56064 19888 57088
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 54976 19888 56000
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 53888 19888 54912
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 52800 19888 53824
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 51712 19888 52736
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 50624 19888 51648
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 49536 19888 50560
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 48448 19888 49472
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 47360 19888 48384
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 4208 2128 4528 2144
rect 19568 2128 19888 2688
rect 20228 2176 20548 97376
rect 20888 2176 21208 97376
rect 21548 2176 21868 97376
rect 34928 96864 35248 97424
rect 50288 97408 50608 97424
rect 34928 96800 34936 96864
rect 35000 96800 35016 96864
rect 35080 96800 35096 96864
rect 35160 96800 35176 96864
rect 35240 96800 35248 96864
rect 34928 95776 35248 96800
rect 34928 95712 34936 95776
rect 35000 95712 35016 95776
rect 35080 95712 35096 95776
rect 35160 95712 35176 95776
rect 35240 95712 35248 95776
rect 34928 94688 35248 95712
rect 34928 94624 34936 94688
rect 35000 94624 35016 94688
rect 35080 94624 35096 94688
rect 35160 94624 35176 94688
rect 35240 94624 35248 94688
rect 34928 93600 35248 94624
rect 34928 93536 34936 93600
rect 35000 93536 35016 93600
rect 35080 93536 35096 93600
rect 35160 93536 35176 93600
rect 35240 93536 35248 93600
rect 34928 92512 35248 93536
rect 34928 92448 34936 92512
rect 35000 92448 35016 92512
rect 35080 92448 35096 92512
rect 35160 92448 35176 92512
rect 35240 92448 35248 92512
rect 34928 91424 35248 92448
rect 34928 91360 34936 91424
rect 35000 91360 35016 91424
rect 35080 91360 35096 91424
rect 35160 91360 35176 91424
rect 35240 91360 35248 91424
rect 34928 90336 35248 91360
rect 34928 90272 34936 90336
rect 35000 90272 35016 90336
rect 35080 90272 35096 90336
rect 35160 90272 35176 90336
rect 35240 90272 35248 90336
rect 34928 89248 35248 90272
rect 34928 89184 34936 89248
rect 35000 89184 35016 89248
rect 35080 89184 35096 89248
rect 35160 89184 35176 89248
rect 35240 89184 35248 89248
rect 34928 88160 35248 89184
rect 34928 88096 34936 88160
rect 35000 88096 35016 88160
rect 35080 88096 35096 88160
rect 35160 88096 35176 88160
rect 35240 88096 35248 88160
rect 34928 87072 35248 88096
rect 34928 87008 34936 87072
rect 35000 87008 35016 87072
rect 35080 87008 35096 87072
rect 35160 87008 35176 87072
rect 35240 87008 35248 87072
rect 34928 85984 35248 87008
rect 34928 85920 34936 85984
rect 35000 85920 35016 85984
rect 35080 85920 35096 85984
rect 35160 85920 35176 85984
rect 35240 85920 35248 85984
rect 34928 84896 35248 85920
rect 34928 84832 34936 84896
rect 35000 84832 35016 84896
rect 35080 84832 35096 84896
rect 35160 84832 35176 84896
rect 35240 84832 35248 84896
rect 34928 83808 35248 84832
rect 34928 83744 34936 83808
rect 35000 83744 35016 83808
rect 35080 83744 35096 83808
rect 35160 83744 35176 83808
rect 35240 83744 35248 83808
rect 34928 82720 35248 83744
rect 34928 82656 34936 82720
rect 35000 82656 35016 82720
rect 35080 82656 35096 82720
rect 35160 82656 35176 82720
rect 35240 82656 35248 82720
rect 34928 81632 35248 82656
rect 34928 81568 34936 81632
rect 35000 81568 35016 81632
rect 35080 81568 35096 81632
rect 35160 81568 35176 81632
rect 35240 81568 35248 81632
rect 34928 80544 35248 81568
rect 34928 80480 34936 80544
rect 35000 80480 35016 80544
rect 35080 80480 35096 80544
rect 35160 80480 35176 80544
rect 35240 80480 35248 80544
rect 34928 79456 35248 80480
rect 34928 79392 34936 79456
rect 35000 79392 35016 79456
rect 35080 79392 35096 79456
rect 35160 79392 35176 79456
rect 35240 79392 35248 79456
rect 34928 78368 35248 79392
rect 34928 78304 34936 78368
rect 35000 78304 35016 78368
rect 35080 78304 35096 78368
rect 35160 78304 35176 78368
rect 35240 78304 35248 78368
rect 34928 77280 35248 78304
rect 34928 77216 34936 77280
rect 35000 77216 35016 77280
rect 35080 77216 35096 77280
rect 35160 77216 35176 77280
rect 35240 77216 35248 77280
rect 34928 76192 35248 77216
rect 34928 76128 34936 76192
rect 35000 76128 35016 76192
rect 35080 76128 35096 76192
rect 35160 76128 35176 76192
rect 35240 76128 35248 76192
rect 34928 75104 35248 76128
rect 34928 75040 34936 75104
rect 35000 75040 35016 75104
rect 35080 75040 35096 75104
rect 35160 75040 35176 75104
rect 35240 75040 35248 75104
rect 34928 74016 35248 75040
rect 34928 73952 34936 74016
rect 35000 73952 35016 74016
rect 35080 73952 35096 74016
rect 35160 73952 35176 74016
rect 35240 73952 35248 74016
rect 34928 72928 35248 73952
rect 34928 72864 34936 72928
rect 35000 72864 35016 72928
rect 35080 72864 35096 72928
rect 35160 72864 35176 72928
rect 35240 72864 35248 72928
rect 34928 71840 35248 72864
rect 34928 71776 34936 71840
rect 35000 71776 35016 71840
rect 35080 71776 35096 71840
rect 35160 71776 35176 71840
rect 35240 71776 35248 71840
rect 34928 70752 35248 71776
rect 34928 70688 34936 70752
rect 35000 70688 35016 70752
rect 35080 70688 35096 70752
rect 35160 70688 35176 70752
rect 35240 70688 35248 70752
rect 34928 69664 35248 70688
rect 34928 69600 34936 69664
rect 35000 69600 35016 69664
rect 35080 69600 35096 69664
rect 35160 69600 35176 69664
rect 35240 69600 35248 69664
rect 34928 68576 35248 69600
rect 34928 68512 34936 68576
rect 35000 68512 35016 68576
rect 35080 68512 35096 68576
rect 35160 68512 35176 68576
rect 35240 68512 35248 68576
rect 34928 67488 35248 68512
rect 34928 67424 34936 67488
rect 35000 67424 35016 67488
rect 35080 67424 35096 67488
rect 35160 67424 35176 67488
rect 35240 67424 35248 67488
rect 34928 66400 35248 67424
rect 34928 66336 34936 66400
rect 35000 66336 35016 66400
rect 35080 66336 35096 66400
rect 35160 66336 35176 66400
rect 35240 66336 35248 66400
rect 34928 65312 35248 66336
rect 34928 65248 34936 65312
rect 35000 65248 35016 65312
rect 35080 65248 35096 65312
rect 35160 65248 35176 65312
rect 35240 65248 35248 65312
rect 34928 64224 35248 65248
rect 34928 64160 34936 64224
rect 35000 64160 35016 64224
rect 35080 64160 35096 64224
rect 35160 64160 35176 64224
rect 35240 64160 35248 64224
rect 34928 63136 35248 64160
rect 34928 63072 34936 63136
rect 35000 63072 35016 63136
rect 35080 63072 35096 63136
rect 35160 63072 35176 63136
rect 35240 63072 35248 63136
rect 34928 62048 35248 63072
rect 34928 61984 34936 62048
rect 35000 61984 35016 62048
rect 35080 61984 35096 62048
rect 35160 61984 35176 62048
rect 35240 61984 35248 62048
rect 34928 60960 35248 61984
rect 34928 60896 34936 60960
rect 35000 60896 35016 60960
rect 35080 60896 35096 60960
rect 35160 60896 35176 60960
rect 35240 60896 35248 60960
rect 34928 59872 35248 60896
rect 34928 59808 34936 59872
rect 35000 59808 35016 59872
rect 35080 59808 35096 59872
rect 35160 59808 35176 59872
rect 35240 59808 35248 59872
rect 34928 58784 35248 59808
rect 34928 58720 34936 58784
rect 35000 58720 35016 58784
rect 35080 58720 35096 58784
rect 35160 58720 35176 58784
rect 35240 58720 35248 58784
rect 34928 57696 35248 58720
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 56608 35248 57632
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 55520 35248 56544
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 54432 35248 55456
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 53344 35248 54368
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 52256 35248 53280
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 51168 35248 52192
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 50080 35248 51104
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 48992 35248 50016
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 47904 35248 48928
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 46816 35248 47840
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 35588 2176 35908 97376
rect 36248 2176 36568 97376
rect 36908 2176 37228 97376
rect 50288 97344 50296 97408
rect 50360 97344 50376 97408
rect 50440 97344 50456 97408
rect 50520 97344 50536 97408
rect 50600 97344 50608 97408
rect 50288 96320 50608 97344
rect 50288 96256 50296 96320
rect 50360 96256 50376 96320
rect 50440 96256 50456 96320
rect 50520 96256 50536 96320
rect 50600 96256 50608 96320
rect 50288 95232 50608 96256
rect 50288 95168 50296 95232
rect 50360 95168 50376 95232
rect 50440 95168 50456 95232
rect 50520 95168 50536 95232
rect 50600 95168 50608 95232
rect 50288 94144 50608 95168
rect 50288 94080 50296 94144
rect 50360 94080 50376 94144
rect 50440 94080 50456 94144
rect 50520 94080 50536 94144
rect 50600 94080 50608 94144
rect 50288 93056 50608 94080
rect 50288 92992 50296 93056
rect 50360 92992 50376 93056
rect 50440 92992 50456 93056
rect 50520 92992 50536 93056
rect 50600 92992 50608 93056
rect 50288 91968 50608 92992
rect 50288 91904 50296 91968
rect 50360 91904 50376 91968
rect 50440 91904 50456 91968
rect 50520 91904 50536 91968
rect 50600 91904 50608 91968
rect 50288 90880 50608 91904
rect 50288 90816 50296 90880
rect 50360 90816 50376 90880
rect 50440 90816 50456 90880
rect 50520 90816 50536 90880
rect 50600 90816 50608 90880
rect 50288 89792 50608 90816
rect 50288 89728 50296 89792
rect 50360 89728 50376 89792
rect 50440 89728 50456 89792
rect 50520 89728 50536 89792
rect 50600 89728 50608 89792
rect 50288 88704 50608 89728
rect 50288 88640 50296 88704
rect 50360 88640 50376 88704
rect 50440 88640 50456 88704
rect 50520 88640 50536 88704
rect 50600 88640 50608 88704
rect 50288 87616 50608 88640
rect 50288 87552 50296 87616
rect 50360 87552 50376 87616
rect 50440 87552 50456 87616
rect 50520 87552 50536 87616
rect 50600 87552 50608 87616
rect 50288 86528 50608 87552
rect 50288 86464 50296 86528
rect 50360 86464 50376 86528
rect 50440 86464 50456 86528
rect 50520 86464 50536 86528
rect 50600 86464 50608 86528
rect 50288 85440 50608 86464
rect 50288 85376 50296 85440
rect 50360 85376 50376 85440
rect 50440 85376 50456 85440
rect 50520 85376 50536 85440
rect 50600 85376 50608 85440
rect 50288 84352 50608 85376
rect 50288 84288 50296 84352
rect 50360 84288 50376 84352
rect 50440 84288 50456 84352
rect 50520 84288 50536 84352
rect 50600 84288 50608 84352
rect 50288 83264 50608 84288
rect 50288 83200 50296 83264
rect 50360 83200 50376 83264
rect 50440 83200 50456 83264
rect 50520 83200 50536 83264
rect 50600 83200 50608 83264
rect 50288 82176 50608 83200
rect 50288 82112 50296 82176
rect 50360 82112 50376 82176
rect 50440 82112 50456 82176
rect 50520 82112 50536 82176
rect 50600 82112 50608 82176
rect 50288 81088 50608 82112
rect 50288 81024 50296 81088
rect 50360 81024 50376 81088
rect 50440 81024 50456 81088
rect 50520 81024 50536 81088
rect 50600 81024 50608 81088
rect 50288 80000 50608 81024
rect 50288 79936 50296 80000
rect 50360 79936 50376 80000
rect 50440 79936 50456 80000
rect 50520 79936 50536 80000
rect 50600 79936 50608 80000
rect 50288 78912 50608 79936
rect 50288 78848 50296 78912
rect 50360 78848 50376 78912
rect 50440 78848 50456 78912
rect 50520 78848 50536 78912
rect 50600 78848 50608 78912
rect 50288 77824 50608 78848
rect 50288 77760 50296 77824
rect 50360 77760 50376 77824
rect 50440 77760 50456 77824
rect 50520 77760 50536 77824
rect 50600 77760 50608 77824
rect 50288 76736 50608 77760
rect 50288 76672 50296 76736
rect 50360 76672 50376 76736
rect 50440 76672 50456 76736
rect 50520 76672 50536 76736
rect 50600 76672 50608 76736
rect 50288 75648 50608 76672
rect 50288 75584 50296 75648
rect 50360 75584 50376 75648
rect 50440 75584 50456 75648
rect 50520 75584 50536 75648
rect 50600 75584 50608 75648
rect 50288 74560 50608 75584
rect 50288 74496 50296 74560
rect 50360 74496 50376 74560
rect 50440 74496 50456 74560
rect 50520 74496 50536 74560
rect 50600 74496 50608 74560
rect 50288 73472 50608 74496
rect 50288 73408 50296 73472
rect 50360 73408 50376 73472
rect 50440 73408 50456 73472
rect 50520 73408 50536 73472
rect 50600 73408 50608 73472
rect 50288 72384 50608 73408
rect 50288 72320 50296 72384
rect 50360 72320 50376 72384
rect 50440 72320 50456 72384
rect 50520 72320 50536 72384
rect 50600 72320 50608 72384
rect 50288 71296 50608 72320
rect 50288 71232 50296 71296
rect 50360 71232 50376 71296
rect 50440 71232 50456 71296
rect 50520 71232 50536 71296
rect 50600 71232 50608 71296
rect 50288 70208 50608 71232
rect 50288 70144 50296 70208
rect 50360 70144 50376 70208
rect 50440 70144 50456 70208
rect 50520 70144 50536 70208
rect 50600 70144 50608 70208
rect 50288 69120 50608 70144
rect 50288 69056 50296 69120
rect 50360 69056 50376 69120
rect 50440 69056 50456 69120
rect 50520 69056 50536 69120
rect 50600 69056 50608 69120
rect 50288 68032 50608 69056
rect 50288 67968 50296 68032
rect 50360 67968 50376 68032
rect 50440 67968 50456 68032
rect 50520 67968 50536 68032
rect 50600 67968 50608 68032
rect 50288 66944 50608 67968
rect 50288 66880 50296 66944
rect 50360 66880 50376 66944
rect 50440 66880 50456 66944
rect 50520 66880 50536 66944
rect 50600 66880 50608 66944
rect 50288 65856 50608 66880
rect 50288 65792 50296 65856
rect 50360 65792 50376 65856
rect 50440 65792 50456 65856
rect 50520 65792 50536 65856
rect 50600 65792 50608 65856
rect 50288 64768 50608 65792
rect 50288 64704 50296 64768
rect 50360 64704 50376 64768
rect 50440 64704 50456 64768
rect 50520 64704 50536 64768
rect 50600 64704 50608 64768
rect 50288 63680 50608 64704
rect 50288 63616 50296 63680
rect 50360 63616 50376 63680
rect 50440 63616 50456 63680
rect 50520 63616 50536 63680
rect 50600 63616 50608 63680
rect 50288 62592 50608 63616
rect 50288 62528 50296 62592
rect 50360 62528 50376 62592
rect 50440 62528 50456 62592
rect 50520 62528 50536 62592
rect 50600 62528 50608 62592
rect 50288 61504 50608 62528
rect 50288 61440 50296 61504
rect 50360 61440 50376 61504
rect 50440 61440 50456 61504
rect 50520 61440 50536 61504
rect 50600 61440 50608 61504
rect 50288 60416 50608 61440
rect 50288 60352 50296 60416
rect 50360 60352 50376 60416
rect 50440 60352 50456 60416
rect 50520 60352 50536 60416
rect 50600 60352 50608 60416
rect 50288 59328 50608 60352
rect 50288 59264 50296 59328
rect 50360 59264 50376 59328
rect 50440 59264 50456 59328
rect 50520 59264 50536 59328
rect 50600 59264 50608 59328
rect 50288 58240 50608 59264
rect 50288 58176 50296 58240
rect 50360 58176 50376 58240
rect 50440 58176 50456 58240
rect 50520 58176 50536 58240
rect 50600 58176 50608 58240
rect 50288 57152 50608 58176
rect 50288 57088 50296 57152
rect 50360 57088 50376 57152
rect 50440 57088 50456 57152
rect 50520 57088 50536 57152
rect 50600 57088 50608 57152
rect 50288 56064 50608 57088
rect 50288 56000 50296 56064
rect 50360 56000 50376 56064
rect 50440 56000 50456 56064
rect 50520 56000 50536 56064
rect 50600 56000 50608 56064
rect 50288 54976 50608 56000
rect 50288 54912 50296 54976
rect 50360 54912 50376 54976
rect 50440 54912 50456 54976
rect 50520 54912 50536 54976
rect 50600 54912 50608 54976
rect 50288 53888 50608 54912
rect 50288 53824 50296 53888
rect 50360 53824 50376 53888
rect 50440 53824 50456 53888
rect 50520 53824 50536 53888
rect 50600 53824 50608 53888
rect 50288 52800 50608 53824
rect 50288 52736 50296 52800
rect 50360 52736 50376 52800
rect 50440 52736 50456 52800
rect 50520 52736 50536 52800
rect 50600 52736 50608 52800
rect 50288 51712 50608 52736
rect 50288 51648 50296 51712
rect 50360 51648 50376 51712
rect 50440 51648 50456 51712
rect 50520 51648 50536 51712
rect 50600 51648 50608 51712
rect 50288 50624 50608 51648
rect 50288 50560 50296 50624
rect 50360 50560 50376 50624
rect 50440 50560 50456 50624
rect 50520 50560 50536 50624
rect 50600 50560 50608 50624
rect 50288 49536 50608 50560
rect 50288 49472 50296 49536
rect 50360 49472 50376 49536
rect 50440 49472 50456 49536
rect 50520 49472 50536 49536
rect 50600 49472 50608 49536
rect 50288 48448 50608 49472
rect 50288 48384 50296 48448
rect 50360 48384 50376 48448
rect 50440 48384 50456 48448
rect 50520 48384 50536 48448
rect 50600 48384 50608 48448
rect 50288 47360 50608 48384
rect 50288 47296 50296 47360
rect 50360 47296 50376 47360
rect 50440 47296 50456 47360
rect 50520 47296 50536 47360
rect 50600 47296 50608 47360
rect 50288 46272 50608 47296
rect 50288 46208 50296 46272
rect 50360 46208 50376 46272
rect 50440 46208 50456 46272
rect 50520 46208 50536 46272
rect 50600 46208 50608 46272
rect 50288 45184 50608 46208
rect 50288 45120 50296 45184
rect 50360 45120 50376 45184
rect 50440 45120 50456 45184
rect 50520 45120 50536 45184
rect 50600 45120 50608 45184
rect 50288 44096 50608 45120
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 43008 50608 44032
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 41920 50608 42944
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 40832 50608 41856
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 39744 50608 40768
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 38656 50608 39680
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 37568 50608 38592
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 36480 50608 37504
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 35392 50608 36416
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 34304 50608 35328
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 33216 50608 34240
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 32128 50608 33152
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 31040 50608 32064
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 29952 50608 30976
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 28864 50608 29888
rect 50288 28800 50296 28864
rect 50360 28800 50376 28864
rect 50440 28800 50456 28864
rect 50520 28800 50536 28864
rect 50600 28800 50608 28864
rect 50288 27776 50608 28800
rect 50288 27712 50296 27776
rect 50360 27712 50376 27776
rect 50440 27712 50456 27776
rect 50520 27712 50536 27776
rect 50600 27712 50608 27776
rect 50288 26688 50608 27712
rect 50288 26624 50296 26688
rect 50360 26624 50376 26688
rect 50440 26624 50456 26688
rect 50520 26624 50536 26688
rect 50600 26624 50608 26688
rect 50288 25600 50608 26624
rect 50288 25536 50296 25600
rect 50360 25536 50376 25600
rect 50440 25536 50456 25600
rect 50520 25536 50536 25600
rect 50600 25536 50608 25600
rect 50288 24512 50608 25536
rect 50288 24448 50296 24512
rect 50360 24448 50376 24512
rect 50440 24448 50456 24512
rect 50520 24448 50536 24512
rect 50600 24448 50608 24512
rect 50288 23424 50608 24448
rect 50288 23360 50296 23424
rect 50360 23360 50376 23424
rect 50440 23360 50456 23424
rect 50520 23360 50536 23424
rect 50600 23360 50608 23424
rect 50288 22336 50608 23360
rect 50288 22272 50296 22336
rect 50360 22272 50376 22336
rect 50440 22272 50456 22336
rect 50520 22272 50536 22336
rect 50600 22272 50608 22336
rect 50288 21248 50608 22272
rect 50288 21184 50296 21248
rect 50360 21184 50376 21248
rect 50440 21184 50456 21248
rect 50520 21184 50536 21248
rect 50600 21184 50608 21248
rect 50288 20160 50608 21184
rect 50288 20096 50296 20160
rect 50360 20096 50376 20160
rect 50440 20096 50456 20160
rect 50520 20096 50536 20160
rect 50600 20096 50608 20160
rect 50288 19072 50608 20096
rect 50288 19008 50296 19072
rect 50360 19008 50376 19072
rect 50440 19008 50456 19072
rect 50520 19008 50536 19072
rect 50600 19008 50608 19072
rect 50288 17984 50608 19008
rect 50288 17920 50296 17984
rect 50360 17920 50376 17984
rect 50440 17920 50456 17984
rect 50520 17920 50536 17984
rect 50600 17920 50608 17984
rect 50288 16896 50608 17920
rect 50288 16832 50296 16896
rect 50360 16832 50376 16896
rect 50440 16832 50456 16896
rect 50520 16832 50536 16896
rect 50600 16832 50608 16896
rect 50288 15808 50608 16832
rect 50288 15744 50296 15808
rect 50360 15744 50376 15808
rect 50440 15744 50456 15808
rect 50520 15744 50536 15808
rect 50600 15744 50608 15808
rect 50288 14720 50608 15744
rect 50288 14656 50296 14720
rect 50360 14656 50376 14720
rect 50440 14656 50456 14720
rect 50520 14656 50536 14720
rect 50600 14656 50608 14720
rect 50288 13632 50608 14656
rect 50288 13568 50296 13632
rect 50360 13568 50376 13632
rect 50440 13568 50456 13632
rect 50520 13568 50536 13632
rect 50600 13568 50608 13632
rect 50288 12544 50608 13568
rect 50288 12480 50296 12544
rect 50360 12480 50376 12544
rect 50440 12480 50456 12544
rect 50520 12480 50536 12544
rect 50600 12480 50608 12544
rect 50288 11456 50608 12480
rect 50288 11392 50296 11456
rect 50360 11392 50376 11456
rect 50440 11392 50456 11456
rect 50520 11392 50536 11456
rect 50600 11392 50608 11456
rect 50288 10368 50608 11392
rect 50288 10304 50296 10368
rect 50360 10304 50376 10368
rect 50440 10304 50456 10368
rect 50520 10304 50536 10368
rect 50600 10304 50608 10368
rect 50288 9280 50608 10304
rect 50288 9216 50296 9280
rect 50360 9216 50376 9280
rect 50440 9216 50456 9280
rect 50520 9216 50536 9280
rect 50600 9216 50608 9280
rect 50288 8192 50608 9216
rect 50288 8128 50296 8192
rect 50360 8128 50376 8192
rect 50440 8128 50456 8192
rect 50520 8128 50536 8192
rect 50600 8128 50608 8192
rect 50288 7104 50608 8128
rect 50288 7040 50296 7104
rect 50360 7040 50376 7104
rect 50440 7040 50456 7104
rect 50520 7040 50536 7104
rect 50600 7040 50608 7104
rect 50288 6016 50608 7040
rect 50288 5952 50296 6016
rect 50360 5952 50376 6016
rect 50440 5952 50456 6016
rect 50520 5952 50536 6016
rect 50600 5952 50608 6016
rect 50288 4928 50608 5952
rect 50288 4864 50296 4928
rect 50360 4864 50376 4928
rect 50440 4864 50456 4928
rect 50520 4864 50536 4928
rect 50600 4864 50608 4928
rect 50288 3840 50608 4864
rect 50288 3776 50296 3840
rect 50360 3776 50376 3840
rect 50440 3776 50456 3840
rect 50520 3776 50536 3840
rect 50600 3776 50608 3840
rect 50288 2752 50608 3776
rect 50288 2688 50296 2752
rect 50360 2688 50376 2752
rect 50440 2688 50456 2752
rect 50520 2688 50536 2752
rect 50600 2688 50608 2752
rect 34928 2128 35248 2144
rect 50288 2128 50608 2688
rect 50948 2176 51268 97376
rect 51608 2176 51928 97376
rect 52268 2176 52588 97376
rect 65648 96864 65968 97424
rect 81008 97408 81328 97424
rect 65648 96800 65656 96864
rect 65720 96800 65736 96864
rect 65800 96800 65816 96864
rect 65880 96800 65896 96864
rect 65960 96800 65968 96864
rect 65648 95776 65968 96800
rect 65648 95712 65656 95776
rect 65720 95712 65736 95776
rect 65800 95712 65816 95776
rect 65880 95712 65896 95776
rect 65960 95712 65968 95776
rect 65648 94688 65968 95712
rect 65648 94624 65656 94688
rect 65720 94624 65736 94688
rect 65800 94624 65816 94688
rect 65880 94624 65896 94688
rect 65960 94624 65968 94688
rect 65648 93600 65968 94624
rect 65648 93536 65656 93600
rect 65720 93536 65736 93600
rect 65800 93536 65816 93600
rect 65880 93536 65896 93600
rect 65960 93536 65968 93600
rect 65648 92512 65968 93536
rect 65648 92448 65656 92512
rect 65720 92448 65736 92512
rect 65800 92448 65816 92512
rect 65880 92448 65896 92512
rect 65960 92448 65968 92512
rect 65648 91424 65968 92448
rect 65648 91360 65656 91424
rect 65720 91360 65736 91424
rect 65800 91360 65816 91424
rect 65880 91360 65896 91424
rect 65960 91360 65968 91424
rect 65648 90336 65968 91360
rect 65648 90272 65656 90336
rect 65720 90272 65736 90336
rect 65800 90272 65816 90336
rect 65880 90272 65896 90336
rect 65960 90272 65968 90336
rect 65648 89248 65968 90272
rect 65648 89184 65656 89248
rect 65720 89184 65736 89248
rect 65800 89184 65816 89248
rect 65880 89184 65896 89248
rect 65960 89184 65968 89248
rect 65648 88160 65968 89184
rect 65648 88096 65656 88160
rect 65720 88096 65736 88160
rect 65800 88096 65816 88160
rect 65880 88096 65896 88160
rect 65960 88096 65968 88160
rect 65648 87072 65968 88096
rect 65648 87008 65656 87072
rect 65720 87008 65736 87072
rect 65800 87008 65816 87072
rect 65880 87008 65896 87072
rect 65960 87008 65968 87072
rect 65648 85984 65968 87008
rect 65648 85920 65656 85984
rect 65720 85920 65736 85984
rect 65800 85920 65816 85984
rect 65880 85920 65896 85984
rect 65960 85920 65968 85984
rect 65648 84896 65968 85920
rect 65648 84832 65656 84896
rect 65720 84832 65736 84896
rect 65800 84832 65816 84896
rect 65880 84832 65896 84896
rect 65960 84832 65968 84896
rect 65648 83808 65968 84832
rect 65648 83744 65656 83808
rect 65720 83744 65736 83808
rect 65800 83744 65816 83808
rect 65880 83744 65896 83808
rect 65960 83744 65968 83808
rect 65648 82720 65968 83744
rect 65648 82656 65656 82720
rect 65720 82656 65736 82720
rect 65800 82656 65816 82720
rect 65880 82656 65896 82720
rect 65960 82656 65968 82720
rect 65648 81632 65968 82656
rect 65648 81568 65656 81632
rect 65720 81568 65736 81632
rect 65800 81568 65816 81632
rect 65880 81568 65896 81632
rect 65960 81568 65968 81632
rect 65648 80544 65968 81568
rect 65648 80480 65656 80544
rect 65720 80480 65736 80544
rect 65800 80480 65816 80544
rect 65880 80480 65896 80544
rect 65960 80480 65968 80544
rect 65648 79456 65968 80480
rect 65648 79392 65656 79456
rect 65720 79392 65736 79456
rect 65800 79392 65816 79456
rect 65880 79392 65896 79456
rect 65960 79392 65968 79456
rect 65648 78368 65968 79392
rect 65648 78304 65656 78368
rect 65720 78304 65736 78368
rect 65800 78304 65816 78368
rect 65880 78304 65896 78368
rect 65960 78304 65968 78368
rect 65648 77280 65968 78304
rect 65648 77216 65656 77280
rect 65720 77216 65736 77280
rect 65800 77216 65816 77280
rect 65880 77216 65896 77280
rect 65960 77216 65968 77280
rect 65648 76192 65968 77216
rect 65648 76128 65656 76192
rect 65720 76128 65736 76192
rect 65800 76128 65816 76192
rect 65880 76128 65896 76192
rect 65960 76128 65968 76192
rect 65648 75104 65968 76128
rect 65648 75040 65656 75104
rect 65720 75040 65736 75104
rect 65800 75040 65816 75104
rect 65880 75040 65896 75104
rect 65960 75040 65968 75104
rect 65648 74016 65968 75040
rect 65648 73952 65656 74016
rect 65720 73952 65736 74016
rect 65800 73952 65816 74016
rect 65880 73952 65896 74016
rect 65960 73952 65968 74016
rect 65648 72928 65968 73952
rect 65648 72864 65656 72928
rect 65720 72864 65736 72928
rect 65800 72864 65816 72928
rect 65880 72864 65896 72928
rect 65960 72864 65968 72928
rect 65648 71840 65968 72864
rect 65648 71776 65656 71840
rect 65720 71776 65736 71840
rect 65800 71776 65816 71840
rect 65880 71776 65896 71840
rect 65960 71776 65968 71840
rect 65648 70752 65968 71776
rect 65648 70688 65656 70752
rect 65720 70688 65736 70752
rect 65800 70688 65816 70752
rect 65880 70688 65896 70752
rect 65960 70688 65968 70752
rect 65648 69664 65968 70688
rect 65648 69600 65656 69664
rect 65720 69600 65736 69664
rect 65800 69600 65816 69664
rect 65880 69600 65896 69664
rect 65960 69600 65968 69664
rect 65648 68576 65968 69600
rect 65648 68512 65656 68576
rect 65720 68512 65736 68576
rect 65800 68512 65816 68576
rect 65880 68512 65896 68576
rect 65960 68512 65968 68576
rect 65648 67488 65968 68512
rect 65648 67424 65656 67488
rect 65720 67424 65736 67488
rect 65800 67424 65816 67488
rect 65880 67424 65896 67488
rect 65960 67424 65968 67488
rect 65648 66400 65968 67424
rect 65648 66336 65656 66400
rect 65720 66336 65736 66400
rect 65800 66336 65816 66400
rect 65880 66336 65896 66400
rect 65960 66336 65968 66400
rect 65648 65312 65968 66336
rect 65648 65248 65656 65312
rect 65720 65248 65736 65312
rect 65800 65248 65816 65312
rect 65880 65248 65896 65312
rect 65960 65248 65968 65312
rect 65648 64224 65968 65248
rect 65648 64160 65656 64224
rect 65720 64160 65736 64224
rect 65800 64160 65816 64224
rect 65880 64160 65896 64224
rect 65960 64160 65968 64224
rect 65648 63136 65968 64160
rect 65648 63072 65656 63136
rect 65720 63072 65736 63136
rect 65800 63072 65816 63136
rect 65880 63072 65896 63136
rect 65960 63072 65968 63136
rect 65648 62048 65968 63072
rect 65648 61984 65656 62048
rect 65720 61984 65736 62048
rect 65800 61984 65816 62048
rect 65880 61984 65896 62048
rect 65960 61984 65968 62048
rect 65648 60960 65968 61984
rect 65648 60896 65656 60960
rect 65720 60896 65736 60960
rect 65800 60896 65816 60960
rect 65880 60896 65896 60960
rect 65960 60896 65968 60960
rect 65648 59872 65968 60896
rect 65648 59808 65656 59872
rect 65720 59808 65736 59872
rect 65800 59808 65816 59872
rect 65880 59808 65896 59872
rect 65960 59808 65968 59872
rect 65648 58784 65968 59808
rect 65648 58720 65656 58784
rect 65720 58720 65736 58784
rect 65800 58720 65816 58784
rect 65880 58720 65896 58784
rect 65960 58720 65968 58784
rect 65648 57696 65968 58720
rect 65648 57632 65656 57696
rect 65720 57632 65736 57696
rect 65800 57632 65816 57696
rect 65880 57632 65896 57696
rect 65960 57632 65968 57696
rect 65648 56608 65968 57632
rect 65648 56544 65656 56608
rect 65720 56544 65736 56608
rect 65800 56544 65816 56608
rect 65880 56544 65896 56608
rect 65960 56544 65968 56608
rect 65648 55520 65968 56544
rect 65648 55456 65656 55520
rect 65720 55456 65736 55520
rect 65800 55456 65816 55520
rect 65880 55456 65896 55520
rect 65960 55456 65968 55520
rect 65648 54432 65968 55456
rect 65648 54368 65656 54432
rect 65720 54368 65736 54432
rect 65800 54368 65816 54432
rect 65880 54368 65896 54432
rect 65960 54368 65968 54432
rect 65648 53344 65968 54368
rect 65648 53280 65656 53344
rect 65720 53280 65736 53344
rect 65800 53280 65816 53344
rect 65880 53280 65896 53344
rect 65960 53280 65968 53344
rect 65648 52256 65968 53280
rect 65648 52192 65656 52256
rect 65720 52192 65736 52256
rect 65800 52192 65816 52256
rect 65880 52192 65896 52256
rect 65960 52192 65968 52256
rect 65648 51168 65968 52192
rect 65648 51104 65656 51168
rect 65720 51104 65736 51168
rect 65800 51104 65816 51168
rect 65880 51104 65896 51168
rect 65960 51104 65968 51168
rect 65648 50080 65968 51104
rect 65648 50016 65656 50080
rect 65720 50016 65736 50080
rect 65800 50016 65816 50080
rect 65880 50016 65896 50080
rect 65960 50016 65968 50080
rect 65648 48992 65968 50016
rect 65648 48928 65656 48992
rect 65720 48928 65736 48992
rect 65800 48928 65816 48992
rect 65880 48928 65896 48992
rect 65960 48928 65968 48992
rect 65648 47904 65968 48928
rect 65648 47840 65656 47904
rect 65720 47840 65736 47904
rect 65800 47840 65816 47904
rect 65880 47840 65896 47904
rect 65960 47840 65968 47904
rect 65648 46816 65968 47840
rect 65648 46752 65656 46816
rect 65720 46752 65736 46816
rect 65800 46752 65816 46816
rect 65880 46752 65896 46816
rect 65960 46752 65968 46816
rect 65648 45728 65968 46752
rect 65648 45664 65656 45728
rect 65720 45664 65736 45728
rect 65800 45664 65816 45728
rect 65880 45664 65896 45728
rect 65960 45664 65968 45728
rect 65648 44640 65968 45664
rect 65648 44576 65656 44640
rect 65720 44576 65736 44640
rect 65800 44576 65816 44640
rect 65880 44576 65896 44640
rect 65960 44576 65968 44640
rect 65648 43552 65968 44576
rect 65648 43488 65656 43552
rect 65720 43488 65736 43552
rect 65800 43488 65816 43552
rect 65880 43488 65896 43552
rect 65960 43488 65968 43552
rect 65648 42464 65968 43488
rect 65648 42400 65656 42464
rect 65720 42400 65736 42464
rect 65800 42400 65816 42464
rect 65880 42400 65896 42464
rect 65960 42400 65968 42464
rect 65648 41376 65968 42400
rect 65648 41312 65656 41376
rect 65720 41312 65736 41376
rect 65800 41312 65816 41376
rect 65880 41312 65896 41376
rect 65960 41312 65968 41376
rect 65648 40288 65968 41312
rect 65648 40224 65656 40288
rect 65720 40224 65736 40288
rect 65800 40224 65816 40288
rect 65880 40224 65896 40288
rect 65960 40224 65968 40288
rect 65648 39200 65968 40224
rect 65648 39136 65656 39200
rect 65720 39136 65736 39200
rect 65800 39136 65816 39200
rect 65880 39136 65896 39200
rect 65960 39136 65968 39200
rect 65648 38112 65968 39136
rect 65648 38048 65656 38112
rect 65720 38048 65736 38112
rect 65800 38048 65816 38112
rect 65880 38048 65896 38112
rect 65960 38048 65968 38112
rect 65648 37024 65968 38048
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 35936 65968 36960
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 34848 65968 35872
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 33760 65968 34784
rect 65648 33696 65656 33760
rect 65720 33696 65736 33760
rect 65800 33696 65816 33760
rect 65880 33696 65896 33760
rect 65960 33696 65968 33760
rect 65648 32672 65968 33696
rect 65648 32608 65656 32672
rect 65720 32608 65736 32672
rect 65800 32608 65816 32672
rect 65880 32608 65896 32672
rect 65960 32608 65968 32672
rect 65648 31584 65968 32608
rect 65648 31520 65656 31584
rect 65720 31520 65736 31584
rect 65800 31520 65816 31584
rect 65880 31520 65896 31584
rect 65960 31520 65968 31584
rect 65648 30496 65968 31520
rect 65648 30432 65656 30496
rect 65720 30432 65736 30496
rect 65800 30432 65816 30496
rect 65880 30432 65896 30496
rect 65960 30432 65968 30496
rect 65648 29408 65968 30432
rect 65648 29344 65656 29408
rect 65720 29344 65736 29408
rect 65800 29344 65816 29408
rect 65880 29344 65896 29408
rect 65960 29344 65968 29408
rect 65648 28320 65968 29344
rect 65648 28256 65656 28320
rect 65720 28256 65736 28320
rect 65800 28256 65816 28320
rect 65880 28256 65896 28320
rect 65960 28256 65968 28320
rect 65648 27232 65968 28256
rect 65648 27168 65656 27232
rect 65720 27168 65736 27232
rect 65800 27168 65816 27232
rect 65880 27168 65896 27232
rect 65960 27168 65968 27232
rect 65648 26144 65968 27168
rect 65648 26080 65656 26144
rect 65720 26080 65736 26144
rect 65800 26080 65816 26144
rect 65880 26080 65896 26144
rect 65960 26080 65968 26144
rect 65648 25056 65968 26080
rect 65648 24992 65656 25056
rect 65720 24992 65736 25056
rect 65800 24992 65816 25056
rect 65880 24992 65896 25056
rect 65960 24992 65968 25056
rect 65648 23968 65968 24992
rect 65648 23904 65656 23968
rect 65720 23904 65736 23968
rect 65800 23904 65816 23968
rect 65880 23904 65896 23968
rect 65960 23904 65968 23968
rect 65648 22880 65968 23904
rect 65648 22816 65656 22880
rect 65720 22816 65736 22880
rect 65800 22816 65816 22880
rect 65880 22816 65896 22880
rect 65960 22816 65968 22880
rect 65648 21792 65968 22816
rect 65648 21728 65656 21792
rect 65720 21728 65736 21792
rect 65800 21728 65816 21792
rect 65880 21728 65896 21792
rect 65960 21728 65968 21792
rect 65648 20704 65968 21728
rect 65648 20640 65656 20704
rect 65720 20640 65736 20704
rect 65800 20640 65816 20704
rect 65880 20640 65896 20704
rect 65960 20640 65968 20704
rect 65648 19616 65968 20640
rect 65648 19552 65656 19616
rect 65720 19552 65736 19616
rect 65800 19552 65816 19616
rect 65880 19552 65896 19616
rect 65960 19552 65968 19616
rect 65648 18528 65968 19552
rect 65648 18464 65656 18528
rect 65720 18464 65736 18528
rect 65800 18464 65816 18528
rect 65880 18464 65896 18528
rect 65960 18464 65968 18528
rect 65648 17440 65968 18464
rect 65648 17376 65656 17440
rect 65720 17376 65736 17440
rect 65800 17376 65816 17440
rect 65880 17376 65896 17440
rect 65960 17376 65968 17440
rect 65648 16352 65968 17376
rect 65648 16288 65656 16352
rect 65720 16288 65736 16352
rect 65800 16288 65816 16352
rect 65880 16288 65896 16352
rect 65960 16288 65968 16352
rect 65648 15264 65968 16288
rect 65648 15200 65656 15264
rect 65720 15200 65736 15264
rect 65800 15200 65816 15264
rect 65880 15200 65896 15264
rect 65960 15200 65968 15264
rect 65648 14176 65968 15200
rect 65648 14112 65656 14176
rect 65720 14112 65736 14176
rect 65800 14112 65816 14176
rect 65880 14112 65896 14176
rect 65960 14112 65968 14176
rect 65648 13088 65968 14112
rect 65648 13024 65656 13088
rect 65720 13024 65736 13088
rect 65800 13024 65816 13088
rect 65880 13024 65896 13088
rect 65960 13024 65968 13088
rect 65648 12000 65968 13024
rect 65648 11936 65656 12000
rect 65720 11936 65736 12000
rect 65800 11936 65816 12000
rect 65880 11936 65896 12000
rect 65960 11936 65968 12000
rect 65648 10912 65968 11936
rect 65648 10848 65656 10912
rect 65720 10848 65736 10912
rect 65800 10848 65816 10912
rect 65880 10848 65896 10912
rect 65960 10848 65968 10912
rect 65648 9824 65968 10848
rect 65648 9760 65656 9824
rect 65720 9760 65736 9824
rect 65800 9760 65816 9824
rect 65880 9760 65896 9824
rect 65960 9760 65968 9824
rect 65648 8736 65968 9760
rect 65648 8672 65656 8736
rect 65720 8672 65736 8736
rect 65800 8672 65816 8736
rect 65880 8672 65896 8736
rect 65960 8672 65968 8736
rect 65648 7648 65968 8672
rect 65648 7584 65656 7648
rect 65720 7584 65736 7648
rect 65800 7584 65816 7648
rect 65880 7584 65896 7648
rect 65960 7584 65968 7648
rect 65648 6560 65968 7584
rect 65648 6496 65656 6560
rect 65720 6496 65736 6560
rect 65800 6496 65816 6560
rect 65880 6496 65896 6560
rect 65960 6496 65968 6560
rect 65648 5472 65968 6496
rect 65648 5408 65656 5472
rect 65720 5408 65736 5472
rect 65800 5408 65816 5472
rect 65880 5408 65896 5472
rect 65960 5408 65968 5472
rect 65648 4384 65968 5408
rect 65648 4320 65656 4384
rect 65720 4320 65736 4384
rect 65800 4320 65816 4384
rect 65880 4320 65896 4384
rect 65960 4320 65968 4384
rect 65648 3296 65968 4320
rect 65648 3232 65656 3296
rect 65720 3232 65736 3296
rect 65800 3232 65816 3296
rect 65880 3232 65896 3296
rect 65960 3232 65968 3296
rect 65648 2208 65968 3232
rect 65648 2144 65656 2208
rect 65720 2144 65736 2208
rect 65800 2144 65816 2208
rect 65880 2144 65896 2208
rect 65960 2144 65968 2208
rect 66308 2176 66628 97376
rect 66968 2176 67288 97376
rect 67628 2176 67948 97376
rect 81008 97344 81016 97408
rect 81080 97344 81096 97408
rect 81160 97344 81176 97408
rect 81240 97344 81256 97408
rect 81320 97344 81328 97408
rect 81008 96320 81328 97344
rect 81008 96256 81016 96320
rect 81080 96256 81096 96320
rect 81160 96256 81176 96320
rect 81240 96256 81256 96320
rect 81320 96256 81328 96320
rect 81008 95232 81328 96256
rect 81008 95168 81016 95232
rect 81080 95168 81096 95232
rect 81160 95168 81176 95232
rect 81240 95168 81256 95232
rect 81320 95168 81328 95232
rect 81008 94144 81328 95168
rect 81008 94080 81016 94144
rect 81080 94080 81096 94144
rect 81160 94080 81176 94144
rect 81240 94080 81256 94144
rect 81320 94080 81328 94144
rect 81008 93056 81328 94080
rect 81008 92992 81016 93056
rect 81080 92992 81096 93056
rect 81160 92992 81176 93056
rect 81240 92992 81256 93056
rect 81320 92992 81328 93056
rect 81008 91968 81328 92992
rect 81008 91904 81016 91968
rect 81080 91904 81096 91968
rect 81160 91904 81176 91968
rect 81240 91904 81256 91968
rect 81320 91904 81328 91968
rect 81008 90880 81328 91904
rect 81008 90816 81016 90880
rect 81080 90816 81096 90880
rect 81160 90816 81176 90880
rect 81240 90816 81256 90880
rect 81320 90816 81328 90880
rect 81008 89792 81328 90816
rect 81008 89728 81016 89792
rect 81080 89728 81096 89792
rect 81160 89728 81176 89792
rect 81240 89728 81256 89792
rect 81320 89728 81328 89792
rect 81008 88704 81328 89728
rect 81008 88640 81016 88704
rect 81080 88640 81096 88704
rect 81160 88640 81176 88704
rect 81240 88640 81256 88704
rect 81320 88640 81328 88704
rect 81008 87616 81328 88640
rect 81008 87552 81016 87616
rect 81080 87552 81096 87616
rect 81160 87552 81176 87616
rect 81240 87552 81256 87616
rect 81320 87552 81328 87616
rect 81008 86528 81328 87552
rect 81008 86464 81016 86528
rect 81080 86464 81096 86528
rect 81160 86464 81176 86528
rect 81240 86464 81256 86528
rect 81320 86464 81328 86528
rect 81008 85440 81328 86464
rect 81008 85376 81016 85440
rect 81080 85376 81096 85440
rect 81160 85376 81176 85440
rect 81240 85376 81256 85440
rect 81320 85376 81328 85440
rect 81008 84352 81328 85376
rect 81008 84288 81016 84352
rect 81080 84288 81096 84352
rect 81160 84288 81176 84352
rect 81240 84288 81256 84352
rect 81320 84288 81328 84352
rect 81008 83264 81328 84288
rect 81008 83200 81016 83264
rect 81080 83200 81096 83264
rect 81160 83200 81176 83264
rect 81240 83200 81256 83264
rect 81320 83200 81328 83264
rect 81008 82176 81328 83200
rect 81008 82112 81016 82176
rect 81080 82112 81096 82176
rect 81160 82112 81176 82176
rect 81240 82112 81256 82176
rect 81320 82112 81328 82176
rect 81008 81088 81328 82112
rect 81008 81024 81016 81088
rect 81080 81024 81096 81088
rect 81160 81024 81176 81088
rect 81240 81024 81256 81088
rect 81320 81024 81328 81088
rect 81008 80000 81328 81024
rect 81008 79936 81016 80000
rect 81080 79936 81096 80000
rect 81160 79936 81176 80000
rect 81240 79936 81256 80000
rect 81320 79936 81328 80000
rect 81008 78912 81328 79936
rect 81008 78848 81016 78912
rect 81080 78848 81096 78912
rect 81160 78848 81176 78912
rect 81240 78848 81256 78912
rect 81320 78848 81328 78912
rect 81008 77824 81328 78848
rect 81008 77760 81016 77824
rect 81080 77760 81096 77824
rect 81160 77760 81176 77824
rect 81240 77760 81256 77824
rect 81320 77760 81328 77824
rect 81008 76736 81328 77760
rect 81008 76672 81016 76736
rect 81080 76672 81096 76736
rect 81160 76672 81176 76736
rect 81240 76672 81256 76736
rect 81320 76672 81328 76736
rect 81008 75648 81328 76672
rect 81008 75584 81016 75648
rect 81080 75584 81096 75648
rect 81160 75584 81176 75648
rect 81240 75584 81256 75648
rect 81320 75584 81328 75648
rect 81008 74560 81328 75584
rect 81008 74496 81016 74560
rect 81080 74496 81096 74560
rect 81160 74496 81176 74560
rect 81240 74496 81256 74560
rect 81320 74496 81328 74560
rect 81008 73472 81328 74496
rect 81008 73408 81016 73472
rect 81080 73408 81096 73472
rect 81160 73408 81176 73472
rect 81240 73408 81256 73472
rect 81320 73408 81328 73472
rect 81008 72384 81328 73408
rect 81008 72320 81016 72384
rect 81080 72320 81096 72384
rect 81160 72320 81176 72384
rect 81240 72320 81256 72384
rect 81320 72320 81328 72384
rect 81008 71296 81328 72320
rect 81008 71232 81016 71296
rect 81080 71232 81096 71296
rect 81160 71232 81176 71296
rect 81240 71232 81256 71296
rect 81320 71232 81328 71296
rect 81008 70208 81328 71232
rect 81008 70144 81016 70208
rect 81080 70144 81096 70208
rect 81160 70144 81176 70208
rect 81240 70144 81256 70208
rect 81320 70144 81328 70208
rect 81008 69120 81328 70144
rect 81008 69056 81016 69120
rect 81080 69056 81096 69120
rect 81160 69056 81176 69120
rect 81240 69056 81256 69120
rect 81320 69056 81328 69120
rect 81008 68032 81328 69056
rect 81008 67968 81016 68032
rect 81080 67968 81096 68032
rect 81160 67968 81176 68032
rect 81240 67968 81256 68032
rect 81320 67968 81328 68032
rect 81008 66944 81328 67968
rect 81008 66880 81016 66944
rect 81080 66880 81096 66944
rect 81160 66880 81176 66944
rect 81240 66880 81256 66944
rect 81320 66880 81328 66944
rect 81008 65856 81328 66880
rect 81008 65792 81016 65856
rect 81080 65792 81096 65856
rect 81160 65792 81176 65856
rect 81240 65792 81256 65856
rect 81320 65792 81328 65856
rect 81008 64768 81328 65792
rect 81008 64704 81016 64768
rect 81080 64704 81096 64768
rect 81160 64704 81176 64768
rect 81240 64704 81256 64768
rect 81320 64704 81328 64768
rect 81008 63680 81328 64704
rect 81008 63616 81016 63680
rect 81080 63616 81096 63680
rect 81160 63616 81176 63680
rect 81240 63616 81256 63680
rect 81320 63616 81328 63680
rect 81008 62592 81328 63616
rect 81008 62528 81016 62592
rect 81080 62528 81096 62592
rect 81160 62528 81176 62592
rect 81240 62528 81256 62592
rect 81320 62528 81328 62592
rect 81008 61504 81328 62528
rect 81008 61440 81016 61504
rect 81080 61440 81096 61504
rect 81160 61440 81176 61504
rect 81240 61440 81256 61504
rect 81320 61440 81328 61504
rect 81008 60416 81328 61440
rect 81008 60352 81016 60416
rect 81080 60352 81096 60416
rect 81160 60352 81176 60416
rect 81240 60352 81256 60416
rect 81320 60352 81328 60416
rect 81008 59328 81328 60352
rect 81008 59264 81016 59328
rect 81080 59264 81096 59328
rect 81160 59264 81176 59328
rect 81240 59264 81256 59328
rect 81320 59264 81328 59328
rect 81008 58240 81328 59264
rect 81008 58176 81016 58240
rect 81080 58176 81096 58240
rect 81160 58176 81176 58240
rect 81240 58176 81256 58240
rect 81320 58176 81328 58240
rect 81008 57152 81328 58176
rect 81008 57088 81016 57152
rect 81080 57088 81096 57152
rect 81160 57088 81176 57152
rect 81240 57088 81256 57152
rect 81320 57088 81328 57152
rect 81008 56064 81328 57088
rect 81008 56000 81016 56064
rect 81080 56000 81096 56064
rect 81160 56000 81176 56064
rect 81240 56000 81256 56064
rect 81320 56000 81328 56064
rect 81008 54976 81328 56000
rect 81008 54912 81016 54976
rect 81080 54912 81096 54976
rect 81160 54912 81176 54976
rect 81240 54912 81256 54976
rect 81320 54912 81328 54976
rect 81008 53888 81328 54912
rect 81008 53824 81016 53888
rect 81080 53824 81096 53888
rect 81160 53824 81176 53888
rect 81240 53824 81256 53888
rect 81320 53824 81328 53888
rect 81008 52800 81328 53824
rect 81008 52736 81016 52800
rect 81080 52736 81096 52800
rect 81160 52736 81176 52800
rect 81240 52736 81256 52800
rect 81320 52736 81328 52800
rect 81008 51712 81328 52736
rect 81008 51648 81016 51712
rect 81080 51648 81096 51712
rect 81160 51648 81176 51712
rect 81240 51648 81256 51712
rect 81320 51648 81328 51712
rect 81008 50624 81328 51648
rect 81008 50560 81016 50624
rect 81080 50560 81096 50624
rect 81160 50560 81176 50624
rect 81240 50560 81256 50624
rect 81320 50560 81328 50624
rect 81008 49536 81328 50560
rect 81008 49472 81016 49536
rect 81080 49472 81096 49536
rect 81160 49472 81176 49536
rect 81240 49472 81256 49536
rect 81320 49472 81328 49536
rect 81008 48448 81328 49472
rect 81008 48384 81016 48448
rect 81080 48384 81096 48448
rect 81160 48384 81176 48448
rect 81240 48384 81256 48448
rect 81320 48384 81328 48448
rect 81008 47360 81328 48384
rect 81008 47296 81016 47360
rect 81080 47296 81096 47360
rect 81160 47296 81176 47360
rect 81240 47296 81256 47360
rect 81320 47296 81328 47360
rect 81008 46272 81328 47296
rect 81008 46208 81016 46272
rect 81080 46208 81096 46272
rect 81160 46208 81176 46272
rect 81240 46208 81256 46272
rect 81320 46208 81328 46272
rect 81008 45184 81328 46208
rect 81008 45120 81016 45184
rect 81080 45120 81096 45184
rect 81160 45120 81176 45184
rect 81240 45120 81256 45184
rect 81320 45120 81328 45184
rect 81008 44096 81328 45120
rect 81008 44032 81016 44096
rect 81080 44032 81096 44096
rect 81160 44032 81176 44096
rect 81240 44032 81256 44096
rect 81320 44032 81328 44096
rect 81008 43008 81328 44032
rect 81008 42944 81016 43008
rect 81080 42944 81096 43008
rect 81160 42944 81176 43008
rect 81240 42944 81256 43008
rect 81320 42944 81328 43008
rect 81008 41920 81328 42944
rect 81008 41856 81016 41920
rect 81080 41856 81096 41920
rect 81160 41856 81176 41920
rect 81240 41856 81256 41920
rect 81320 41856 81328 41920
rect 81008 40832 81328 41856
rect 81008 40768 81016 40832
rect 81080 40768 81096 40832
rect 81160 40768 81176 40832
rect 81240 40768 81256 40832
rect 81320 40768 81328 40832
rect 81008 39744 81328 40768
rect 81008 39680 81016 39744
rect 81080 39680 81096 39744
rect 81160 39680 81176 39744
rect 81240 39680 81256 39744
rect 81320 39680 81328 39744
rect 81008 38656 81328 39680
rect 81008 38592 81016 38656
rect 81080 38592 81096 38656
rect 81160 38592 81176 38656
rect 81240 38592 81256 38656
rect 81320 38592 81328 38656
rect 81008 37568 81328 38592
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 36480 81328 37504
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 35392 81328 36416
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 34304 81328 35328
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 33216 81328 34240
rect 81008 33152 81016 33216
rect 81080 33152 81096 33216
rect 81160 33152 81176 33216
rect 81240 33152 81256 33216
rect 81320 33152 81328 33216
rect 81008 32128 81328 33152
rect 81008 32064 81016 32128
rect 81080 32064 81096 32128
rect 81160 32064 81176 32128
rect 81240 32064 81256 32128
rect 81320 32064 81328 32128
rect 81008 31040 81328 32064
rect 81008 30976 81016 31040
rect 81080 30976 81096 31040
rect 81160 30976 81176 31040
rect 81240 30976 81256 31040
rect 81320 30976 81328 31040
rect 81008 29952 81328 30976
rect 81008 29888 81016 29952
rect 81080 29888 81096 29952
rect 81160 29888 81176 29952
rect 81240 29888 81256 29952
rect 81320 29888 81328 29952
rect 81008 28864 81328 29888
rect 81008 28800 81016 28864
rect 81080 28800 81096 28864
rect 81160 28800 81176 28864
rect 81240 28800 81256 28864
rect 81320 28800 81328 28864
rect 81008 27776 81328 28800
rect 81008 27712 81016 27776
rect 81080 27712 81096 27776
rect 81160 27712 81176 27776
rect 81240 27712 81256 27776
rect 81320 27712 81328 27776
rect 81008 26688 81328 27712
rect 81008 26624 81016 26688
rect 81080 26624 81096 26688
rect 81160 26624 81176 26688
rect 81240 26624 81256 26688
rect 81320 26624 81328 26688
rect 81008 25600 81328 26624
rect 81008 25536 81016 25600
rect 81080 25536 81096 25600
rect 81160 25536 81176 25600
rect 81240 25536 81256 25600
rect 81320 25536 81328 25600
rect 81008 24512 81328 25536
rect 81008 24448 81016 24512
rect 81080 24448 81096 24512
rect 81160 24448 81176 24512
rect 81240 24448 81256 24512
rect 81320 24448 81328 24512
rect 81008 23424 81328 24448
rect 81008 23360 81016 23424
rect 81080 23360 81096 23424
rect 81160 23360 81176 23424
rect 81240 23360 81256 23424
rect 81320 23360 81328 23424
rect 81008 22336 81328 23360
rect 81008 22272 81016 22336
rect 81080 22272 81096 22336
rect 81160 22272 81176 22336
rect 81240 22272 81256 22336
rect 81320 22272 81328 22336
rect 81008 21248 81328 22272
rect 81008 21184 81016 21248
rect 81080 21184 81096 21248
rect 81160 21184 81176 21248
rect 81240 21184 81256 21248
rect 81320 21184 81328 21248
rect 81008 20160 81328 21184
rect 81008 20096 81016 20160
rect 81080 20096 81096 20160
rect 81160 20096 81176 20160
rect 81240 20096 81256 20160
rect 81320 20096 81328 20160
rect 81008 19072 81328 20096
rect 81008 19008 81016 19072
rect 81080 19008 81096 19072
rect 81160 19008 81176 19072
rect 81240 19008 81256 19072
rect 81320 19008 81328 19072
rect 81008 17984 81328 19008
rect 81008 17920 81016 17984
rect 81080 17920 81096 17984
rect 81160 17920 81176 17984
rect 81240 17920 81256 17984
rect 81320 17920 81328 17984
rect 81008 16896 81328 17920
rect 81008 16832 81016 16896
rect 81080 16832 81096 16896
rect 81160 16832 81176 16896
rect 81240 16832 81256 16896
rect 81320 16832 81328 16896
rect 81008 15808 81328 16832
rect 81008 15744 81016 15808
rect 81080 15744 81096 15808
rect 81160 15744 81176 15808
rect 81240 15744 81256 15808
rect 81320 15744 81328 15808
rect 81008 14720 81328 15744
rect 81008 14656 81016 14720
rect 81080 14656 81096 14720
rect 81160 14656 81176 14720
rect 81240 14656 81256 14720
rect 81320 14656 81328 14720
rect 81008 13632 81328 14656
rect 81008 13568 81016 13632
rect 81080 13568 81096 13632
rect 81160 13568 81176 13632
rect 81240 13568 81256 13632
rect 81320 13568 81328 13632
rect 81008 12544 81328 13568
rect 81008 12480 81016 12544
rect 81080 12480 81096 12544
rect 81160 12480 81176 12544
rect 81240 12480 81256 12544
rect 81320 12480 81328 12544
rect 81008 11456 81328 12480
rect 81008 11392 81016 11456
rect 81080 11392 81096 11456
rect 81160 11392 81176 11456
rect 81240 11392 81256 11456
rect 81320 11392 81328 11456
rect 81008 10368 81328 11392
rect 81008 10304 81016 10368
rect 81080 10304 81096 10368
rect 81160 10304 81176 10368
rect 81240 10304 81256 10368
rect 81320 10304 81328 10368
rect 81008 9280 81328 10304
rect 81008 9216 81016 9280
rect 81080 9216 81096 9280
rect 81160 9216 81176 9280
rect 81240 9216 81256 9280
rect 81320 9216 81328 9280
rect 81008 8192 81328 9216
rect 81008 8128 81016 8192
rect 81080 8128 81096 8192
rect 81160 8128 81176 8192
rect 81240 8128 81256 8192
rect 81320 8128 81328 8192
rect 81008 7104 81328 8128
rect 81008 7040 81016 7104
rect 81080 7040 81096 7104
rect 81160 7040 81176 7104
rect 81240 7040 81256 7104
rect 81320 7040 81328 7104
rect 81008 6016 81328 7040
rect 81008 5952 81016 6016
rect 81080 5952 81096 6016
rect 81160 5952 81176 6016
rect 81240 5952 81256 6016
rect 81320 5952 81328 6016
rect 81008 4928 81328 5952
rect 81008 4864 81016 4928
rect 81080 4864 81096 4928
rect 81160 4864 81176 4928
rect 81240 4864 81256 4928
rect 81320 4864 81328 4928
rect 81008 3840 81328 4864
rect 81008 3776 81016 3840
rect 81080 3776 81096 3840
rect 81160 3776 81176 3840
rect 81240 3776 81256 3840
rect 81320 3776 81328 3840
rect 81008 2752 81328 3776
rect 81008 2688 81016 2752
rect 81080 2688 81096 2752
rect 81160 2688 81176 2752
rect 81240 2688 81256 2752
rect 81320 2688 81328 2752
rect 65648 2128 65968 2144
rect 81008 2128 81328 2688
rect 81668 2176 81988 97376
rect 82328 2176 82648 97376
rect 82988 2176 83308 97376
rect 96368 96864 96688 97424
rect 96368 96800 96376 96864
rect 96440 96800 96456 96864
rect 96520 96800 96536 96864
rect 96600 96800 96616 96864
rect 96680 96800 96688 96864
rect 96368 95776 96688 96800
rect 96368 95712 96376 95776
rect 96440 95712 96456 95776
rect 96520 95712 96536 95776
rect 96600 95712 96616 95776
rect 96680 95712 96688 95776
rect 96368 94688 96688 95712
rect 96368 94624 96376 94688
rect 96440 94624 96456 94688
rect 96520 94624 96536 94688
rect 96600 94624 96616 94688
rect 96680 94624 96688 94688
rect 96368 93600 96688 94624
rect 96368 93536 96376 93600
rect 96440 93536 96456 93600
rect 96520 93536 96536 93600
rect 96600 93536 96616 93600
rect 96680 93536 96688 93600
rect 96368 92512 96688 93536
rect 96368 92448 96376 92512
rect 96440 92448 96456 92512
rect 96520 92448 96536 92512
rect 96600 92448 96616 92512
rect 96680 92448 96688 92512
rect 96368 91424 96688 92448
rect 96368 91360 96376 91424
rect 96440 91360 96456 91424
rect 96520 91360 96536 91424
rect 96600 91360 96616 91424
rect 96680 91360 96688 91424
rect 96368 90336 96688 91360
rect 96368 90272 96376 90336
rect 96440 90272 96456 90336
rect 96520 90272 96536 90336
rect 96600 90272 96616 90336
rect 96680 90272 96688 90336
rect 96368 89248 96688 90272
rect 96368 89184 96376 89248
rect 96440 89184 96456 89248
rect 96520 89184 96536 89248
rect 96600 89184 96616 89248
rect 96680 89184 96688 89248
rect 96368 88160 96688 89184
rect 96368 88096 96376 88160
rect 96440 88096 96456 88160
rect 96520 88096 96536 88160
rect 96600 88096 96616 88160
rect 96680 88096 96688 88160
rect 96368 87072 96688 88096
rect 96368 87008 96376 87072
rect 96440 87008 96456 87072
rect 96520 87008 96536 87072
rect 96600 87008 96616 87072
rect 96680 87008 96688 87072
rect 96368 85984 96688 87008
rect 96368 85920 96376 85984
rect 96440 85920 96456 85984
rect 96520 85920 96536 85984
rect 96600 85920 96616 85984
rect 96680 85920 96688 85984
rect 96368 84896 96688 85920
rect 96368 84832 96376 84896
rect 96440 84832 96456 84896
rect 96520 84832 96536 84896
rect 96600 84832 96616 84896
rect 96680 84832 96688 84896
rect 96368 83808 96688 84832
rect 96368 83744 96376 83808
rect 96440 83744 96456 83808
rect 96520 83744 96536 83808
rect 96600 83744 96616 83808
rect 96680 83744 96688 83808
rect 96368 82720 96688 83744
rect 96368 82656 96376 82720
rect 96440 82656 96456 82720
rect 96520 82656 96536 82720
rect 96600 82656 96616 82720
rect 96680 82656 96688 82720
rect 96368 81632 96688 82656
rect 96368 81568 96376 81632
rect 96440 81568 96456 81632
rect 96520 81568 96536 81632
rect 96600 81568 96616 81632
rect 96680 81568 96688 81632
rect 96368 80544 96688 81568
rect 96368 80480 96376 80544
rect 96440 80480 96456 80544
rect 96520 80480 96536 80544
rect 96600 80480 96616 80544
rect 96680 80480 96688 80544
rect 96368 79456 96688 80480
rect 96368 79392 96376 79456
rect 96440 79392 96456 79456
rect 96520 79392 96536 79456
rect 96600 79392 96616 79456
rect 96680 79392 96688 79456
rect 96368 78368 96688 79392
rect 96368 78304 96376 78368
rect 96440 78304 96456 78368
rect 96520 78304 96536 78368
rect 96600 78304 96616 78368
rect 96680 78304 96688 78368
rect 96368 77280 96688 78304
rect 96368 77216 96376 77280
rect 96440 77216 96456 77280
rect 96520 77216 96536 77280
rect 96600 77216 96616 77280
rect 96680 77216 96688 77280
rect 96368 76192 96688 77216
rect 96368 76128 96376 76192
rect 96440 76128 96456 76192
rect 96520 76128 96536 76192
rect 96600 76128 96616 76192
rect 96680 76128 96688 76192
rect 96368 75104 96688 76128
rect 96368 75040 96376 75104
rect 96440 75040 96456 75104
rect 96520 75040 96536 75104
rect 96600 75040 96616 75104
rect 96680 75040 96688 75104
rect 96368 74016 96688 75040
rect 96368 73952 96376 74016
rect 96440 73952 96456 74016
rect 96520 73952 96536 74016
rect 96600 73952 96616 74016
rect 96680 73952 96688 74016
rect 96368 72928 96688 73952
rect 96368 72864 96376 72928
rect 96440 72864 96456 72928
rect 96520 72864 96536 72928
rect 96600 72864 96616 72928
rect 96680 72864 96688 72928
rect 96368 71840 96688 72864
rect 96368 71776 96376 71840
rect 96440 71776 96456 71840
rect 96520 71776 96536 71840
rect 96600 71776 96616 71840
rect 96680 71776 96688 71840
rect 96368 70752 96688 71776
rect 96368 70688 96376 70752
rect 96440 70688 96456 70752
rect 96520 70688 96536 70752
rect 96600 70688 96616 70752
rect 96680 70688 96688 70752
rect 96368 69664 96688 70688
rect 96368 69600 96376 69664
rect 96440 69600 96456 69664
rect 96520 69600 96536 69664
rect 96600 69600 96616 69664
rect 96680 69600 96688 69664
rect 96368 68576 96688 69600
rect 96368 68512 96376 68576
rect 96440 68512 96456 68576
rect 96520 68512 96536 68576
rect 96600 68512 96616 68576
rect 96680 68512 96688 68576
rect 96368 67488 96688 68512
rect 96368 67424 96376 67488
rect 96440 67424 96456 67488
rect 96520 67424 96536 67488
rect 96600 67424 96616 67488
rect 96680 67424 96688 67488
rect 96368 66400 96688 67424
rect 96368 66336 96376 66400
rect 96440 66336 96456 66400
rect 96520 66336 96536 66400
rect 96600 66336 96616 66400
rect 96680 66336 96688 66400
rect 96368 65312 96688 66336
rect 96368 65248 96376 65312
rect 96440 65248 96456 65312
rect 96520 65248 96536 65312
rect 96600 65248 96616 65312
rect 96680 65248 96688 65312
rect 96368 64224 96688 65248
rect 96368 64160 96376 64224
rect 96440 64160 96456 64224
rect 96520 64160 96536 64224
rect 96600 64160 96616 64224
rect 96680 64160 96688 64224
rect 96368 63136 96688 64160
rect 96368 63072 96376 63136
rect 96440 63072 96456 63136
rect 96520 63072 96536 63136
rect 96600 63072 96616 63136
rect 96680 63072 96688 63136
rect 96368 62048 96688 63072
rect 96368 61984 96376 62048
rect 96440 61984 96456 62048
rect 96520 61984 96536 62048
rect 96600 61984 96616 62048
rect 96680 61984 96688 62048
rect 96368 60960 96688 61984
rect 96368 60896 96376 60960
rect 96440 60896 96456 60960
rect 96520 60896 96536 60960
rect 96600 60896 96616 60960
rect 96680 60896 96688 60960
rect 96368 59872 96688 60896
rect 96368 59808 96376 59872
rect 96440 59808 96456 59872
rect 96520 59808 96536 59872
rect 96600 59808 96616 59872
rect 96680 59808 96688 59872
rect 96368 58784 96688 59808
rect 96368 58720 96376 58784
rect 96440 58720 96456 58784
rect 96520 58720 96536 58784
rect 96600 58720 96616 58784
rect 96680 58720 96688 58784
rect 96368 57696 96688 58720
rect 96368 57632 96376 57696
rect 96440 57632 96456 57696
rect 96520 57632 96536 57696
rect 96600 57632 96616 57696
rect 96680 57632 96688 57696
rect 96368 56608 96688 57632
rect 96368 56544 96376 56608
rect 96440 56544 96456 56608
rect 96520 56544 96536 56608
rect 96600 56544 96616 56608
rect 96680 56544 96688 56608
rect 96368 55520 96688 56544
rect 96368 55456 96376 55520
rect 96440 55456 96456 55520
rect 96520 55456 96536 55520
rect 96600 55456 96616 55520
rect 96680 55456 96688 55520
rect 96368 54432 96688 55456
rect 96368 54368 96376 54432
rect 96440 54368 96456 54432
rect 96520 54368 96536 54432
rect 96600 54368 96616 54432
rect 96680 54368 96688 54432
rect 96368 53344 96688 54368
rect 96368 53280 96376 53344
rect 96440 53280 96456 53344
rect 96520 53280 96536 53344
rect 96600 53280 96616 53344
rect 96680 53280 96688 53344
rect 96368 52256 96688 53280
rect 96368 52192 96376 52256
rect 96440 52192 96456 52256
rect 96520 52192 96536 52256
rect 96600 52192 96616 52256
rect 96680 52192 96688 52256
rect 96368 51168 96688 52192
rect 96368 51104 96376 51168
rect 96440 51104 96456 51168
rect 96520 51104 96536 51168
rect 96600 51104 96616 51168
rect 96680 51104 96688 51168
rect 96368 50080 96688 51104
rect 96368 50016 96376 50080
rect 96440 50016 96456 50080
rect 96520 50016 96536 50080
rect 96600 50016 96616 50080
rect 96680 50016 96688 50080
rect 96368 48992 96688 50016
rect 96368 48928 96376 48992
rect 96440 48928 96456 48992
rect 96520 48928 96536 48992
rect 96600 48928 96616 48992
rect 96680 48928 96688 48992
rect 96368 47904 96688 48928
rect 96368 47840 96376 47904
rect 96440 47840 96456 47904
rect 96520 47840 96536 47904
rect 96600 47840 96616 47904
rect 96680 47840 96688 47904
rect 96368 46816 96688 47840
rect 96368 46752 96376 46816
rect 96440 46752 96456 46816
rect 96520 46752 96536 46816
rect 96600 46752 96616 46816
rect 96680 46752 96688 46816
rect 96368 45728 96688 46752
rect 96368 45664 96376 45728
rect 96440 45664 96456 45728
rect 96520 45664 96536 45728
rect 96600 45664 96616 45728
rect 96680 45664 96688 45728
rect 96368 44640 96688 45664
rect 96368 44576 96376 44640
rect 96440 44576 96456 44640
rect 96520 44576 96536 44640
rect 96600 44576 96616 44640
rect 96680 44576 96688 44640
rect 96368 43552 96688 44576
rect 96368 43488 96376 43552
rect 96440 43488 96456 43552
rect 96520 43488 96536 43552
rect 96600 43488 96616 43552
rect 96680 43488 96688 43552
rect 96368 42464 96688 43488
rect 96368 42400 96376 42464
rect 96440 42400 96456 42464
rect 96520 42400 96536 42464
rect 96600 42400 96616 42464
rect 96680 42400 96688 42464
rect 96368 41376 96688 42400
rect 96368 41312 96376 41376
rect 96440 41312 96456 41376
rect 96520 41312 96536 41376
rect 96600 41312 96616 41376
rect 96680 41312 96688 41376
rect 96368 40288 96688 41312
rect 96368 40224 96376 40288
rect 96440 40224 96456 40288
rect 96520 40224 96536 40288
rect 96600 40224 96616 40288
rect 96680 40224 96688 40288
rect 96368 39200 96688 40224
rect 96368 39136 96376 39200
rect 96440 39136 96456 39200
rect 96520 39136 96536 39200
rect 96600 39136 96616 39200
rect 96680 39136 96688 39200
rect 96368 38112 96688 39136
rect 96368 38048 96376 38112
rect 96440 38048 96456 38112
rect 96520 38048 96536 38112
rect 96600 38048 96616 38112
rect 96680 38048 96688 38112
rect 96368 37024 96688 38048
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 35936 96688 36960
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 34848 96688 35872
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 33760 96688 34784
rect 96368 33696 96376 33760
rect 96440 33696 96456 33760
rect 96520 33696 96536 33760
rect 96600 33696 96616 33760
rect 96680 33696 96688 33760
rect 96368 32672 96688 33696
rect 96368 32608 96376 32672
rect 96440 32608 96456 32672
rect 96520 32608 96536 32672
rect 96600 32608 96616 32672
rect 96680 32608 96688 32672
rect 96368 31584 96688 32608
rect 96368 31520 96376 31584
rect 96440 31520 96456 31584
rect 96520 31520 96536 31584
rect 96600 31520 96616 31584
rect 96680 31520 96688 31584
rect 96368 30496 96688 31520
rect 96368 30432 96376 30496
rect 96440 30432 96456 30496
rect 96520 30432 96536 30496
rect 96600 30432 96616 30496
rect 96680 30432 96688 30496
rect 96368 29408 96688 30432
rect 96368 29344 96376 29408
rect 96440 29344 96456 29408
rect 96520 29344 96536 29408
rect 96600 29344 96616 29408
rect 96680 29344 96688 29408
rect 96368 28320 96688 29344
rect 96368 28256 96376 28320
rect 96440 28256 96456 28320
rect 96520 28256 96536 28320
rect 96600 28256 96616 28320
rect 96680 28256 96688 28320
rect 96368 27232 96688 28256
rect 96368 27168 96376 27232
rect 96440 27168 96456 27232
rect 96520 27168 96536 27232
rect 96600 27168 96616 27232
rect 96680 27168 96688 27232
rect 96368 26144 96688 27168
rect 96368 26080 96376 26144
rect 96440 26080 96456 26144
rect 96520 26080 96536 26144
rect 96600 26080 96616 26144
rect 96680 26080 96688 26144
rect 96368 25056 96688 26080
rect 96368 24992 96376 25056
rect 96440 24992 96456 25056
rect 96520 24992 96536 25056
rect 96600 24992 96616 25056
rect 96680 24992 96688 25056
rect 96368 23968 96688 24992
rect 96368 23904 96376 23968
rect 96440 23904 96456 23968
rect 96520 23904 96536 23968
rect 96600 23904 96616 23968
rect 96680 23904 96688 23968
rect 96368 22880 96688 23904
rect 96368 22816 96376 22880
rect 96440 22816 96456 22880
rect 96520 22816 96536 22880
rect 96600 22816 96616 22880
rect 96680 22816 96688 22880
rect 96368 21792 96688 22816
rect 96368 21728 96376 21792
rect 96440 21728 96456 21792
rect 96520 21728 96536 21792
rect 96600 21728 96616 21792
rect 96680 21728 96688 21792
rect 96368 20704 96688 21728
rect 96368 20640 96376 20704
rect 96440 20640 96456 20704
rect 96520 20640 96536 20704
rect 96600 20640 96616 20704
rect 96680 20640 96688 20704
rect 96368 19616 96688 20640
rect 96368 19552 96376 19616
rect 96440 19552 96456 19616
rect 96520 19552 96536 19616
rect 96600 19552 96616 19616
rect 96680 19552 96688 19616
rect 96368 18528 96688 19552
rect 96368 18464 96376 18528
rect 96440 18464 96456 18528
rect 96520 18464 96536 18528
rect 96600 18464 96616 18528
rect 96680 18464 96688 18528
rect 96368 17440 96688 18464
rect 96368 17376 96376 17440
rect 96440 17376 96456 17440
rect 96520 17376 96536 17440
rect 96600 17376 96616 17440
rect 96680 17376 96688 17440
rect 96368 16352 96688 17376
rect 96368 16288 96376 16352
rect 96440 16288 96456 16352
rect 96520 16288 96536 16352
rect 96600 16288 96616 16352
rect 96680 16288 96688 16352
rect 96368 15264 96688 16288
rect 96368 15200 96376 15264
rect 96440 15200 96456 15264
rect 96520 15200 96536 15264
rect 96600 15200 96616 15264
rect 96680 15200 96688 15264
rect 96368 14176 96688 15200
rect 96368 14112 96376 14176
rect 96440 14112 96456 14176
rect 96520 14112 96536 14176
rect 96600 14112 96616 14176
rect 96680 14112 96688 14176
rect 96368 13088 96688 14112
rect 96368 13024 96376 13088
rect 96440 13024 96456 13088
rect 96520 13024 96536 13088
rect 96600 13024 96616 13088
rect 96680 13024 96688 13088
rect 96368 12000 96688 13024
rect 96368 11936 96376 12000
rect 96440 11936 96456 12000
rect 96520 11936 96536 12000
rect 96600 11936 96616 12000
rect 96680 11936 96688 12000
rect 96368 10912 96688 11936
rect 96368 10848 96376 10912
rect 96440 10848 96456 10912
rect 96520 10848 96536 10912
rect 96600 10848 96616 10912
rect 96680 10848 96688 10912
rect 96368 9824 96688 10848
rect 96368 9760 96376 9824
rect 96440 9760 96456 9824
rect 96520 9760 96536 9824
rect 96600 9760 96616 9824
rect 96680 9760 96688 9824
rect 96368 8736 96688 9760
rect 96368 8672 96376 8736
rect 96440 8672 96456 8736
rect 96520 8672 96536 8736
rect 96600 8672 96616 8736
rect 96680 8672 96688 8736
rect 96368 7648 96688 8672
rect 96368 7584 96376 7648
rect 96440 7584 96456 7648
rect 96520 7584 96536 7648
rect 96600 7584 96616 7648
rect 96680 7584 96688 7648
rect 96368 6560 96688 7584
rect 96368 6496 96376 6560
rect 96440 6496 96456 6560
rect 96520 6496 96536 6560
rect 96600 6496 96616 6560
rect 96680 6496 96688 6560
rect 96368 5472 96688 6496
rect 96368 5408 96376 5472
rect 96440 5408 96456 5472
rect 96520 5408 96536 5472
rect 96600 5408 96616 5472
rect 96680 5408 96688 5472
rect 96368 4384 96688 5408
rect 96368 4320 96376 4384
rect 96440 4320 96456 4384
rect 96520 4320 96536 4384
rect 96600 4320 96616 4384
rect 96680 4320 96688 4384
rect 96368 3296 96688 4320
rect 96368 3232 96376 3296
rect 96440 3232 96456 3296
rect 96520 3232 96536 3296
rect 96600 3232 96616 3296
rect 96680 3232 96688 3296
rect 96368 2208 96688 3232
rect 96368 2144 96376 2208
rect 96440 2144 96456 2208
rect 96520 2144 96536 2208
rect 96600 2144 96616 2208
rect 96680 2144 96688 2208
rect 97028 2176 97348 97376
rect 97688 2176 98008 97376
rect 96368 2128 96688 2144
<< labels >>
rlabel metal2 s 386 99200 442 100000 6 io_in[0]
port 0 nsew signal input
rlabel metal2 s 26422 99200 26478 100000 6 io_in[10]
port 1 nsew signal input
rlabel metal2 s 28998 99200 29054 100000 6 io_in[11]
port 2 nsew signal input
rlabel metal2 s 31666 99200 31722 100000 6 io_in[12]
port 3 nsew signal input
rlabel metal2 s 34242 99200 34298 100000 6 io_in[13]
port 4 nsew signal input
rlabel metal2 s 36818 99200 36874 100000 6 io_in[14]
port 5 nsew signal input
rlabel metal2 s 39486 99200 39542 100000 6 io_in[15]
port 6 nsew signal input
rlabel metal2 s 42062 99200 42118 100000 6 io_in[16]
port 7 nsew signal input
rlabel metal2 s 44730 99200 44786 100000 6 io_in[17]
port 8 nsew signal input
rlabel metal2 s 47306 99200 47362 100000 6 io_in[18]
port 9 nsew signal input
rlabel metal2 s 49882 99200 49938 100000 6 io_in[19]
port 10 nsew signal input
rlabel metal2 s 2962 99200 3018 100000 6 io_in[1]
port 11 nsew signal input
rlabel metal2 s 52550 99200 52606 100000 6 io_in[20]
port 12 nsew signal input
rlabel metal2 s 55126 99200 55182 100000 6 io_in[21]
port 13 nsew signal input
rlabel metal2 s 57702 99200 57758 100000 6 io_in[22]
port 14 nsew signal input
rlabel metal2 s 60370 99200 60426 100000 6 io_in[23]
port 15 nsew signal input
rlabel metal2 s 62946 99200 63002 100000 6 io_in[24]
port 16 nsew signal input
rlabel metal2 s 65522 99200 65578 100000 6 io_in[25]
port 17 nsew signal input
rlabel metal2 s 68190 99200 68246 100000 6 io_in[26]
port 18 nsew signal input
rlabel metal2 s 70766 99200 70822 100000 6 io_in[27]
port 19 nsew signal input
rlabel metal2 s 73342 99200 73398 100000 6 io_in[28]
port 20 nsew signal input
rlabel metal2 s 76010 99200 76066 100000 6 io_in[29]
port 21 nsew signal input
rlabel metal2 s 5538 99200 5594 100000 6 io_in[2]
port 22 nsew signal input
rlabel metal2 s 78586 99200 78642 100000 6 io_in[30]
port 23 nsew signal input
rlabel metal2 s 81254 99200 81310 100000 6 io_in[31]
port 24 nsew signal input
rlabel metal2 s 83830 99200 83886 100000 6 io_in[32]
port 25 nsew signal input
rlabel metal2 s 86406 99200 86462 100000 6 io_in[33]
port 26 nsew signal input
rlabel metal2 s 89074 99200 89130 100000 6 io_in[34]
port 27 nsew signal input
rlabel metal2 s 91650 99200 91706 100000 6 io_in[35]
port 28 nsew signal input
rlabel metal2 s 94226 99200 94282 100000 6 io_in[36]
port 29 nsew signal input
rlabel metal2 s 96894 99200 96950 100000 6 io_in[37]
port 30 nsew signal input
rlabel metal2 s 8206 99200 8262 100000 6 io_in[3]
port 31 nsew signal input
rlabel metal2 s 10782 99200 10838 100000 6 io_in[4]
port 32 nsew signal input
rlabel metal2 s 13358 99200 13414 100000 6 io_in[5]
port 33 nsew signal input
rlabel metal2 s 16026 99200 16082 100000 6 io_in[6]
port 34 nsew signal input
rlabel metal2 s 18602 99200 18658 100000 6 io_in[7]
port 35 nsew signal input
rlabel metal2 s 21178 99200 21234 100000 6 io_in[8]
port 36 nsew signal input
rlabel metal2 s 23846 99200 23902 100000 6 io_in[9]
port 37 nsew signal input
rlabel metal2 s 1214 99200 1270 100000 6 io_oeb[0]
port 38 nsew signal tristate
rlabel metal2 s 27342 99200 27398 100000 6 io_oeb[10]
port 39 nsew signal tristate
rlabel metal2 s 29918 99200 29974 100000 6 io_oeb[11]
port 40 nsew signal tristate
rlabel metal2 s 32494 99200 32550 100000 6 io_oeb[12]
port 41 nsew signal tristate
rlabel metal2 s 35162 99200 35218 100000 6 io_oeb[13]
port 42 nsew signal tristate
rlabel metal2 s 37738 99200 37794 100000 6 io_oeb[14]
port 43 nsew signal tristate
rlabel metal2 s 40314 99200 40370 100000 6 io_oeb[15]
port 44 nsew signal tristate
rlabel metal2 s 42982 99200 43038 100000 6 io_oeb[16]
port 45 nsew signal tristate
rlabel metal2 s 45558 99200 45614 100000 6 io_oeb[17]
port 46 nsew signal tristate
rlabel metal2 s 48134 99200 48190 100000 6 io_oeb[18]
port 47 nsew signal tristate
rlabel metal2 s 50802 99200 50858 100000 6 io_oeb[19]
port 48 nsew signal tristate
rlabel metal2 s 3790 99200 3846 100000 6 io_oeb[1]
port 49 nsew signal tristate
rlabel metal2 s 53378 99200 53434 100000 6 io_oeb[20]
port 50 nsew signal tristate
rlabel metal2 s 55954 99200 56010 100000 6 io_oeb[21]
port 51 nsew signal tristate
rlabel metal2 s 58622 99200 58678 100000 6 io_oeb[22]
port 52 nsew signal tristate
rlabel metal2 s 61198 99200 61254 100000 6 io_oeb[23]
port 53 nsew signal tristate
rlabel metal2 s 63866 99200 63922 100000 6 io_oeb[24]
port 54 nsew signal tristate
rlabel metal2 s 66442 99200 66498 100000 6 io_oeb[25]
port 55 nsew signal tristate
rlabel metal2 s 69018 99200 69074 100000 6 io_oeb[26]
port 56 nsew signal tristate
rlabel metal2 s 71686 99200 71742 100000 6 io_oeb[27]
port 57 nsew signal tristate
rlabel metal2 s 74262 99200 74318 100000 6 io_oeb[28]
port 58 nsew signal tristate
rlabel metal2 s 76838 99200 76894 100000 6 io_oeb[29]
port 59 nsew signal tristate
rlabel metal2 s 6458 99200 6514 100000 6 io_oeb[2]
port 60 nsew signal tristate
rlabel metal2 s 79506 99200 79562 100000 6 io_oeb[30]
port 61 nsew signal tristate
rlabel metal2 s 82082 99200 82138 100000 6 io_oeb[31]
port 62 nsew signal tristate
rlabel metal2 s 84658 99200 84714 100000 6 io_oeb[32]
port 63 nsew signal tristate
rlabel metal2 s 87326 99200 87382 100000 6 io_oeb[33]
port 64 nsew signal tristate
rlabel metal2 s 89902 99200 89958 100000 6 io_oeb[34]
port 65 nsew signal tristate
rlabel metal2 s 92478 99200 92534 100000 6 io_oeb[35]
port 66 nsew signal tristate
rlabel metal2 s 95146 99200 95202 100000 6 io_oeb[36]
port 67 nsew signal tristate
rlabel metal2 s 97722 99200 97778 100000 6 io_oeb[37]
port 68 nsew signal tristate
rlabel metal2 s 9034 99200 9090 100000 6 io_oeb[3]
port 69 nsew signal tristate
rlabel metal2 s 11610 99200 11666 100000 6 io_oeb[4]
port 70 nsew signal tristate
rlabel metal2 s 14278 99200 14334 100000 6 io_oeb[5]
port 71 nsew signal tristate
rlabel metal2 s 16854 99200 16910 100000 6 io_oeb[6]
port 72 nsew signal tristate
rlabel metal2 s 19430 99200 19486 100000 6 io_oeb[7]
port 73 nsew signal tristate
rlabel metal2 s 22098 99200 22154 100000 6 io_oeb[8]
port 74 nsew signal tristate
rlabel metal2 s 24674 99200 24730 100000 6 io_oeb[9]
port 75 nsew signal tristate
rlabel metal2 s 2042 99200 2098 100000 6 io_out[0]
port 76 nsew signal tristate
rlabel metal2 s 28170 99200 28226 100000 6 io_out[10]
port 77 nsew signal tristate
rlabel metal2 s 30746 99200 30802 100000 6 io_out[11]
port 78 nsew signal tristate
rlabel metal2 s 33414 99200 33470 100000 6 io_out[12]
port 79 nsew signal tristate
rlabel metal2 s 35990 99200 36046 100000 6 io_out[13]
port 80 nsew signal tristate
rlabel metal2 s 38566 99200 38622 100000 6 io_out[14]
port 81 nsew signal tristate
rlabel metal2 s 41234 99200 41290 100000 6 io_out[15]
port 82 nsew signal tristate
rlabel metal2 s 43810 99200 43866 100000 6 io_out[16]
port 83 nsew signal tristate
rlabel metal2 s 46386 99200 46442 100000 6 io_out[17]
port 84 nsew signal tristate
rlabel metal2 s 49054 99200 49110 100000 6 io_out[18]
port 85 nsew signal tristate
rlabel metal2 s 51630 99200 51686 100000 6 io_out[19]
port 86 nsew signal tristate
rlabel metal2 s 4710 99200 4766 100000 6 io_out[1]
port 87 nsew signal tristate
rlabel metal2 s 54298 99200 54354 100000 6 io_out[20]
port 88 nsew signal tristate
rlabel metal2 s 56874 99200 56930 100000 6 io_out[21]
port 89 nsew signal tristate
rlabel metal2 s 59450 99200 59506 100000 6 io_out[22]
port 90 nsew signal tristate
rlabel metal2 s 62118 99200 62174 100000 6 io_out[23]
port 91 nsew signal tristate
rlabel metal2 s 64694 99200 64750 100000 6 io_out[24]
port 92 nsew signal tristate
rlabel metal2 s 67270 99200 67326 100000 6 io_out[25]
port 93 nsew signal tristate
rlabel metal2 s 69938 99200 69994 100000 6 io_out[26]
port 94 nsew signal tristate
rlabel metal2 s 72514 99200 72570 100000 6 io_out[27]
port 95 nsew signal tristate
rlabel metal2 s 75090 99200 75146 100000 6 io_out[28]
port 96 nsew signal tristate
rlabel metal2 s 77758 99200 77814 100000 6 io_out[29]
port 97 nsew signal tristate
rlabel metal2 s 7286 99200 7342 100000 6 io_out[2]
port 98 nsew signal tristate
rlabel metal2 s 80334 99200 80390 100000 6 io_out[30]
port 99 nsew signal tristate
rlabel metal2 s 82910 99200 82966 100000 6 io_out[31]
port 100 nsew signal tristate
rlabel metal2 s 85578 99200 85634 100000 6 io_out[32]
port 101 nsew signal tristate
rlabel metal2 s 88154 99200 88210 100000 6 io_out[33]
port 102 nsew signal tristate
rlabel metal2 s 90822 99200 90878 100000 6 io_out[34]
port 103 nsew signal tristate
rlabel metal2 s 93398 99200 93454 100000 6 io_out[35]
port 104 nsew signal tristate
rlabel metal2 s 95974 99200 96030 100000 6 io_out[36]
port 105 nsew signal tristate
rlabel metal2 s 98642 99200 98698 100000 6 io_out[37]
port 106 nsew signal tristate
rlabel metal2 s 9862 99200 9918 100000 6 io_out[3]
port 107 nsew signal tristate
rlabel metal2 s 12530 99200 12586 100000 6 io_out[4]
port 108 nsew signal tristate
rlabel metal2 s 15106 99200 15162 100000 6 io_out[5]
port 109 nsew signal tristate
rlabel metal2 s 17774 99200 17830 100000 6 io_out[6]
port 110 nsew signal tristate
rlabel metal2 s 20350 99200 20406 100000 6 io_out[7]
port 111 nsew signal tristate
rlabel metal2 s 22926 99200 22982 100000 6 io_out[8]
port 112 nsew signal tristate
rlabel metal2 s 25594 99200 25650 100000 6 io_out[9]
port 113 nsew signal tristate
rlabel metal2 s 99654 0 99710 800 6 irq[0]
port 114 nsew signal tristate
rlabel metal2 s 99470 99200 99526 100000 6 irq[1]
port 115 nsew signal tristate
rlabel metal2 s 99838 0 99894 800 6 irq[2]
port 116 nsew signal tristate
rlabel metal2 s 21638 0 21694 800 6 la_data_in[0]
port 117 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[100]
port 118 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_data_in[101]
port 119 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[102]
port 120 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[103]
port 121 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[104]
port 122 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_data_in[105]
port 123 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[106]
port 124 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[107]
port 125 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[108]
port 126 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[109]
port 127 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[10]
port 128 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[110]
port 129 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_data_in[111]
port 130 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[112]
port 131 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[113]
port 132 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[114]
port 133 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[115]
port 134 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[116]
port 135 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[117]
port 136 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[118]
port 137 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[119]
port 138 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_in[11]
port 139 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[120]
port 140 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[121]
port 141 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[122]
port 142 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[123]
port 143 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[124]
port 144 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[125]
port 145 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[126]
port 146 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[127]
port 147 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in[12]
port 148 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[13]
port 149 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[14]
port 150 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in[15]
port 151 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_data_in[16]
port 152 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[17]
port 153 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[18]
port 154 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_data_in[19]
port 155 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[1]
port 156 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_data_in[20]
port 157 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[21]
port 158 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[22]
port 159 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_data_in[23]
port 160 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[24]
port 161 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[25]
port 162 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_in[26]
port 163 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[27]
port 164 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_data_in[28]
port 165 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[29]
port 166 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_data_in[2]
port 167 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[30]
port 168 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[31]
port 169 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[32]
port 170 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[33]
port 171 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[34]
port 172 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_data_in[35]
port 173 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[36]
port 174 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[37]
port 175 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[38]
port 176 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[39]
port 177 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[3]
port 178 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[40]
port 179 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[41]
port 180 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[42]
port 181 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[43]
port 182 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_data_in[44]
port 183 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[45]
port 184 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[46]
port 185 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[47]
port 186 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_data_in[48]
port 187 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[49]
port 188 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[4]
port 189 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_data_in[50]
port 190 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[51]
port 191 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[52]
port 192 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[53]
port 193 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[54]
port 194 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[55]
port 195 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[56]
port 196 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[57]
port 197 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[58]
port 198 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[59]
port 199 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 la_data_in[5]
port 200 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_data_in[60]
port 201 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[61]
port 202 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[62]
port 203 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[63]
port 204 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[64]
port 205 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[65]
port 206 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[66]
port 207 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_data_in[67]
port 208 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[68]
port 209 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[69]
port 210 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[6]
port 211 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[70]
port 212 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[71]
port 213 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_data_in[72]
port 214 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[73]
port 215 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[74]
port 216 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[75]
port 217 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[76]
port 218 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[77]
port 219 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[78]
port 220 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[79]
port 221 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[7]
port 222 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[80]
port 223 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[81]
port 224 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[82]
port 225 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[83]
port 226 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[84]
port 227 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[85]
port 228 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[86]
port 229 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[87]
port 230 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[88]
port 231 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[89]
port 232 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_data_in[8]
port 233 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[90]
port 234 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[91]
port 235 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[92]
port 236 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[93]
port 237 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[94]
port 238 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[95]
port 239 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[96]
port 240 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[97]
port 241 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[98]
port 242 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[99]
port 243 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[9]
port 244 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_out[0]
port 245 nsew signal tristate
rlabel metal2 s 82818 0 82874 800 6 la_data_out[100]
port 246 nsew signal tristate
rlabel metal2 s 83370 0 83426 800 6 la_data_out[101]
port 247 nsew signal tristate
rlabel metal2 s 84014 0 84070 800 6 la_data_out[102]
port 248 nsew signal tristate
rlabel metal2 s 84658 0 84714 800 6 la_data_out[103]
port 249 nsew signal tristate
rlabel metal2 s 85210 0 85266 800 6 la_data_out[104]
port 250 nsew signal tristate
rlabel metal2 s 85854 0 85910 800 6 la_data_out[105]
port 251 nsew signal tristate
rlabel metal2 s 86406 0 86462 800 6 la_data_out[106]
port 252 nsew signal tristate
rlabel metal2 s 87050 0 87106 800 6 la_data_out[107]
port 253 nsew signal tristate
rlabel metal2 s 87694 0 87750 800 6 la_data_out[108]
port 254 nsew signal tristate
rlabel metal2 s 88246 0 88302 800 6 la_data_out[109]
port 255 nsew signal tristate
rlabel metal2 s 27894 0 27950 800 6 la_data_out[10]
port 256 nsew signal tristate
rlabel metal2 s 88890 0 88946 800 6 la_data_out[110]
port 257 nsew signal tristate
rlabel metal2 s 89534 0 89590 800 6 la_data_out[111]
port 258 nsew signal tristate
rlabel metal2 s 90086 0 90142 800 6 la_data_out[112]
port 259 nsew signal tristate
rlabel metal2 s 90730 0 90786 800 6 la_data_out[113]
port 260 nsew signal tristate
rlabel metal2 s 91282 0 91338 800 6 la_data_out[114]
port 261 nsew signal tristate
rlabel metal2 s 91926 0 91982 800 6 la_data_out[115]
port 262 nsew signal tristate
rlabel metal2 s 92570 0 92626 800 6 la_data_out[116]
port 263 nsew signal tristate
rlabel metal2 s 93122 0 93178 800 6 la_data_out[117]
port 264 nsew signal tristate
rlabel metal2 s 93766 0 93822 800 6 la_data_out[118]
port 265 nsew signal tristate
rlabel metal2 s 94410 0 94466 800 6 la_data_out[119]
port 266 nsew signal tristate
rlabel metal2 s 28538 0 28594 800 6 la_data_out[11]
port 267 nsew signal tristate
rlabel metal2 s 94962 0 95018 800 6 la_data_out[120]
port 268 nsew signal tristate
rlabel metal2 s 95606 0 95662 800 6 la_data_out[121]
port 269 nsew signal tristate
rlabel metal2 s 96250 0 96306 800 6 la_data_out[122]
port 270 nsew signal tristate
rlabel metal2 s 96802 0 96858 800 6 la_data_out[123]
port 271 nsew signal tristate
rlabel metal2 s 97446 0 97502 800 6 la_data_out[124]
port 272 nsew signal tristate
rlabel metal2 s 97998 0 98054 800 6 la_data_out[125]
port 273 nsew signal tristate
rlabel metal2 s 98642 0 98698 800 6 la_data_out[126]
port 274 nsew signal tristate
rlabel metal2 s 99286 0 99342 800 6 la_data_out[127]
port 275 nsew signal tristate
rlabel metal2 s 29090 0 29146 800 6 la_data_out[12]
port 276 nsew signal tristate
rlabel metal2 s 29734 0 29790 800 6 la_data_out[13]
port 277 nsew signal tristate
rlabel metal2 s 30378 0 30434 800 6 la_data_out[14]
port 278 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 la_data_out[15]
port 279 nsew signal tristate
rlabel metal2 s 31574 0 31630 800 6 la_data_out[16]
port 280 nsew signal tristate
rlabel metal2 s 32218 0 32274 800 6 la_data_out[17]
port 281 nsew signal tristate
rlabel metal2 s 32770 0 32826 800 6 la_data_out[18]
port 282 nsew signal tristate
rlabel metal2 s 33414 0 33470 800 6 la_data_out[19]
port 283 nsew signal tristate
rlabel metal2 s 22466 0 22522 800 6 la_data_out[1]
port 284 nsew signal tristate
rlabel metal2 s 33966 0 34022 800 6 la_data_out[20]
port 285 nsew signal tristate
rlabel metal2 s 34610 0 34666 800 6 la_data_out[21]
port 286 nsew signal tristate
rlabel metal2 s 35254 0 35310 800 6 la_data_out[22]
port 287 nsew signal tristate
rlabel metal2 s 35806 0 35862 800 6 la_data_out[23]
port 288 nsew signal tristate
rlabel metal2 s 36450 0 36506 800 6 la_data_out[24]
port 289 nsew signal tristate
rlabel metal2 s 37094 0 37150 800 6 la_data_out[25]
port 290 nsew signal tristate
rlabel metal2 s 37646 0 37702 800 6 la_data_out[26]
port 291 nsew signal tristate
rlabel metal2 s 38290 0 38346 800 6 la_data_out[27]
port 292 nsew signal tristate
rlabel metal2 s 38842 0 38898 800 6 la_data_out[28]
port 293 nsew signal tristate
rlabel metal2 s 39486 0 39542 800 6 la_data_out[29]
port 294 nsew signal tristate
rlabel metal2 s 23018 0 23074 800 6 la_data_out[2]
port 295 nsew signal tristate
rlabel metal2 s 40130 0 40186 800 6 la_data_out[30]
port 296 nsew signal tristate
rlabel metal2 s 40682 0 40738 800 6 la_data_out[31]
port 297 nsew signal tristate
rlabel metal2 s 41326 0 41382 800 6 la_data_out[32]
port 298 nsew signal tristate
rlabel metal2 s 41970 0 42026 800 6 la_data_out[33]
port 299 nsew signal tristate
rlabel metal2 s 42522 0 42578 800 6 la_data_out[34]
port 300 nsew signal tristate
rlabel metal2 s 43166 0 43222 800 6 la_data_out[35]
port 301 nsew signal tristate
rlabel metal2 s 43810 0 43866 800 6 la_data_out[36]
port 302 nsew signal tristate
rlabel metal2 s 44362 0 44418 800 6 la_data_out[37]
port 303 nsew signal tristate
rlabel metal2 s 45006 0 45062 800 6 la_data_out[38]
port 304 nsew signal tristate
rlabel metal2 s 45558 0 45614 800 6 la_data_out[39]
port 305 nsew signal tristate
rlabel metal2 s 23662 0 23718 800 6 la_data_out[3]
port 306 nsew signal tristate
rlabel metal2 s 46202 0 46258 800 6 la_data_out[40]
port 307 nsew signal tristate
rlabel metal2 s 46846 0 46902 800 6 la_data_out[41]
port 308 nsew signal tristate
rlabel metal2 s 47398 0 47454 800 6 la_data_out[42]
port 309 nsew signal tristate
rlabel metal2 s 48042 0 48098 800 6 la_data_out[43]
port 310 nsew signal tristate
rlabel metal2 s 48686 0 48742 800 6 la_data_out[44]
port 311 nsew signal tristate
rlabel metal2 s 49238 0 49294 800 6 la_data_out[45]
port 312 nsew signal tristate
rlabel metal2 s 49882 0 49938 800 6 la_data_out[46]
port 313 nsew signal tristate
rlabel metal2 s 50434 0 50490 800 6 la_data_out[47]
port 314 nsew signal tristate
rlabel metal2 s 51078 0 51134 800 6 la_data_out[48]
port 315 nsew signal tristate
rlabel metal2 s 51722 0 51778 800 6 la_data_out[49]
port 316 nsew signal tristate
rlabel metal2 s 24214 0 24270 800 6 la_data_out[4]
port 317 nsew signal tristate
rlabel metal2 s 52274 0 52330 800 6 la_data_out[50]
port 318 nsew signal tristate
rlabel metal2 s 52918 0 52974 800 6 la_data_out[51]
port 319 nsew signal tristate
rlabel metal2 s 53562 0 53618 800 6 la_data_out[52]
port 320 nsew signal tristate
rlabel metal2 s 54114 0 54170 800 6 la_data_out[53]
port 321 nsew signal tristate
rlabel metal2 s 54758 0 54814 800 6 la_data_out[54]
port 322 nsew signal tristate
rlabel metal2 s 55310 0 55366 800 6 la_data_out[55]
port 323 nsew signal tristate
rlabel metal2 s 55954 0 56010 800 6 la_data_out[56]
port 324 nsew signal tristate
rlabel metal2 s 56598 0 56654 800 6 la_data_out[57]
port 325 nsew signal tristate
rlabel metal2 s 57150 0 57206 800 6 la_data_out[58]
port 326 nsew signal tristate
rlabel metal2 s 57794 0 57850 800 6 la_data_out[59]
port 327 nsew signal tristate
rlabel metal2 s 24858 0 24914 800 6 la_data_out[5]
port 328 nsew signal tristate
rlabel metal2 s 58438 0 58494 800 6 la_data_out[60]
port 329 nsew signal tristate
rlabel metal2 s 58990 0 59046 800 6 la_data_out[61]
port 330 nsew signal tristate
rlabel metal2 s 59634 0 59690 800 6 la_data_out[62]
port 331 nsew signal tristate
rlabel metal2 s 60186 0 60242 800 6 la_data_out[63]
port 332 nsew signal tristate
rlabel metal2 s 60830 0 60886 800 6 la_data_out[64]
port 333 nsew signal tristate
rlabel metal2 s 61474 0 61530 800 6 la_data_out[65]
port 334 nsew signal tristate
rlabel metal2 s 62026 0 62082 800 6 la_data_out[66]
port 335 nsew signal tristate
rlabel metal2 s 62670 0 62726 800 6 la_data_out[67]
port 336 nsew signal tristate
rlabel metal2 s 63314 0 63370 800 6 la_data_out[68]
port 337 nsew signal tristate
rlabel metal2 s 63866 0 63922 800 6 la_data_out[69]
port 338 nsew signal tristate
rlabel metal2 s 25502 0 25558 800 6 la_data_out[6]
port 339 nsew signal tristate
rlabel metal2 s 64510 0 64566 800 6 la_data_out[70]
port 340 nsew signal tristate
rlabel metal2 s 65062 0 65118 800 6 la_data_out[71]
port 341 nsew signal tristate
rlabel metal2 s 65706 0 65762 800 6 la_data_out[72]
port 342 nsew signal tristate
rlabel metal2 s 66350 0 66406 800 6 la_data_out[73]
port 343 nsew signal tristate
rlabel metal2 s 66902 0 66958 800 6 la_data_out[74]
port 344 nsew signal tristate
rlabel metal2 s 67546 0 67602 800 6 la_data_out[75]
port 345 nsew signal tristate
rlabel metal2 s 68190 0 68246 800 6 la_data_out[76]
port 346 nsew signal tristate
rlabel metal2 s 68742 0 68798 800 6 la_data_out[77]
port 347 nsew signal tristate
rlabel metal2 s 69386 0 69442 800 6 la_data_out[78]
port 348 nsew signal tristate
rlabel metal2 s 70030 0 70086 800 6 la_data_out[79]
port 349 nsew signal tristate
rlabel metal2 s 26054 0 26110 800 6 la_data_out[7]
port 350 nsew signal tristate
rlabel metal2 s 70582 0 70638 800 6 la_data_out[80]
port 351 nsew signal tristate
rlabel metal2 s 71226 0 71282 800 6 la_data_out[81]
port 352 nsew signal tristate
rlabel metal2 s 71778 0 71834 800 6 la_data_out[82]
port 353 nsew signal tristate
rlabel metal2 s 72422 0 72478 800 6 la_data_out[83]
port 354 nsew signal tristate
rlabel metal2 s 73066 0 73122 800 6 la_data_out[84]
port 355 nsew signal tristate
rlabel metal2 s 73618 0 73674 800 6 la_data_out[85]
port 356 nsew signal tristate
rlabel metal2 s 74262 0 74318 800 6 la_data_out[86]
port 357 nsew signal tristate
rlabel metal2 s 74906 0 74962 800 6 la_data_out[87]
port 358 nsew signal tristate
rlabel metal2 s 75458 0 75514 800 6 la_data_out[88]
port 359 nsew signal tristate
rlabel metal2 s 76102 0 76158 800 6 la_data_out[89]
port 360 nsew signal tristate
rlabel metal2 s 26698 0 26754 800 6 la_data_out[8]
port 361 nsew signal tristate
rlabel metal2 s 76654 0 76710 800 6 la_data_out[90]
port 362 nsew signal tristate
rlabel metal2 s 77298 0 77354 800 6 la_data_out[91]
port 363 nsew signal tristate
rlabel metal2 s 77942 0 77998 800 6 la_data_out[92]
port 364 nsew signal tristate
rlabel metal2 s 78494 0 78550 800 6 la_data_out[93]
port 365 nsew signal tristate
rlabel metal2 s 79138 0 79194 800 6 la_data_out[94]
port 366 nsew signal tristate
rlabel metal2 s 79782 0 79838 800 6 la_data_out[95]
port 367 nsew signal tristate
rlabel metal2 s 80334 0 80390 800 6 la_data_out[96]
port 368 nsew signal tristate
rlabel metal2 s 80978 0 81034 800 6 la_data_out[97]
port 369 nsew signal tristate
rlabel metal2 s 81530 0 81586 800 6 la_data_out[98]
port 370 nsew signal tristate
rlabel metal2 s 82174 0 82230 800 6 la_data_out[99]
port 371 nsew signal tristate
rlabel metal2 s 27342 0 27398 800 6 la_data_out[9]
port 372 nsew signal tristate
rlabel metal2 s 22006 0 22062 800 6 la_oenb[0]
port 373 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[100]
port 374 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[101]
port 375 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[102]
port 376 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_oenb[103]
port 377 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[104]
port 378 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[105]
port 379 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[106]
port 380 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[107]
port 381 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[108]
port 382 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[109]
port 383 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[10]
port 384 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oenb[110]
port 385 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[111]
port 386 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[112]
port 387 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[113]
port 388 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[114]
port 389 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[115]
port 390 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[116]
port 391 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[117]
port 392 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[118]
port 393 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[119]
port 394 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[11]
port 395 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[120]
port 396 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[121]
port 397 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[122]
port 398 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[123]
port 399 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[124]
port 400 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_oenb[125]
port 401 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[126]
port 402 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[127]
port 403 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[12]
port 404 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[13]
port 405 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_oenb[14]
port 406 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_oenb[15]
port 407 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_oenb[16]
port 408 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_oenb[17]
port 409 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[18]
port 410 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_oenb[19]
port 411 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_oenb[1]
port 412 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_oenb[20]
port 413 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_oenb[21]
port 414 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_oenb[22]
port 415 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[23]
port 416 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_oenb[24]
port 417 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_oenb[25]
port 418 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[26]
port 419 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_oenb[27]
port 420 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[28]
port 421 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_oenb[29]
port 422 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 la_oenb[2]
port 423 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_oenb[30]
port 424 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[31]
port 425 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_oenb[32]
port 426 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_oenb[33]
port 427 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[34]
port 428 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[35]
port 429 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[36]
port 430 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[37]
port 431 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[38]
port 432 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[39]
port 433 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_oenb[3]
port 434 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[40]
port 435 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[41]
port 436 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[42]
port 437 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[43]
port 438 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[44]
port 439 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_oenb[45]
port 440 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_oenb[46]
port 441 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[47]
port 442 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[48]
port 443 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[49]
port 444 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_oenb[4]
port 445 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[50]
port 446 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[51]
port 447 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[52]
port 448 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_oenb[53]
port 449 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[54]
port 450 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[55]
port 451 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[56]
port 452 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[57]
port 453 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[58]
port 454 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_oenb[59]
port 455 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_oenb[5]
port 456 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[60]
port 457 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[61]
port 458 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[62]
port 459 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[63]
port 460 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[64]
port 461 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[65]
port 462 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oenb[66]
port 463 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[67]
port 464 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[68]
port 465 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_oenb[69]
port 466 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_oenb[6]
port 467 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[70]
port 468 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oenb[71]
port 469 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[72]
port 470 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[73]
port 471 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[74]
port 472 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[75]
port 473 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[76]
port 474 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[77]
port 475 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oenb[78]
port 476 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[79]
port 477 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[7]
port 478 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[80]
port 479 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[81]
port 480 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[82]
port 481 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_oenb[83]
port 482 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oenb[84]
port 483 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[85]
port 484 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_oenb[86]
port 485 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[87]
port 486 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[88]
port 487 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[89]
port 488 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_oenb[8]
port 489 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[90]
port 490 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_oenb[91]
port 491 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[92]
port 492 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[93]
port 493 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[94]
port 494 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[95]
port 495 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[96]
port 496 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_oenb[97]
port 497 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[98]
port 498 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[99]
port 499 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[9]
port 500 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 user_clock2
port 501 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 504 nsew signal tristate
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 570 nsew signal tristate
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[10]
port 571 nsew signal tristate
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[11]
port 572 nsew signal tristate
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[12]
port 573 nsew signal tristate
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[13]
port 574 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[14]
port 575 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[15]
port 576 nsew signal tristate
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[16]
port 577 nsew signal tristate
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[17]
port 578 nsew signal tristate
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[18]
port 579 nsew signal tristate
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[19]
port 580 nsew signal tristate
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[1]
port 581 nsew signal tristate
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[20]
port 582 nsew signal tristate
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[21]
port 583 nsew signal tristate
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[22]
port 584 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[23]
port 585 nsew signal tristate
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[24]
port 586 nsew signal tristate
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[25]
port 587 nsew signal tristate
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[26]
port 588 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[27]
port 589 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[28]
port 590 nsew signal tristate
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[29]
port 591 nsew signal tristate
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[2]
port 592 nsew signal tristate
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[30]
port 593 nsew signal tristate
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[31]
port 594 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[3]
port 595 nsew signal tristate
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[4]
port 596 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[5]
port 597 nsew signal tristate
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[6]
port 598 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[7]
port 599 nsew signal tristate
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[8]
port 600 nsew signal tristate
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[9]
port 601 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 612 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 613 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 97028 2176 97348 97376 6 vccd2
port 615 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 97376 6 vccd2
port 616 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 97376 6 vccd2
port 617 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 97376 6 vccd2
port 618 nsew power bidirectional
rlabel metal4 s 81668 2176 81988 97376 6 vssd2
port 619 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 97376 6 vssd2
port 620 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 97376 6 vssd2
port 621 nsew ground bidirectional
rlabel metal4 s 97688 2176 98008 97376 6 vdda1
port 622 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 97376 6 vdda1
port 623 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 97376 6 vdda1
port 624 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 97376 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 82328 2176 82648 97376 6 vssa1
port 626 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 97376 6 vssa1
port 627 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 97376 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 67628 2176 67948 97376 6 vdda2
port 629 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 97376 6 vdda2
port 630 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 97376 6 vdda2
port 631 nsew power bidirectional
rlabel metal4 s 82988 2176 83308 97376 6 vssa2
port 632 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 97376 6 vssa2
port 633 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 97376 6 vssa2
port 634 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 100000
<< end >>
