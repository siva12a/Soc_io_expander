magic
tech sky130A
magscale 1 2
timestamp 1623855685
<< obsli1 >>
rect 1409 2261 98227 97291
<< obsm1 >>
rect 106 1164 99898 97640
<< metal2 >>
rect 386 99200 442 100000
rect 1214 99200 1270 100000
rect 2042 99200 2098 100000
rect 2962 99200 3018 100000
rect 3790 99200 3846 100000
rect 4710 99200 4766 100000
rect 5538 99200 5594 100000
rect 6458 99200 6514 100000
rect 7286 99200 7342 100000
rect 8206 99200 8262 100000
rect 9034 99200 9090 100000
rect 9862 99200 9918 100000
rect 10782 99200 10838 100000
rect 11610 99200 11666 100000
rect 12530 99200 12586 100000
rect 13358 99200 13414 100000
rect 14278 99200 14334 100000
rect 15106 99200 15162 100000
rect 16026 99200 16082 100000
rect 16854 99200 16910 100000
rect 17774 99200 17830 100000
rect 18602 99200 18658 100000
rect 19430 99200 19486 100000
rect 20350 99200 20406 100000
rect 21178 99200 21234 100000
rect 22098 99200 22154 100000
rect 22926 99200 22982 100000
rect 23846 99200 23902 100000
rect 24674 99200 24730 100000
rect 25594 99200 25650 100000
rect 26422 99200 26478 100000
rect 27342 99200 27398 100000
rect 28170 99200 28226 100000
rect 28998 99200 29054 100000
rect 29918 99200 29974 100000
rect 30746 99200 30802 100000
rect 31666 99200 31722 100000
rect 32494 99200 32550 100000
rect 33414 99200 33470 100000
rect 34242 99200 34298 100000
rect 35162 99200 35218 100000
rect 35990 99200 36046 100000
rect 36818 99200 36874 100000
rect 37738 99200 37794 100000
rect 38566 99200 38622 100000
rect 39486 99200 39542 100000
rect 40314 99200 40370 100000
rect 41234 99200 41290 100000
rect 42062 99200 42118 100000
rect 42982 99200 43038 100000
rect 43810 99200 43866 100000
rect 44730 99200 44786 100000
rect 45558 99200 45614 100000
rect 46386 99200 46442 100000
rect 47306 99200 47362 100000
rect 48134 99200 48190 100000
rect 49054 99200 49110 100000
rect 49882 99200 49938 100000
rect 50802 99200 50858 100000
rect 51630 99200 51686 100000
rect 52550 99200 52606 100000
rect 53378 99200 53434 100000
rect 54298 99200 54354 100000
rect 55126 99200 55182 100000
rect 55954 99200 56010 100000
rect 56874 99200 56930 100000
rect 57702 99200 57758 100000
rect 58622 99200 58678 100000
rect 59450 99200 59506 100000
rect 60370 99200 60426 100000
rect 61198 99200 61254 100000
rect 62118 99200 62174 100000
rect 62946 99200 63002 100000
rect 63866 99200 63922 100000
rect 64694 99200 64750 100000
rect 65522 99200 65578 100000
rect 66442 99200 66498 100000
rect 67270 99200 67326 100000
rect 68190 99200 68246 100000
rect 69018 99200 69074 100000
rect 69938 99200 69994 100000
rect 70766 99200 70822 100000
rect 71686 99200 71742 100000
rect 72514 99200 72570 100000
rect 73342 99200 73398 100000
rect 74262 99200 74318 100000
rect 75090 99200 75146 100000
rect 76010 99200 76066 100000
rect 76838 99200 76894 100000
rect 77758 99200 77814 100000
rect 78586 99200 78642 100000
rect 79506 99200 79562 100000
rect 80334 99200 80390 100000
rect 81254 99200 81310 100000
rect 82082 99200 82138 100000
rect 82910 99200 82966 100000
rect 83830 99200 83886 100000
rect 84658 99200 84714 100000
rect 85578 99200 85634 100000
rect 86406 99200 86462 100000
rect 87326 99200 87382 100000
rect 88154 99200 88210 100000
rect 89074 99200 89130 100000
rect 89902 99200 89958 100000
rect 90822 99200 90878 100000
rect 91650 99200 91706 100000
rect 92478 99200 92534 100000
rect 93398 99200 93454 100000
rect 94226 99200 94282 100000
rect 95146 99200 95202 100000
rect 95974 99200 96030 100000
rect 96894 99200 96950 100000
rect 97722 99200 97778 100000
rect 98642 99200 98698 100000
rect 99470 99200 99526 100000
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 13910 0 13966 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19338 0 19394 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36450 0 36506 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38658 0 38714 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40130 0 40186 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62026 0 62082 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63498 0 63554 800
rect 63682 0 63738 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65338 0 65394 800
rect 65522 0 65578 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67546 0 67602 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70766 0 70822 800
rect 71042 0 71098 800
rect 71226 0 71282 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73250 0 73306 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73802 0 73858 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74906 0 74962 800
rect 75090 0 75146 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76286 0 76342 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78770 0 78826 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81346 0 81402 800
rect 81530 0 81586 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83002 0 83058 800
rect 83186 0 83242 800
rect 83370 0 83426 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85026 0 85082 800
rect 85210 0 85266 800
rect 85394 0 85450 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88522 0 88578 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89258 0 89314 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 92938 0 92994 800
rect 93122 0 93178 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95146 0 95202 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< obsm2 >>
rect 112 99144 330 99200
rect 498 99144 1158 99200
rect 1326 99144 1986 99200
rect 2154 99144 2906 99200
rect 3074 99144 3734 99200
rect 3902 99144 4654 99200
rect 4822 99144 5482 99200
rect 5650 99144 6402 99200
rect 6570 99144 7230 99200
rect 7398 99144 8150 99200
rect 8318 99144 8978 99200
rect 9146 99144 9806 99200
rect 9974 99144 10726 99200
rect 10894 99144 11554 99200
rect 11722 99144 12474 99200
rect 12642 99144 13302 99200
rect 13470 99144 14222 99200
rect 14390 99144 15050 99200
rect 15218 99144 15970 99200
rect 16138 99144 16798 99200
rect 16966 99144 17718 99200
rect 17886 99144 18546 99200
rect 18714 99144 19374 99200
rect 19542 99144 20294 99200
rect 20462 99144 21122 99200
rect 21290 99144 22042 99200
rect 22210 99144 22870 99200
rect 23038 99144 23790 99200
rect 23958 99144 24618 99200
rect 24786 99144 25538 99200
rect 25706 99144 26366 99200
rect 26534 99144 27286 99200
rect 27454 99144 28114 99200
rect 28282 99144 28942 99200
rect 29110 99144 29862 99200
rect 30030 99144 30690 99200
rect 30858 99144 31610 99200
rect 31778 99144 32438 99200
rect 32606 99144 33358 99200
rect 33526 99144 34186 99200
rect 34354 99144 35106 99200
rect 35274 99144 35934 99200
rect 36102 99144 36762 99200
rect 36930 99144 37682 99200
rect 37850 99144 38510 99200
rect 38678 99144 39430 99200
rect 39598 99144 40258 99200
rect 40426 99144 41178 99200
rect 41346 99144 42006 99200
rect 42174 99144 42926 99200
rect 43094 99144 43754 99200
rect 43922 99144 44674 99200
rect 44842 99144 45502 99200
rect 45670 99144 46330 99200
rect 46498 99144 47250 99200
rect 47418 99144 48078 99200
rect 48246 99144 48998 99200
rect 49166 99144 49826 99200
rect 49994 99144 50746 99200
rect 50914 99144 51574 99200
rect 51742 99144 52494 99200
rect 52662 99144 53322 99200
rect 53490 99144 54242 99200
rect 54410 99144 55070 99200
rect 55238 99144 55898 99200
rect 56066 99144 56818 99200
rect 56986 99144 57646 99200
rect 57814 99144 58566 99200
rect 58734 99144 59394 99200
rect 59562 99144 60314 99200
rect 60482 99144 61142 99200
rect 61310 99144 62062 99200
rect 62230 99144 62890 99200
rect 63058 99144 63810 99200
rect 63978 99144 64638 99200
rect 64806 99144 65466 99200
rect 65634 99144 66386 99200
rect 66554 99144 67214 99200
rect 67382 99144 68134 99200
rect 68302 99144 68962 99200
rect 69130 99144 69882 99200
rect 70050 99144 70710 99200
rect 70878 99144 71630 99200
rect 71798 99144 72458 99200
rect 72626 99144 73286 99200
rect 73454 99144 74206 99200
rect 74374 99144 75034 99200
rect 75202 99144 75954 99200
rect 76122 99144 76782 99200
rect 76950 99144 77702 99200
rect 77870 99144 78530 99200
rect 78698 99144 79450 99200
rect 79618 99144 80278 99200
rect 80446 99144 81198 99200
rect 81366 99144 82026 99200
rect 82194 99144 82854 99200
rect 83022 99144 83774 99200
rect 83942 99144 84602 99200
rect 84770 99144 85522 99200
rect 85690 99144 86350 99200
rect 86518 99144 87270 99200
rect 87438 99144 88098 99200
rect 88266 99144 89018 99200
rect 89186 99144 89846 99200
rect 90014 99144 90766 99200
rect 90934 99144 91594 99200
rect 91762 99144 92422 99200
rect 92590 99144 93342 99200
rect 93510 99144 94170 99200
rect 94338 99144 95090 99200
rect 95258 99144 95918 99200
rect 96086 99144 96838 99200
rect 97006 99144 97666 99200
rect 97834 99144 98586 99200
rect 98754 99144 99414 99200
rect 99582 99144 99892 99200
rect 112 856 99892 99144
rect 222 800 238 856
rect 406 800 422 856
rect 590 800 606 856
rect 774 800 790 856
rect 958 800 1066 856
rect 1234 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1618 856
rect 1786 800 1802 856
rect 1970 800 2078 856
rect 2246 800 2262 856
rect 2430 800 2446 856
rect 2614 800 2630 856
rect 2798 800 2814 856
rect 2982 800 3090 856
rect 3258 800 3274 856
rect 3442 800 3458 856
rect 3626 800 3642 856
rect 3810 800 3826 856
rect 3994 800 4102 856
rect 4270 800 4286 856
rect 4454 800 4470 856
rect 4638 800 4654 856
rect 4822 800 4930 856
rect 5098 800 5114 856
rect 5282 800 5298 856
rect 5466 800 5482 856
rect 5650 800 5666 856
rect 5834 800 5942 856
rect 6110 800 6126 856
rect 6294 800 6310 856
rect 6478 800 6494 856
rect 6662 800 6678 856
rect 6846 800 6954 856
rect 7122 800 7138 856
rect 7306 800 7322 856
rect 7490 800 7506 856
rect 7674 800 7690 856
rect 7858 800 7966 856
rect 8134 800 8150 856
rect 8318 800 8334 856
rect 8502 800 8518 856
rect 8686 800 8794 856
rect 8962 800 8978 856
rect 9146 800 9162 856
rect 9330 800 9346 856
rect 9514 800 9530 856
rect 9698 800 9806 856
rect 9974 800 9990 856
rect 10158 800 10174 856
rect 10342 800 10358 856
rect 10526 800 10542 856
rect 10710 800 10818 856
rect 10986 800 11002 856
rect 11170 800 11186 856
rect 11354 800 11370 856
rect 11538 800 11554 856
rect 11722 800 11830 856
rect 11998 800 12014 856
rect 12182 800 12198 856
rect 12366 800 12382 856
rect 12550 800 12566 856
rect 12734 800 12842 856
rect 13010 800 13026 856
rect 13194 800 13210 856
rect 13378 800 13394 856
rect 13562 800 13670 856
rect 13838 800 13854 856
rect 14022 800 14038 856
rect 14206 800 14222 856
rect 14390 800 14406 856
rect 14574 800 14682 856
rect 14850 800 14866 856
rect 15034 800 15050 856
rect 15218 800 15234 856
rect 15402 800 15418 856
rect 15586 800 15694 856
rect 15862 800 15878 856
rect 16046 800 16062 856
rect 16230 800 16246 856
rect 16414 800 16430 856
rect 16598 800 16706 856
rect 16874 800 16890 856
rect 17058 800 17074 856
rect 17242 800 17258 856
rect 17426 800 17534 856
rect 17702 800 17718 856
rect 17886 800 17902 856
rect 18070 800 18086 856
rect 18254 800 18270 856
rect 18438 800 18546 856
rect 18714 800 18730 856
rect 18898 800 18914 856
rect 19082 800 19098 856
rect 19266 800 19282 856
rect 19450 800 19558 856
rect 19726 800 19742 856
rect 19910 800 19926 856
rect 20094 800 20110 856
rect 20278 800 20294 856
rect 20462 800 20570 856
rect 20738 800 20754 856
rect 20922 800 20938 856
rect 21106 800 21122 856
rect 21290 800 21306 856
rect 21474 800 21582 856
rect 21750 800 21766 856
rect 21934 800 21950 856
rect 22118 800 22134 856
rect 22302 800 22410 856
rect 22578 800 22594 856
rect 22762 800 22778 856
rect 22946 800 22962 856
rect 23130 800 23146 856
rect 23314 800 23422 856
rect 23590 800 23606 856
rect 23774 800 23790 856
rect 23958 800 23974 856
rect 24142 800 24158 856
rect 24326 800 24434 856
rect 24602 800 24618 856
rect 24786 800 24802 856
rect 24970 800 24986 856
rect 25154 800 25170 856
rect 25338 800 25446 856
rect 25614 800 25630 856
rect 25798 800 25814 856
rect 25982 800 25998 856
rect 26166 800 26274 856
rect 26442 800 26458 856
rect 26626 800 26642 856
rect 26810 800 26826 856
rect 26994 800 27010 856
rect 27178 800 27286 856
rect 27454 800 27470 856
rect 27638 800 27654 856
rect 27822 800 27838 856
rect 28006 800 28022 856
rect 28190 800 28298 856
rect 28466 800 28482 856
rect 28650 800 28666 856
rect 28834 800 28850 856
rect 29018 800 29034 856
rect 29202 800 29310 856
rect 29478 800 29494 856
rect 29662 800 29678 856
rect 29846 800 29862 856
rect 30030 800 30046 856
rect 30214 800 30322 856
rect 30490 800 30506 856
rect 30674 800 30690 856
rect 30858 800 30874 856
rect 31042 800 31150 856
rect 31318 800 31334 856
rect 31502 800 31518 856
rect 31686 800 31702 856
rect 31870 800 31886 856
rect 32054 800 32162 856
rect 32330 800 32346 856
rect 32514 800 32530 856
rect 32698 800 32714 856
rect 32882 800 32898 856
rect 33066 800 33174 856
rect 33342 800 33358 856
rect 33526 800 33542 856
rect 33710 800 33726 856
rect 33894 800 33910 856
rect 34078 800 34186 856
rect 34354 800 34370 856
rect 34538 800 34554 856
rect 34722 800 34738 856
rect 34906 800 35014 856
rect 35182 800 35198 856
rect 35366 800 35382 856
rect 35550 800 35566 856
rect 35734 800 35750 856
rect 35918 800 36026 856
rect 36194 800 36210 856
rect 36378 800 36394 856
rect 36562 800 36578 856
rect 36746 800 36762 856
rect 36930 800 37038 856
rect 37206 800 37222 856
rect 37390 800 37406 856
rect 37574 800 37590 856
rect 37758 800 37774 856
rect 37942 800 38050 856
rect 38218 800 38234 856
rect 38402 800 38418 856
rect 38586 800 38602 856
rect 38770 800 38786 856
rect 38954 800 39062 856
rect 39230 800 39246 856
rect 39414 800 39430 856
rect 39598 800 39614 856
rect 39782 800 39890 856
rect 40058 800 40074 856
rect 40242 800 40258 856
rect 40426 800 40442 856
rect 40610 800 40626 856
rect 40794 800 40902 856
rect 41070 800 41086 856
rect 41254 800 41270 856
rect 41438 800 41454 856
rect 41622 800 41638 856
rect 41806 800 41914 856
rect 42082 800 42098 856
rect 42266 800 42282 856
rect 42450 800 42466 856
rect 42634 800 42650 856
rect 42818 800 42926 856
rect 43094 800 43110 856
rect 43278 800 43294 856
rect 43462 800 43478 856
rect 43646 800 43754 856
rect 43922 800 43938 856
rect 44106 800 44122 856
rect 44290 800 44306 856
rect 44474 800 44490 856
rect 44658 800 44766 856
rect 44934 800 44950 856
rect 45118 800 45134 856
rect 45302 800 45318 856
rect 45486 800 45502 856
rect 45670 800 45778 856
rect 45946 800 45962 856
rect 46130 800 46146 856
rect 46314 800 46330 856
rect 46498 800 46514 856
rect 46682 800 46790 856
rect 46958 800 46974 856
rect 47142 800 47158 856
rect 47326 800 47342 856
rect 47510 800 47526 856
rect 47694 800 47802 856
rect 47970 800 47986 856
rect 48154 800 48170 856
rect 48338 800 48354 856
rect 48522 800 48630 856
rect 48798 800 48814 856
rect 48982 800 48998 856
rect 49166 800 49182 856
rect 49350 800 49366 856
rect 49534 800 49642 856
rect 49810 800 49826 856
rect 49994 800 50010 856
rect 50178 800 50194 856
rect 50362 800 50378 856
rect 50546 800 50654 856
rect 50822 800 50838 856
rect 51006 800 51022 856
rect 51190 800 51206 856
rect 51374 800 51390 856
rect 51558 800 51666 856
rect 51834 800 51850 856
rect 52018 800 52034 856
rect 52202 800 52218 856
rect 52386 800 52494 856
rect 52662 800 52678 856
rect 52846 800 52862 856
rect 53030 800 53046 856
rect 53214 800 53230 856
rect 53398 800 53506 856
rect 53674 800 53690 856
rect 53858 800 53874 856
rect 54042 800 54058 856
rect 54226 800 54242 856
rect 54410 800 54518 856
rect 54686 800 54702 856
rect 54870 800 54886 856
rect 55054 800 55070 856
rect 55238 800 55254 856
rect 55422 800 55530 856
rect 55698 800 55714 856
rect 55882 800 55898 856
rect 56066 800 56082 856
rect 56250 800 56266 856
rect 56434 800 56542 856
rect 56710 800 56726 856
rect 56894 800 56910 856
rect 57078 800 57094 856
rect 57262 800 57370 856
rect 57538 800 57554 856
rect 57722 800 57738 856
rect 57906 800 57922 856
rect 58090 800 58106 856
rect 58274 800 58382 856
rect 58550 800 58566 856
rect 58734 800 58750 856
rect 58918 800 58934 856
rect 59102 800 59118 856
rect 59286 800 59394 856
rect 59562 800 59578 856
rect 59746 800 59762 856
rect 59930 800 59946 856
rect 60114 800 60130 856
rect 60298 800 60406 856
rect 60574 800 60590 856
rect 60758 800 60774 856
rect 60942 800 60958 856
rect 61126 800 61234 856
rect 61402 800 61418 856
rect 61586 800 61602 856
rect 61770 800 61786 856
rect 61954 800 61970 856
rect 62138 800 62246 856
rect 62414 800 62430 856
rect 62598 800 62614 856
rect 62782 800 62798 856
rect 62966 800 62982 856
rect 63150 800 63258 856
rect 63426 800 63442 856
rect 63610 800 63626 856
rect 63794 800 63810 856
rect 63978 800 63994 856
rect 64162 800 64270 856
rect 64438 800 64454 856
rect 64622 800 64638 856
rect 64806 800 64822 856
rect 64990 800 65006 856
rect 65174 800 65282 856
rect 65450 800 65466 856
rect 65634 800 65650 856
rect 65818 800 65834 856
rect 66002 800 66110 856
rect 66278 800 66294 856
rect 66462 800 66478 856
rect 66646 800 66662 856
rect 66830 800 66846 856
rect 67014 800 67122 856
rect 67290 800 67306 856
rect 67474 800 67490 856
rect 67658 800 67674 856
rect 67842 800 67858 856
rect 68026 800 68134 856
rect 68302 800 68318 856
rect 68486 800 68502 856
rect 68670 800 68686 856
rect 68854 800 68870 856
rect 69038 800 69146 856
rect 69314 800 69330 856
rect 69498 800 69514 856
rect 69682 800 69698 856
rect 69866 800 69974 856
rect 70142 800 70158 856
rect 70326 800 70342 856
rect 70510 800 70526 856
rect 70694 800 70710 856
rect 70878 800 70986 856
rect 71154 800 71170 856
rect 71338 800 71354 856
rect 71522 800 71538 856
rect 71706 800 71722 856
rect 71890 800 71998 856
rect 72166 800 72182 856
rect 72350 800 72366 856
rect 72534 800 72550 856
rect 72718 800 72734 856
rect 72902 800 73010 856
rect 73178 800 73194 856
rect 73362 800 73378 856
rect 73546 800 73562 856
rect 73730 800 73746 856
rect 73914 800 74022 856
rect 74190 800 74206 856
rect 74374 800 74390 856
rect 74558 800 74574 856
rect 74742 800 74850 856
rect 75018 800 75034 856
rect 75202 800 75218 856
rect 75386 800 75402 856
rect 75570 800 75586 856
rect 75754 800 75862 856
rect 76030 800 76046 856
rect 76214 800 76230 856
rect 76398 800 76414 856
rect 76582 800 76598 856
rect 76766 800 76874 856
rect 77042 800 77058 856
rect 77226 800 77242 856
rect 77410 800 77426 856
rect 77594 800 77610 856
rect 77778 800 77886 856
rect 78054 800 78070 856
rect 78238 800 78254 856
rect 78422 800 78438 856
rect 78606 800 78714 856
rect 78882 800 78898 856
rect 79066 800 79082 856
rect 79250 800 79266 856
rect 79434 800 79450 856
rect 79618 800 79726 856
rect 79894 800 79910 856
rect 80078 800 80094 856
rect 80262 800 80278 856
rect 80446 800 80462 856
rect 80630 800 80738 856
rect 80906 800 80922 856
rect 81090 800 81106 856
rect 81274 800 81290 856
rect 81458 800 81474 856
rect 81642 800 81750 856
rect 81918 800 81934 856
rect 82102 800 82118 856
rect 82286 800 82302 856
rect 82470 800 82486 856
rect 82654 800 82762 856
rect 82930 800 82946 856
rect 83114 800 83130 856
rect 83298 800 83314 856
rect 83482 800 83590 856
rect 83758 800 83774 856
rect 83942 800 83958 856
rect 84126 800 84142 856
rect 84310 800 84326 856
rect 84494 800 84602 856
rect 84770 800 84786 856
rect 84954 800 84970 856
rect 85138 800 85154 856
rect 85322 800 85338 856
rect 85506 800 85614 856
rect 85782 800 85798 856
rect 85966 800 85982 856
rect 86150 800 86166 856
rect 86334 800 86350 856
rect 86518 800 86626 856
rect 86794 800 86810 856
rect 86978 800 86994 856
rect 87162 800 87178 856
rect 87346 800 87454 856
rect 87622 800 87638 856
rect 87806 800 87822 856
rect 87990 800 88006 856
rect 88174 800 88190 856
rect 88358 800 88466 856
rect 88634 800 88650 856
rect 88818 800 88834 856
rect 89002 800 89018 856
rect 89186 800 89202 856
rect 89370 800 89478 856
rect 89646 800 89662 856
rect 89830 800 89846 856
rect 90014 800 90030 856
rect 90198 800 90214 856
rect 90382 800 90490 856
rect 90658 800 90674 856
rect 90842 800 90858 856
rect 91026 800 91042 856
rect 91210 800 91226 856
rect 91394 800 91502 856
rect 91670 800 91686 856
rect 91854 800 91870 856
rect 92038 800 92054 856
rect 92222 800 92330 856
rect 92498 800 92514 856
rect 92682 800 92698 856
rect 92866 800 92882 856
rect 93050 800 93066 856
rect 93234 800 93342 856
rect 93510 800 93526 856
rect 93694 800 93710 856
rect 93878 800 93894 856
rect 94062 800 94078 856
rect 94246 800 94354 856
rect 94522 800 94538 856
rect 94706 800 94722 856
rect 94890 800 94906 856
rect 95074 800 95090 856
rect 95258 800 95366 856
rect 95534 800 95550 856
rect 95718 800 95734 856
rect 95902 800 95918 856
rect 96086 800 96194 856
rect 96362 800 96378 856
rect 96546 800 96562 856
rect 96730 800 96746 856
rect 96914 800 96930 856
rect 97098 800 97206 856
rect 97374 800 97390 856
rect 97558 800 97574 856
rect 97742 800 97758 856
rect 97926 800 97942 856
rect 98110 800 98218 856
rect 98386 800 98402 856
rect 98570 800 98586 856
rect 98754 800 98770 856
rect 98938 800 98954 856
rect 99122 800 99230 856
rect 99398 800 99414 856
rect 99582 800 99598 856
rect 99766 800 99782 856
<< metal3 >>
rect 0 49920 800 50040
<< obsm3 >>
rect 800 50120 96688 97409
rect 880 49840 96688 50120
rect 800 2143 96688 49840
<< metal4 >>
rect 4208 2128 4528 97424
rect 4868 2176 5188 97376
rect 5528 2176 5848 97376
rect 6188 2176 6508 97376
rect 19568 2128 19888 97424
rect 20228 2176 20548 97376
rect 20888 2176 21208 97376
rect 21548 2176 21868 97376
rect 34928 2128 35248 97424
rect 35588 2176 35908 97376
rect 36248 2176 36568 97376
rect 36908 2176 37228 97376
rect 50288 2128 50608 97424
rect 50948 2176 51268 97376
rect 51608 2176 51928 97376
rect 52268 2176 52588 97376
rect 65648 2128 65968 97424
rect 66308 2176 66628 97376
rect 66968 2176 67288 97376
rect 67628 2176 67948 97376
rect 81008 2128 81328 97424
rect 81668 2176 81988 97376
rect 82328 2176 82648 97376
rect 82988 2176 83308 97376
rect 96368 2128 96688 97424
rect 97028 2176 97348 97376
rect 97688 2176 98008 97376
<< labels >>
rlabel metal2 s 386 99200 442 100000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 26422 99200 26478 100000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 28998 99200 29054 100000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 31666 99200 31722 100000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 34242 99200 34298 100000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 36818 99200 36874 100000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 39486 99200 39542 100000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 42062 99200 42118 100000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 44730 99200 44786 100000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 47306 99200 47362 100000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 49882 99200 49938 100000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2962 99200 3018 100000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 52550 99200 52606 100000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 55126 99200 55182 100000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 57702 99200 57758 100000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 60370 99200 60426 100000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 62946 99200 63002 100000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 65522 99200 65578 100000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 68190 99200 68246 100000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 70766 99200 70822 100000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 73342 99200 73398 100000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 76010 99200 76066 100000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5538 99200 5594 100000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 78586 99200 78642 100000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 81254 99200 81310 100000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 83830 99200 83886 100000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 86406 99200 86462 100000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 89074 99200 89130 100000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 91650 99200 91706 100000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 94226 99200 94282 100000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 96894 99200 96950 100000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8206 99200 8262 100000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10782 99200 10838 100000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13358 99200 13414 100000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 16026 99200 16082 100000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 18602 99200 18658 100000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 21178 99200 21234 100000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 23846 99200 23902 100000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1214 99200 1270 100000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 27342 99200 27398 100000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 29918 99200 29974 100000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 32494 99200 32550 100000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 35162 99200 35218 100000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 37738 99200 37794 100000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 40314 99200 40370 100000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 42982 99200 43038 100000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 45558 99200 45614 100000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 48134 99200 48190 100000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 50802 99200 50858 100000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3790 99200 3846 100000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 53378 99200 53434 100000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 55954 99200 56010 100000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 58622 99200 58678 100000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 61198 99200 61254 100000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 63866 99200 63922 100000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 66442 99200 66498 100000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 69018 99200 69074 100000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 71686 99200 71742 100000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 74262 99200 74318 100000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 76838 99200 76894 100000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6458 99200 6514 100000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 79506 99200 79562 100000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 82082 99200 82138 100000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 84658 99200 84714 100000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 87326 99200 87382 100000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 89902 99200 89958 100000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 92478 99200 92534 100000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 95146 99200 95202 100000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 97722 99200 97778 100000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9034 99200 9090 100000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 11610 99200 11666 100000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 14278 99200 14334 100000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 16854 99200 16910 100000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 19430 99200 19486 100000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 22098 99200 22154 100000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 24674 99200 24730 100000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2042 99200 2098 100000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 28170 99200 28226 100000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 30746 99200 30802 100000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 33414 99200 33470 100000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 35990 99200 36046 100000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 38566 99200 38622 100000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 41234 99200 41290 100000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 43810 99200 43866 100000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 46386 99200 46442 100000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 49054 99200 49110 100000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 51630 99200 51686 100000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4710 99200 4766 100000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 54298 99200 54354 100000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 56874 99200 56930 100000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 59450 99200 59506 100000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 62118 99200 62174 100000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 64694 99200 64750 100000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 67270 99200 67326 100000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 69938 99200 69994 100000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 72514 99200 72570 100000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 75090 99200 75146 100000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 77758 99200 77814 100000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7286 99200 7342 100000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 80334 99200 80390 100000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 82910 99200 82966 100000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 85578 99200 85634 100000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 88154 99200 88210 100000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 90822 99200 90878 100000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 93398 99200 93454 100000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 95974 99200 96030 100000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 98642 99200 98698 100000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9862 99200 9918 100000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 12530 99200 12586 100000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 15106 99200 15162 100000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 17774 99200 17830 100000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 20350 99200 20406 100000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 22926 99200 22982 100000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 25594 99200 25650 100000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 99470 99200 99526 100000 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 97446 0 97502 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 80334 0 80390 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 user_clock2
port 502 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 503 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 504 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 505 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[0]
port 506 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[10]
port 507 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[11]
port 508 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[12]
port 509 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[13]
port 510 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[14]
port 511 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[15]
port 512 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[16]
port 513 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[17]
port 514 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[18]
port 515 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_adr_i[19]
port 516 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[1]
port 517 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[20]
port 518 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[21]
port 519 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[22]
port 520 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[23]
port 521 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[24]
port 522 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[25]
port 523 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[26]
port 524 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[27]
port 525 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[28]
port 526 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[29]
port 527 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 528 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[30]
port 529 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[31]
port 530 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[3]
port 531 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[4]
port 532 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[5]
port 533 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[6]
port 534 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[7]
port 535 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[8]
port 536 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[9]
port 537 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 538 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 539 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[10]
port 540 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[11]
port 541 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[12]
port 542 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[13]
port 543 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[14]
port 544 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[15]
port 545 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[16]
port 546 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[17]
port 547 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[18]
port 548 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[19]
port 549 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[1]
port 550 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[20]
port 551 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[21]
port 552 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[22]
port 553 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[23]
port 554 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[24]
port 555 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[25]
port 556 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[26]
port 557 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[27]
port 558 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[28]
port 559 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[29]
port 560 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[2]
port 561 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[30]
port 562 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[31]
port 563 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[3]
port 564 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[4]
port 565 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[5]
port 566 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[6]
port 567 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[7]
port 568 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[8]
port 569 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[9]
port 570 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 571 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[10]
port 572 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[11]
port 573 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[12]
port 574 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[13]
port 575 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[14]
port 576 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[15]
port 577 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[16]
port 578 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[17]
port 579 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[18]
port 580 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[19]
port 581 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[1]
port 582 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[20]
port 583 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[21]
port 584 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[22]
port 585 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[23]
port 586 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[24]
port 587 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[25]
port 588 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[26]
port 589 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[27]
port 590 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[28]
port 591 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[29]
port 592 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[2]
port 593 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[30]
port 594 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[31]
port 595 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[3]
port 596 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[4]
port 597 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[5]
port 598 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[6]
port 599 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[7]
port 600 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[8]
port 601 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[9]
port 602 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 603 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 604 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[2]
port 605 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_sel_i[3]
port 606 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 607 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 608 nsew signal input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 613 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 97028 2176 97348 97376 6 vccd2
port 616 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 97376 6 vccd2
port 617 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 97376 6 vccd2
port 618 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 97376 6 vccd2
port 619 nsew power bidirectional
rlabel metal4 s 81668 2176 81988 97376 6 vssd2
port 620 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 97376 6 vssd2
port 621 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 97376 6 vssd2
port 622 nsew ground bidirectional
rlabel metal4 s 97688 2176 98008 97376 6 vdda1
port 623 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 97376 6 vdda1
port 624 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 97376 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 97376 6 vdda1
port 626 nsew power bidirectional
rlabel metal4 s 82328 2176 82648 97376 6 vssa1
port 627 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 97376 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 97376 6 vssa1
port 629 nsew ground bidirectional
rlabel metal4 s 67628 2176 67948 97376 6 vdda2
port 630 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 97376 6 vdda2
port 631 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 97376 6 vdda2
port 632 nsew power bidirectional
rlabel metal4 s 82988 2176 83308 97376 6 vssa2
port 633 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 97376 6 vssa2
port 634 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 97376 6 vssa2
port 635 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 100000 100000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 3023528
string GDS_START 126
<< end >>

